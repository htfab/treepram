magic
tech sky130A
magscale 1 2
timestamp 1635763811
<< locali >>
rect 66269 670871 66303 671449
rect 70961 670735 70995 671449
rect 79977 670803 80011 671449
rect 93685 670939 93719 671449
rect 134809 671211 134843 671449
rect 421573 671279 421607 671721
rect 449173 671143 449207 671245
rect 467205 671075 467239 671381
rect 490113 671007 490147 671381
rect 40877 30209 41061 30243
rect 31033 29631 31067 30005
rect 40877 29971 40911 30209
rect 39957 29937 40049 29971
rect 39865 29767 39899 29869
rect 39957 29291 39991 29937
rect 41153 29699 41187 30005
rect 50077 29971 50111 30209
rect 40693 29427 40727 29597
rect 39899 29257 39991 29291
rect 40601 29087 40635 29393
rect 46765 29155 46799 29937
rect 50261 29835 50295 29937
rect 50445 29291 50479 29733
rect 50537 29155 50571 29665
rect 105277 29427 105311 29665
rect 107485 29427 107519 29665
<< viali >>
rect 421573 671721 421607 671755
rect 66269 671449 66303 671483
rect 66269 670837 66303 670871
rect 70961 671449 70995 671483
rect 79977 671449 80011 671483
rect 93685 671449 93719 671483
rect 134809 671449 134843 671483
rect 467205 671381 467239 671415
rect 421573 671245 421607 671279
rect 449173 671245 449207 671279
rect 134809 671177 134843 671211
rect 449173 671109 449207 671143
rect 467205 671041 467239 671075
rect 490113 671381 490147 671415
rect 490113 670973 490147 671007
rect 93685 670905 93719 670939
rect 79977 670769 80011 670803
rect 70961 670701 70995 670735
rect 41061 30209 41095 30243
rect 50077 30209 50111 30243
rect 31033 30005 31067 30039
rect 40049 29937 40083 29971
rect 40877 29937 40911 29971
rect 41153 30005 41187 30039
rect 39865 29869 39899 29903
rect 39865 29733 39899 29767
rect 31033 29597 31067 29631
rect 41153 29665 41187 29699
rect 46765 29937 46799 29971
rect 50077 29937 50111 29971
rect 50261 29937 50295 29971
rect 40693 29597 40727 29631
rect 39865 29257 39899 29291
rect 40601 29393 40635 29427
rect 40693 29393 40727 29427
rect 50261 29801 50295 29835
rect 50445 29733 50479 29767
rect 50445 29257 50479 29291
rect 50537 29665 50571 29699
rect 46765 29121 46799 29155
rect 105277 29665 105311 29699
rect 105277 29393 105311 29427
rect 107485 29665 107519 29699
rect 107485 29393 107519 29427
rect 50537 29121 50571 29155
rect 40601 29053 40635 29087
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 329834 700992 329840 701004
rect 154172 700964 329840 700992
rect 154172 700952 154178 700964
rect 329834 700952 329840 700964
rect 329892 700952 329898 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 325694 700924 325700 700936
rect 137888 700896 325700 700924
rect 137888 700884 137894 700896
rect 325694 700884 325700 700896
rect 325752 700884 325758 700936
rect 257982 700816 257988 700868
rect 258040 700856 258046 700868
rect 462314 700856 462320 700868
rect 258040 700828 462320 700856
rect 258040 700816 258046 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 263502 700748 263508 700800
rect 263560 700788 263566 700800
rect 478506 700788 478512 700800
rect 263560 700760 478512 700788
rect 263560 700748 263566 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 343634 700720 343640 700732
rect 89220 700692 343640 700720
rect 89220 700680 89226 700692
rect 343634 700680 343640 700692
rect 343692 700680 343698 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 339494 700652 339500 700664
rect 73028 700624 339500 700652
rect 73028 700612 73034 700624
rect 339494 700612 339500 700624
rect 339552 700612 339558 700664
rect 244182 700544 244188 700596
rect 244240 700584 244246 700596
rect 527174 700584 527180 700596
rect 244240 700556 527180 700584
rect 244240 700544 244246 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 249702 700476 249708 700528
rect 249760 700516 249766 700528
rect 543458 700516 543464 700528
rect 249760 700488 543464 700516
rect 249760 700476 249766 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 347866 700448 347872 700460
rect 40552 700420 347872 700448
rect 40552 700408 40558 700420
rect 347866 700408 347872 700420
rect 347924 700408 347930 700460
rect 349798 700408 349804 700460
rect 349856 700448 349862 700460
rect 364978 700448 364984 700460
rect 349856 700420 364984 700448
rect 349856 700408 349862 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 357434 700380 357440 700392
rect 24360 700352 357440 700380
rect 24360 700340 24366 700352
rect 357434 700340 357440 700352
rect 357492 700340 357498 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 353294 700312 353300 700324
rect 8168 700284 353300 700312
rect 8168 700272 8174 700284
rect 353294 700272 353300 700284
rect 353352 700272 353358 700324
rect 356698 700272 356704 700324
rect 356756 700312 356762 700324
rect 494790 700312 494796 700324
rect 356756 700284 494796 700312
rect 356756 700272 356762 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 275922 700204 275928 700256
rect 275980 700244 275986 700256
rect 413646 700244 413652 700256
rect 275980 700216 413652 700244
rect 275980 700204 275986 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 271782 700136 271788 700188
rect 271840 700176 271846 700188
rect 397454 700176 397460 700188
rect 271840 700148 397460 700176
rect 271840 700136 271846 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 311894 700108 311900 700120
rect 202840 700080 311900 700108
rect 202840 700068 202846 700080
rect 311894 700068 311900 700080
rect 311952 700068 311958 700120
rect 218974 700000 218980 700052
rect 219032 700040 219038 700052
rect 316034 700040 316040 700052
rect 219032 700012 316040 700040
rect 219032 700000 219038 700012
rect 316034 700000 316040 700012
rect 316092 700000 316098 700052
rect 289722 699932 289728 699984
rect 289780 699972 289786 699984
rect 348786 699972 348792 699984
rect 289780 699944 348792 699972
rect 289780 699932 289786 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 285582 699864 285588 699916
rect 285640 699904 285646 699916
rect 332502 699904 332508 699916
rect 285640 699876 332508 699904
rect 285640 699864 285646 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 235166 699796 235172 699848
rect 235224 699836 235230 699848
rect 238018 699836 238024 699848
rect 235224 699808 238024 699836
rect 235224 699796 235230 699808
rect 238018 699796 238024 699808
rect 238076 699796 238082 699848
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 298094 699836 298100 699848
rect 267700 699808 298100 699836
rect 267700 699796 267706 699808
rect 298094 699796 298100 699808
rect 298152 699796 298158 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 302234 699768 302240 699780
rect 283892 699740 302240 699768
rect 283892 699728 283898 699740
rect 302234 699728 302240 699740
rect 302292 699728 302298 699780
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 555418 699660 555424 699712
rect 555476 699700 555482 699712
rect 559650 699700 559656 699712
rect 555476 699672 559656 699700
rect 555476 699660 555482 699672
rect 559650 699660 559656 699672
rect 559708 699660 559714 699712
rect 230382 696940 230388 696992
rect 230440 696980 230446 696992
rect 580166 696980 580172 696992
rect 230440 696952 580172 696980
rect 230440 696940 230446 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 235902 683204 235908 683256
rect 235960 683244 235966 683256
rect 580166 683244 580172 683256
rect 235960 683216 580172 683244
rect 235960 683204 235966 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 361574 683176 361580 683188
rect 3476 683148 361580 683176
rect 3476 683136 3482 683148
rect 361574 683136 361580 683148
rect 361632 683136 361638 683188
rect 294230 675996 294236 676048
rect 294288 676036 294294 676048
rect 299474 676036 299480 676048
rect 294288 676008 299480 676036
rect 294288 675996 294294 676008
rect 299474 675996 299480 676008
rect 299532 675996 299538 676048
rect 280522 675928 280528 675980
rect 280580 675968 280586 675980
rect 349798 675968 349804 675980
rect 280580 675940 349804 675968
rect 280580 675928 280586 675940
rect 349798 675928 349804 675940
rect 349856 675928 349862 675980
rect 238018 675860 238024 675912
rect 238076 675900 238082 675912
rect 307846 675900 307852 675912
rect 238076 675872 307852 675900
rect 238076 675860 238082 675872
rect 307846 675860 307852 675872
rect 307904 675860 307910 675912
rect 253106 675792 253112 675844
rect 253164 675832 253170 675844
rect 356698 675832 356704 675844
rect 253164 675804 356704 675832
rect 253164 675792 253170 675804
rect 356698 675792 356704 675804
rect 356756 675792 356762 675844
rect 171042 675724 171048 675776
rect 171100 675764 171106 675776
rect 321554 675764 321560 675776
rect 171100 675736 321560 675764
rect 171100 675724 171106 675736
rect 321554 675724 321560 675736
rect 321612 675724 321618 675776
rect 266814 675656 266820 675708
rect 266872 675696 266878 675708
rect 429194 675696 429200 675708
rect 266872 675668 429200 675696
rect 266872 675656 266878 675668
rect 429194 675656 429200 675668
rect 429252 675656 429258 675708
rect 106182 675588 106188 675640
rect 106240 675628 106246 675640
rect 335262 675628 335268 675640
rect 106240 675600 335268 675628
rect 106240 675588 106246 675600
rect 335262 675588 335268 675600
rect 335320 675588 335326 675640
rect 239490 675520 239496 675572
rect 239548 675560 239554 675572
rect 555418 675560 555424 675572
rect 239548 675532 555424 675560
rect 239548 675520 239554 675532
rect 555418 675520 555424 675532
rect 555476 675520 555482 675572
rect 175550 675452 175556 675504
rect 175608 675492 175614 675504
rect 554130 675492 554136 675504
rect 175608 675464 554136 675492
rect 175608 675452 175614 675464
rect 554130 675452 554136 675464
rect 554188 675452 554194 675504
rect 157334 675384 157340 675436
rect 157392 675424 157398 675436
rect 558270 675424 558276 675436
rect 157392 675396 558276 675424
rect 157392 675384 157398 675396
rect 558270 675384 558276 675396
rect 558328 675384 558334 675436
rect 143626 675316 143632 675368
rect 143684 675356 143690 675368
rect 576210 675356 576216 675368
rect 143684 675328 576216 675356
rect 143684 675316 143690 675328
rect 576210 675316 576216 675328
rect 576268 675316 576274 675368
rect 130010 675248 130016 675300
rect 130068 675288 130074 675300
rect 574830 675288 574836 675300
rect 130068 675260 574836 675288
rect 130068 675248 130074 675260
rect 574830 675248 574836 675260
rect 574888 675248 574894 675300
rect 25590 675180 25596 675232
rect 25648 675220 25654 675232
rect 499482 675220 499488 675232
rect 25648 675192 499488 675220
rect 25648 675180 25654 675192
rect 499482 675180 499488 675192
rect 499540 675180 499546 675232
rect 29730 675112 29736 675164
rect 29788 675152 29794 675164
rect 513098 675152 513104 675164
rect 29788 675124 513104 675152
rect 29788 675112 29794 675124
rect 513098 675112 513104 675124
rect 513156 675112 513162 675164
rect 75270 675044 75276 675096
rect 75328 675084 75334 675096
rect 565078 675084 565084 675096
rect 75328 675056 565084 675084
rect 75328 675044 75334 675056
rect 565078 675044 565084 675056
rect 565136 675044 565142 675096
rect 43346 674976 43352 675028
rect 43404 675016 43410 675028
rect 552658 675016 552664 675028
rect 43404 674988 552664 675016
rect 43404 674976 43410 674988
rect 552658 674976 552664 674988
rect 552716 674976 552722 675028
rect 7558 674908 7564 674960
rect 7616 674948 7622 674960
rect 526806 674948 526812 674960
rect 7616 674920 526812 674948
rect 7616 674908 7622 674920
rect 526806 674908 526812 674920
rect 526864 674908 526870 674960
rect 52454 674840 52460 674892
rect 52512 674880 52518 674892
rect 576118 674880 576124 674892
rect 52512 674852 576124 674880
rect 52512 674840 52518 674852
rect 576118 674840 576124 674852
rect 576176 674840 576182 674892
rect 218054 674772 218060 674824
rect 218112 674812 218118 674824
rect 412818 674812 412824 674824
rect 218112 674784 412824 674812
rect 218112 674772 218118 674784
rect 412818 674772 412824 674784
rect 412876 674772 412882 674824
rect 152826 674704 152832 674756
rect 152884 674744 152890 674756
rect 382274 674744 382280 674756
rect 152884 674716 382280 674744
rect 152884 674704 152890 674716
rect 382274 674704 382280 674716
rect 382332 674704 382338 674756
rect 125410 674636 125416 674688
rect 125468 674676 125474 674688
rect 368658 674676 368664 674688
rect 125468 674648 368664 674676
rect 125468 674636 125474 674648
rect 368658 674636 368664 674648
rect 368716 674636 368722 674688
rect 200114 674568 200120 674620
rect 200172 674608 200178 674620
rect 481174 674608 481180 674620
rect 200172 674580 481180 674608
rect 200172 674568 200178 674580
rect 481174 674568 481180 674580
rect 481232 674568 481238 674620
rect 14550 674500 14556 674552
rect 14608 674540 14614 674552
rect 408218 674540 408224 674552
rect 14608 674512 408224 674540
rect 14608 674500 14614 674512
rect 408218 674500 408224 674512
rect 408276 674500 408282 674552
rect 180150 674432 180156 674484
rect 180208 674472 180214 674484
rect 572070 674472 572076 674484
rect 180208 674444 572076 674472
rect 180208 674432 180214 674444
rect 572070 674432 572076 674444
rect 572128 674432 572134 674484
rect 166442 674364 166448 674416
rect 166500 674404 166506 674416
rect 571978 674404 571984 674416
rect 166500 674376 571984 674404
rect 166500 674364 166506 674376
rect 571978 674364 571984 674376
rect 572036 674364 572042 674416
rect 111702 674296 111708 674348
rect 111760 674336 111766 674348
rect 155770 674336 155776 674348
rect 111760 674308 155776 674336
rect 111760 674296 111766 674308
rect 155770 674296 155776 674308
rect 155828 674296 155834 674348
rect 161934 674296 161940 674348
rect 161992 674336 161998 674348
rect 570598 674336 570604 674348
rect 161992 674308 570604 674336
rect 161992 674296 161998 674308
rect 570598 674296 570604 674308
rect 570656 674296 570662 674348
rect 26878 674228 26884 674280
rect 26936 674268 26942 674280
rect 440142 674268 440148 674280
rect 26936 674240 440148 674268
rect 26936 674228 26942 674240
rect 440142 674228 440148 674240
rect 440200 674228 440206 674280
rect 17310 674160 17316 674212
rect 17368 674200 17374 674212
rect 435542 674200 435548 674212
rect 17368 674172 435548 674200
rect 17368 674160 17374 674172
rect 435542 674160 435548 674172
rect 435600 674160 435606 674212
rect 148226 674092 148232 674144
rect 148284 674132 148290 674144
rect 565170 674132 565176 674144
rect 148284 674104 565176 674132
rect 148284 674092 148290 674104
rect 565170 674092 565176 674104
rect 565228 674092 565234 674144
rect 18690 674024 18696 674076
rect 18748 674064 18754 674076
rect 449250 674064 449256 674076
rect 18748 674036 449256 674064
rect 18748 674024 18754 674036
rect 449250 674024 449256 674036
rect 449308 674024 449314 674076
rect 11790 673956 11796 674008
rect 11848 673996 11854 674008
rect 453850 673996 453856 674008
rect 11848 673968 453856 673996
rect 11848 673956 11854 673968
rect 453850 673956 453856 673968
rect 453908 673956 453914 674008
rect 120902 673888 120908 673940
rect 120960 673928 120966 673940
rect 561030 673928 561036 673940
rect 120960 673900 561036 673928
rect 120960 673888 120966 673900
rect 561030 673888 561036 673900
rect 561088 673888 561094 673940
rect 31018 673820 31024 673872
rect 31076 673860 31082 673872
rect 476666 673860 476672 673872
rect 31076 673832 476672 673860
rect 31076 673820 31082 673832
rect 476666 673820 476672 673832
rect 476724 673820 476730 673872
rect 107194 673752 107200 673804
rect 107252 673792 107258 673804
rect 555510 673792 555516 673804
rect 107252 673764 555516 673792
rect 107252 673752 107258 673764
rect 555510 673752 555516 673764
rect 555568 673752 555574 673804
rect 17218 673684 17224 673736
rect 17276 673724 17282 673736
rect 494882 673724 494888 673736
rect 17276 673696 494888 673724
rect 17276 673684 17282 673696
rect 494882 673684 494888 673696
rect 494940 673684 494946 673736
rect 22738 673616 22744 673668
rect 22796 673656 22802 673668
rect 503990 673656 503996 673668
rect 22796 673628 503996 673656
rect 22796 673616 22802 673628
rect 503990 673616 503996 673628
rect 504048 673616 504054 673668
rect 25498 673548 25504 673600
rect 25556 673588 25562 673600
rect 517698 673588 517704 673600
rect 25556 673560 517704 673588
rect 25556 673548 25562 673560
rect 517698 673548 517704 673560
rect 517756 673548 517762 673600
rect 4890 673480 4896 673532
rect 4948 673520 4954 673532
rect 522206 673520 522212 673532
rect 4948 673492 522212 673520
rect 4948 673480 4954 673492
rect 522206 673480 522212 673492
rect 522264 673480 522270 673532
rect 212074 673344 212080 673396
rect 212132 673384 212138 673396
rect 558362 673384 558368 673396
rect 212132 673356 558368 673384
rect 212132 673344 212138 673356
rect 558362 673344 558368 673356
rect 558420 673344 558426 673396
rect 3510 673276 3516 673328
rect 3568 673316 3574 673328
rect 200114 673316 200120 673328
rect 3568 673288 200120 673316
rect 3568 673276 3574 673288
rect 200114 673276 200120 673288
rect 200172 673276 200178 673328
rect 225782 673276 225788 673328
rect 225840 673316 225846 673328
rect 579522 673316 579528 673328
rect 225840 673288 579528 673316
rect 225840 673276 225846 673288
rect 579522 673276 579528 673288
rect 579580 673276 579586 673328
rect 198366 673208 198372 673260
rect 198424 673248 198430 673260
rect 556982 673248 556988 673260
rect 198424 673220 556988 673248
rect 198424 673208 198430 673220
rect 556982 673208 556988 673220
rect 557040 673208 557046 673260
rect 7742 673140 7748 673192
rect 7800 673180 7806 673192
rect 376294 673180 376300 673192
rect 7800 673152 376300 673180
rect 7800 673140 7806 673152
rect 376294 673140 376300 673152
rect 376352 673140 376358 673192
rect 184750 673072 184756 673124
rect 184808 673112 184814 673124
rect 554222 673112 554228 673124
rect 184808 673084 554228 673112
rect 184808 673072 184814 673084
rect 554222 673072 554228 673084
rect 554280 673072 554286 673124
rect 11882 673004 11888 673056
rect 11940 673044 11946 673056
rect 390002 673044 390008 673056
rect 11940 673016 390008 673044
rect 11940 673004 11946 673016
rect 390002 673004 390008 673016
rect 390060 673004 390066 673056
rect 171042 672936 171048 672988
rect 171100 672976 171106 672988
rect 552750 672976 552756 672988
rect 171100 672948 552756 672976
rect 171100 672936 171106 672948
rect 552750 672936 552756 672948
rect 552808 672936 552814 672988
rect 14642 672868 14648 672920
rect 14700 672908 14706 672920
rect 403618 672908 403624 672920
rect 14700 672880 403624 672908
rect 14700 672868 14706 672880
rect 403618 672868 403624 672880
rect 403676 672868 403682 672920
rect 16022 672800 16028 672852
rect 16080 672840 16086 672852
rect 417326 672840 417332 672852
rect 16080 672812 417332 672840
rect 16080 672800 16086 672812
rect 417326 672800 417332 672812
rect 417384 672800 417390 672852
rect 155770 672732 155776 672784
rect 155828 672772 155834 672784
rect 580258 672772 580264 672784
rect 155828 672744 580264 672772
rect 155828 672732 155834 672744
rect 580258 672732 580264 672744
rect 580316 672732 580322 672784
rect 17402 672664 17408 672716
rect 17460 672704 17466 672716
rect 431034 672704 431040 672716
rect 17460 672676 431040 672704
rect 17460 672664 17466 672676
rect 431034 672664 431040 672676
rect 431092 672664 431098 672716
rect 139118 672596 139124 672648
rect 139176 672636 139182 672648
rect 556890 672636 556896 672648
rect 139176 672608 556896 672636
rect 139176 672596 139182 672608
rect 556890 672596 556896 672608
rect 556948 672596 556954 672648
rect 18782 672528 18788 672580
rect 18840 672568 18846 672580
rect 444742 672568 444748 672580
rect 18840 672540 444748 672568
rect 18840 672528 18846 672540
rect 444742 672528 444748 672540
rect 444800 672528 444806 672580
rect 21450 672460 21456 672512
rect 21508 672500 21514 672512
rect 458358 672500 458364 672512
rect 21508 672472 458364 672500
rect 21508 672460 21514 672472
rect 458358 672460 458364 672472
rect 458416 672460 458422 672512
rect 31110 672392 31116 672444
rect 31168 672432 31174 672444
rect 472066 672432 472072 672444
rect 31168 672404 472072 672432
rect 31168 672392 31174 672404
rect 472066 672392 472072 672404
rect 472124 672392 472130 672444
rect 22830 672324 22836 672376
rect 22888 672364 22894 672376
rect 485774 672364 485780 672376
rect 22888 672336 485780 672364
rect 22888 672324 22894 672336
rect 485774 672324 485780 672336
rect 485832 672324 485838 672376
rect 98086 672256 98092 672308
rect 98144 672296 98150 672308
rect 578878 672296 578884 672308
rect 98144 672268 578884 672296
rect 98144 672256 98150 672268
rect 578878 672256 578884 672268
rect 578936 672256 578942 672308
rect 84378 672188 84384 672240
rect 84436 672228 84442 672240
rect 569218 672228 569224 672240
rect 84436 672200 569224 672228
rect 84436 672188 84442 672200
rect 569218 672188 569224 672200
rect 569276 672188 569282 672240
rect 61562 672120 61568 672172
rect 61620 672160 61626 672172
rect 562318 672160 562324 672172
rect 61620 672132 562324 672160
rect 61620 672120 61626 672132
rect 562318 672120 562324 672132
rect 562376 672120 562382 672172
rect 3418 672052 3424 672104
rect 3476 672092 3482 672104
rect 508590 672092 508596 672104
rect 3476 672064 508596 672092
rect 3476 672052 3482 672064
rect 508590 672052 508596 672064
rect 508648 672052 508654 672104
rect 3602 671984 3608 672036
rect 3660 672024 3666 672036
rect 218054 672024 218060 672036
rect 3660 671996 218060 672024
rect 3660 671984 3666 671996
rect 218054 671984 218060 671996
rect 218112 671984 218118 672036
rect 221458 671984 221464 672036
rect 221516 672024 221522 672036
rect 557074 672024 557080 672036
rect 221516 671996 557080 672024
rect 221516 671984 221522 671996
rect 557074 671984 557080 671996
rect 557132 671984 557138 672036
rect 27062 671916 27068 671968
rect 27120 671956 27126 671968
rect 367278 671956 367284 671968
rect 27120 671928 367284 671956
rect 27120 671916 27126 671928
rect 367278 671916 367284 671928
rect 367336 671916 367342 671968
rect 368658 671916 368664 671968
rect 368716 671956 368722 671968
rect 580350 671956 580356 671968
rect 368716 671928 580356 671956
rect 368716 671916 368722 671928
rect 580350 671916 580356 671928
rect 580408 671916 580414 671968
rect 28350 671848 28356 671900
rect 28408 671888 28414 671900
rect 380986 671888 380992 671900
rect 28408 671860 380992 671888
rect 28408 671848 28414 671860
rect 380986 671848 380992 671860
rect 381044 671848 381050 671900
rect 217042 671780 217048 671832
rect 217100 671820 217106 671832
rect 569494 671820 569500 671832
rect 217100 671792 569500 671820
rect 217100 671780 217106 671792
rect 569494 671780 569500 671792
rect 569552 671780 569558 671832
rect 26970 671712 26976 671764
rect 27028 671752 27034 671764
rect 385126 671752 385132 671764
rect 27028 671724 385132 671752
rect 27028 671712 27034 671724
rect 385126 671712 385132 671724
rect 385184 671712 385190 671764
rect 421558 671752 421564 671764
rect 421519 671724 421564 671752
rect 421558 671712 421564 671724
rect 421616 671712 421622 671764
rect 207842 671644 207848 671696
rect 207900 671684 207906 671696
rect 569402 671684 569408 671696
rect 207900 671656 569408 671684
rect 207900 671644 207906 671656
rect 569402 671644 569408 671656
rect 569460 671644 569466 671696
rect 203242 671576 203248 671628
rect 203300 671616 203306 671628
rect 566642 671616 566648 671628
rect 203300 671588 566648 671616
rect 203300 671576 203306 671588
rect 566642 671576 566648 671588
rect 566700 671576 566706 671628
rect 3326 671508 3332 671560
rect 3384 671548 3390 671560
rect 371326 671548 371332 671560
rect 3384 671520 371332 671548
rect 3384 671508 3390 671520
rect 371326 671508 371332 671520
rect 371384 671508 371390 671560
rect 382274 671508 382280 671560
rect 382332 671548 382338 671560
rect 580442 671548 580448 671560
rect 382332 671520 580448 671548
rect 382332 671508 382338 671520
rect 580442 671508 580448 671520
rect 580500 671508 580506 671560
rect 66254 671480 66260 671492
rect 66215 671452 66260 671480
rect 66254 671440 66260 671452
rect 66312 671440 66318 671492
rect 70946 671480 70952 671492
rect 70907 671452 70952 671480
rect 70946 671440 70952 671452
rect 71004 671440 71010 671492
rect 79962 671480 79968 671492
rect 79923 671452 79968 671480
rect 79962 671440 79968 671452
rect 80020 671440 80026 671492
rect 93670 671480 93676 671492
rect 93631 671452 93676 671480
rect 93670 671440 93676 671452
rect 93728 671440 93734 671492
rect 134794 671480 134800 671492
rect 134755 671452 134800 671480
rect 134794 671440 134800 671452
rect 134852 671440 134858 671492
rect 194226 671440 194232 671492
rect 194284 671480 194290 671492
rect 578970 671480 578976 671492
rect 194284 671452 578976 671480
rect 194284 671440 194290 671452
rect 578970 671440 578976 671452
rect 579028 671440 579034 671492
rect 7650 671372 7656 671424
rect 7708 671412 7714 671424
rect 398834 671412 398840 671424
rect 7708 671384 398840 671412
rect 7708 671372 7714 671384
rect 398834 671372 398840 671384
rect 398892 671372 398898 671424
rect 426250 671412 426256 671424
rect 412606 671384 426256 671412
rect 28258 671304 28264 671356
rect 28316 671344 28322 671356
rect 412606 671344 412634 671384
rect 426250 671372 426256 671384
rect 426308 671372 426314 671424
rect 462590 671412 462596 671424
rect 460906 671384 462596 671412
rect 28316 671316 412634 671344
rect 28316 671304 28322 671316
rect 15930 671236 15936 671288
rect 15988 671276 15994 671288
rect 421561 671279 421619 671285
rect 421561 671276 421573 671279
rect 15988 671248 421573 671276
rect 15988 671236 15994 671248
rect 421561 671245 421573 671248
rect 421607 671245 421619 671279
rect 421561 671239 421619 671245
rect 449161 671279 449219 671285
rect 449161 671245 449173 671279
rect 449207 671276 449219 671279
rect 460906 671276 460934 671384
rect 462590 671372 462596 671384
rect 462648 671372 462654 671424
rect 467190 671412 467196 671424
rect 467151 671384 467196 671412
rect 467190 671372 467196 671384
rect 467248 671372 467254 671424
rect 490098 671412 490104 671424
rect 490059 671384 490104 671412
rect 490098 671372 490104 671384
rect 490156 671372 490162 671424
rect 449207 671248 460934 671276
rect 449207 671245 449219 671248
rect 449161 671239 449219 671245
rect 134797 671211 134855 671217
rect 134797 671177 134809 671211
rect 134843 671208 134855 671211
rect 562410 671208 562416 671220
rect 134843 671180 449296 671208
rect 134843 671177 134855 671180
rect 134797 671171 134855 671177
rect 21358 671100 21364 671152
rect 21416 671140 21422 671152
rect 449161 671143 449219 671149
rect 449161 671140 449173 671143
rect 21416 671112 449173 671140
rect 21416 671100 21422 671112
rect 449161 671109 449173 671112
rect 449207 671109 449219 671143
rect 449268 671140 449296 671180
rect 454006 671180 562416 671208
rect 454006 671140 454034 671180
rect 562410 671168 562416 671180
rect 562468 671168 562474 671220
rect 449268 671112 454034 671140
rect 449161 671103 449219 671109
rect 10318 671032 10324 671084
rect 10376 671072 10382 671084
rect 467193 671075 467251 671081
rect 467193 671072 467205 671075
rect 10376 671044 467205 671072
rect 10376 671032 10382 671044
rect 467193 671041 467205 671044
rect 467239 671041 467251 671075
rect 467193 671035 467251 671041
rect 14458 670964 14464 671016
rect 14516 671004 14522 671016
rect 490101 671007 490159 671013
rect 490101 671004 490113 671007
rect 14516 670976 490113 671004
rect 14516 670964 14522 670976
rect 490101 670973 490113 670976
rect 490147 670973 490159 671007
rect 490101 670967 490159 670973
rect 93673 670939 93731 670945
rect 93673 670905 93685 670939
rect 93719 670936 93731 670939
rect 573358 670936 573364 670948
rect 93719 670908 573364 670936
rect 93719 670905 93731 670908
rect 93673 670899 93731 670905
rect 573358 670896 573364 670908
rect 573416 670896 573422 670948
rect 66257 670871 66315 670877
rect 66257 670837 66269 670871
rect 66303 670868 66315 670871
rect 558178 670868 558184 670880
rect 66303 670840 558184 670868
rect 66303 670837 66315 670840
rect 66257 670831 66315 670837
rect 558178 670828 558184 670840
rect 558236 670828 558242 670880
rect 79965 670803 80023 670809
rect 79965 670769 79977 670803
rect 80011 670800 80023 670803
rect 574738 670800 574744 670812
rect 80011 670772 574744 670800
rect 80011 670769 80023 670772
rect 79965 670763 80023 670769
rect 574738 670760 574744 670772
rect 574796 670760 574802 670812
rect 70949 670735 71007 670741
rect 70949 670701 70961 670735
rect 70995 670732 71007 670735
rect 566458 670732 566464 670744
rect 70995 670704 566464 670732
rect 70995 670701 71007 670704
rect 70949 670695 71007 670701
rect 566458 670692 566464 670704
rect 566516 670692 566522 670744
rect 3326 658180 3332 658232
rect 3384 658220 3390 658232
rect 27062 658220 27068 658232
rect 3384 658192 27068 658220
rect 3384 658180 3390 658192
rect 27062 658180 27068 658192
rect 27120 658180 27126 658232
rect 569494 644376 569500 644428
rect 569552 644416 569558 644428
rect 580166 644416 580172 644428
rect 569552 644388 580172 644416
rect 569552 644376 569558 644388
rect 580166 644376 580172 644388
rect 580224 644376 580230 644428
rect 3326 633360 3332 633412
rect 3384 633400 3390 633412
rect 7742 633400 7748 633412
rect 3384 633372 7748 633400
rect 3384 633360 3390 633372
rect 7742 633360 7748 633372
rect 7800 633360 7806 633412
rect 557074 632000 557080 632052
rect 557132 632040 557138 632052
rect 579706 632040 579712 632052
rect 557132 632012 579712 632040
rect 557132 632000 557138 632012
rect 579706 632000 579712 632012
rect 579764 632000 579770 632052
rect 3326 619556 3332 619608
rect 3384 619596 3390 619608
rect 26970 619596 26976 619608
rect 3384 619568 26976 619596
rect 3384 619556 3390 619568
rect 26970 619556 26976 619568
rect 27028 619556 27034 619608
rect 558362 618196 558368 618248
rect 558420 618236 558426 618248
rect 579798 618236 579804 618248
rect 558420 618208 579804 618236
rect 558420 618196 558426 618208
rect 579798 618196 579804 618208
rect 579856 618196 579862 618248
rect 3050 607112 3056 607164
rect 3108 607152 3114 607164
rect 28350 607152 28356 607164
rect 3108 607124 28356 607152
rect 3108 607112 3114 607124
rect 28350 607112 28356 607124
rect 28408 607112 28414 607164
rect 566642 591948 566648 592000
rect 566700 591988 566706 592000
rect 580166 591988 580172 592000
rect 566700 591960 580172 591988
rect 566700 591948 566706 591960
rect 580166 591948 580172 591960
rect 580224 591948 580230 592000
rect 3326 580932 3332 580984
rect 3384 580972 3390 580984
rect 11882 580972 11888 580984
rect 3384 580944 11888 580972
rect 3384 580932 3390 580944
rect 11882 580932 11888 580944
rect 11940 580932 11946 580984
rect 569402 578144 569408 578196
rect 569460 578184 569466 578196
rect 580166 578184 580172 578196
rect 569460 578156 580172 578184
rect 569460 578144 569466 578156
rect 580166 578144 580172 578156
rect 580224 578144 580230 578196
rect 3142 567060 3148 567112
rect 3200 567100 3206 567112
rect 7650 567100 7656 567112
rect 3200 567072 7656 567100
rect 3200 567060 3206 567072
rect 7650 567060 7656 567072
rect 7708 567060 7714 567112
rect 556982 564340 556988 564392
rect 557040 564380 557046 564392
rect 580166 564380 580172 564392
rect 557040 564352 580172 564380
rect 557040 564340 557046 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 2958 554684 2964 554736
rect 3016 554724 3022 554736
rect 10410 554724 10416 554736
rect 3016 554696 10416 554724
rect 3016 554684 3022 554696
rect 10410 554684 10416 554696
rect 10468 554684 10474 554736
rect 552842 538160 552848 538212
rect 552900 538200 552906 538212
rect 580166 538200 580172 538212
rect 552900 538172 580172 538200
rect 552900 538160 552906 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 3142 528504 3148 528556
rect 3200 528544 3206 528556
rect 14642 528544 14648 528556
rect 3200 528516 14648 528544
rect 3200 528504 3206 528516
rect 14642 528504 14648 528516
rect 14700 528504 14706 528556
rect 554222 511912 554228 511964
rect 554280 511952 554286 511964
rect 580166 511952 580172 511964
rect 554280 511924 580172 511952
rect 554280 511912 554286 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 2958 502256 2964 502308
rect 3016 502296 3022 502308
rect 14550 502296 14556 502308
rect 3016 502268 14556 502296
rect 3016 502256 3022 502268
rect 14550 502256 14556 502268
rect 14608 502256 14614 502308
rect 554130 485732 554136 485784
rect 554188 485772 554194 485784
rect 580166 485772 580172 485784
rect 554188 485744 580172 485772
rect 554188 485732 554194 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 3234 476008 3240 476060
rect 3292 476048 3298 476060
rect 16022 476048 16028 476060
rect 3292 476020 16028 476048
rect 3292 476008 3298 476020
rect 16022 476008 16028 476020
rect 16080 476008 16086 476060
rect 572070 471928 572076 471980
rect 572128 471968 572134 471980
rect 580166 471968 580172 471980
rect 572128 471940 580172 471968
rect 572128 471928 572134 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 3050 463632 3056 463684
rect 3108 463672 3114 463684
rect 28258 463672 28264 463684
rect 3108 463644 28264 463672
rect 3108 463632 3114 463644
rect 28258 463632 28264 463644
rect 28316 463632 28322 463684
rect 552750 458124 552756 458176
rect 552808 458164 552814 458176
rect 580166 458164 580172 458176
rect 552808 458136 580172 458164
rect 552808 458124 552814 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 15930 449868 15936 449880
rect 3384 449840 15936 449868
rect 3384 449828 3390 449840
rect 15930 449828 15936 449840
rect 15988 449828 15994 449880
rect 570598 431876 570604 431928
rect 570656 431916 570662 431928
rect 580166 431916 580172 431928
rect 570656 431888 580172 431916
rect 570656 431876 570662 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 17402 423620 17408 423632
rect 3384 423592 17408 423620
rect 3384 423580 3390 423592
rect 17402 423580 17408 423592
rect 17460 423580 17466 423632
rect 571978 419432 571984 419484
rect 572036 419472 572042 419484
rect 579706 419472 579712 419484
rect 572036 419444 579712 419472
rect 572036 419432 572042 419444
rect 579706 419432 579712 419444
rect 579764 419432 579770 419484
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 26878 411244 26884 411256
rect 3016 411216 26884 411244
rect 3016 411204 3022 411216
rect 26878 411204 26884 411216
rect 26936 411204 26942 411256
rect 558270 405628 558276 405680
rect 558328 405668 558334 405680
rect 579798 405668 579804 405680
rect 558328 405640 579804 405668
rect 558328 405628 558334 405640
rect 579798 405628 579804 405640
rect 579856 405628 579862 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 17310 398800 17316 398812
rect 3384 398772 17316 398800
rect 3384 398760 3390 398772
rect 17310 398760 17316 398772
rect 17368 398760 17374 398812
rect 565170 379448 565176 379500
rect 565228 379488 565234 379500
rect 579798 379488 579804 379500
rect 565228 379460 579804 379488
rect 565228 379448 565234 379460
rect 579798 379448 579804 379460
rect 579856 379448 579862 379500
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 18782 372552 18788 372564
rect 3384 372524 18788 372552
rect 3384 372512 3390 372524
rect 18782 372512 18788 372524
rect 18840 372512 18846 372564
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 11790 358748 11796 358760
rect 3384 358720 11796 358748
rect 3384 358708 3390 358720
rect 11790 358708 11796 358720
rect 11848 358708 11854 358760
rect 576210 353200 576216 353252
rect 576268 353240 576274 353252
rect 580166 353240 580172 353252
rect 576268 353212 580172 353240
rect 576268 353200 576274 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 18690 346372 18696 346384
rect 3384 346344 18696 346372
rect 3384 346332 3390 346344
rect 18690 346332 18696 346344
rect 18748 346332 18754 346384
rect 562410 325592 562416 325644
rect 562468 325632 562474 325644
rect 580166 325632 580172 325644
rect 562468 325604 580172 325632
rect 562468 325592 562474 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 21450 320124 21456 320136
rect 3384 320096 21456 320124
rect 3384 320084 3390 320096
rect 21450 320084 21456 320096
rect 21508 320084 21514 320136
rect 556890 313216 556896 313268
rect 556948 313256 556954 313268
rect 580166 313256 580172 313268
rect 556948 313228 580172 313256
rect 556948 313216 556954 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 10318 306320 10324 306332
rect 3384 306292 10324 306320
rect 3384 306280 3390 306292
rect 10318 306280 10324 306292
rect 10376 306280 10382 306332
rect 574830 299412 574836 299464
rect 574888 299452 574894 299464
rect 580166 299452 580172 299464
rect 574888 299424 580172 299452
rect 574888 299412 574894 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3326 293904 3332 293956
rect 3384 293944 3390 293956
rect 21358 293944 21364 293956
rect 3384 293916 21364 293944
rect 3384 293904 3390 293916
rect 21358 293904 21364 293916
rect 21416 293904 21422 293956
rect 561030 273164 561036 273216
rect 561088 273204 561094 273216
rect 580166 273204 580172 273216
rect 561088 273176 580172 273204
rect 561088 273164 561094 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 31110 267696 31116 267708
rect 3016 267668 31116 267696
rect 3016 267656 3022 267668
rect 31110 267656 31116 267668
rect 31168 267656 31174 267708
rect 573450 245556 573456 245608
rect 573508 245596 573514 245608
rect 580166 245596 580172 245608
rect 573508 245568 580172 245596
rect 573508 245556 573514 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 31018 241448 31024 241460
rect 3568 241420 31024 241448
rect 3568 241408 3574 241420
rect 31018 241408 31024 241420
rect 31076 241408 31082 241460
rect 555510 233180 555516 233232
rect 555568 233220 555574 233232
rect 580166 233220 580172 233232
rect 555568 233192 580172 233220
rect 555568 233180 555574 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 22830 215268 22836 215280
rect 3384 215240 22836 215268
rect 3384 215228 3390 215240
rect 22830 215228 22836 215240
rect 22888 215228 22894 215280
rect 569310 206932 569316 206984
rect 569368 206972 569374 206984
rect 579798 206972 579804 206984
rect 569368 206944 579804 206972
rect 569368 206932 569374 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 17218 202824 17224 202836
rect 3108 202796 17224 202824
rect 3108 202784 3114 202796
rect 17218 202784 17224 202796
rect 17276 202784 17282 202836
rect 573358 193128 573364 193180
rect 573416 193168 573422 193180
rect 580166 193168 580172 193180
rect 573416 193140 580172 193168
rect 573416 193128 573422 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 14458 189020 14464 189032
rect 3568 188992 14464 189020
rect 3568 188980 3574 188992
rect 14458 188980 14464 188992
rect 14516 188980 14522 189032
rect 566550 166948 566556 167000
rect 566608 166988 566614 167000
rect 580166 166988 580172 167000
rect 566608 166960 580172 166988
rect 566608 166948 566614 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 25590 164200 25596 164212
rect 3292 164172 25596 164200
rect 3292 164160 3298 164172
rect 25590 164160 25596 164172
rect 25648 164160 25654 164212
rect 574738 153144 574744 153196
rect 574796 153184 574802 153196
rect 580166 153184 580172 153196
rect 574796 153156 580172 153184
rect 574796 153144 574802 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3510 150424 3516 150476
rect 3568 150464 3574 150476
rect 4890 150464 4896 150476
rect 3568 150436 4896 150464
rect 3568 150424 3574 150436
rect 4890 150424 4896 150436
rect 4948 150424 4954 150476
rect 569218 139340 569224 139392
rect 569276 139380 569282 139392
rect 580166 139380 580172 139392
rect 569276 139352 580172 139380
rect 569276 139340 569282 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3418 137912 3424 137964
rect 3476 137952 3482 137964
rect 22738 137952 22744 137964
rect 3476 137924 22744 137952
rect 3476 137912 3482 137924
rect 22738 137912 22744 137924
rect 22796 137912 22802 137964
rect 565078 126896 565084 126948
rect 565136 126936 565142 126948
rect 580166 126936 580172 126948
rect 565136 126908 580172 126936
rect 565136 126896 565142 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 558178 113092 558184 113144
rect 558236 113132 558242 113144
rect 579798 113132 579804 113144
rect 558236 113104 579804 113132
rect 558236 113092 558242 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 29730 111772 29736 111784
rect 3200 111744 29736 111772
rect 3200 111732 3206 111744
rect 29730 111732 29736 111744
rect 29788 111732 29794 111784
rect 566458 100648 566464 100700
rect 566516 100688 566522 100700
rect 580166 100688 580172 100700
rect 566516 100660 580172 100688
rect 566516 100648 566522 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 562318 86912 562324 86964
rect 562376 86952 562382 86964
rect 580166 86952 580172 86964
rect 562376 86924 580172 86952
rect 562376 86912 562382 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 25498 85524 25504 85536
rect 3200 85496 25504 85524
rect 3200 85484 3206 85496
rect 25498 85484 25504 85496
rect 25556 85484 25562 85536
rect 576118 73108 576124 73160
rect 576176 73148 576182 73160
rect 580166 73148 580172 73160
rect 576176 73120 580172 73148
rect 576176 73108 576182 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3418 71612 3424 71664
rect 3476 71652 3482 71664
rect 7558 71652 7564 71664
rect 3476 71624 7564 71652
rect 3476 71612 3482 71624
rect 7558 71612 7564 71624
rect 7616 71612 7622 71664
rect 554038 60664 554044 60716
rect 554096 60704 554102 60716
rect 580166 60704 580172 60716
rect 554096 60676 580172 60704
rect 554096 60664 554102 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 2774 58624 2780 58676
rect 2832 58664 2838 58676
rect 4798 58664 4804 58676
rect 2832 58636 4804 58664
rect 2832 58624 2838 58636
rect 4798 58624 4804 58636
rect 4856 58624 4862 58676
rect 560938 46860 560944 46912
rect 560996 46900 561002 46912
rect 580166 46900 580172 46912
rect 560996 46872 580172 46900
rect 560996 46860 561002 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 29638 45540 29644 45552
rect 3476 45512 29644 45540
rect 3476 45500 3482 45512
rect 29638 45500 29644 45512
rect 29696 45500 29702 45552
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 11698 33096 11704 33108
rect 3200 33068 11704 33096
rect 3200 33056 3206 33068
rect 11698 33056 11704 33068
rect 11756 33056 11762 33108
rect 556798 33056 556804 33108
rect 556856 33096 556862 33108
rect 580166 33096 580172 33108
rect 556856 33068 580172 33096
rect 556856 33056 556862 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 20622 30268 20628 30320
rect 20680 30308 20686 30320
rect 50338 30308 50344 30320
rect 20680 30280 50344 30308
rect 20680 30268 20686 30280
rect 50338 30268 50344 30280
rect 50396 30268 50402 30320
rect 50982 30268 50988 30320
rect 51040 30308 51046 30320
rect 76742 30308 76748 30320
rect 51040 30280 76748 30308
rect 51040 30268 51046 30280
rect 76742 30268 76748 30280
rect 76800 30268 76806 30320
rect 78582 30268 78588 30320
rect 78640 30308 78646 30320
rect 101030 30308 101036 30320
rect 78640 30280 101036 30308
rect 78640 30268 78646 30280
rect 101030 30268 101036 30280
rect 101088 30268 101094 30320
rect 101950 30268 101956 30320
rect 102008 30308 102014 30320
rect 122098 30308 122104 30320
rect 102008 30280 122104 30308
rect 102008 30268 102014 30280
rect 122098 30268 122104 30280
rect 122156 30268 122162 30320
rect 128262 30268 128268 30320
rect 128320 30308 128326 30320
rect 145282 30308 145288 30320
rect 128320 30280 145288 30308
rect 128320 30268 128326 30280
rect 145282 30268 145288 30280
rect 145340 30268 145346 30320
rect 146202 30268 146208 30320
rect 146260 30308 146266 30320
rect 162210 30308 162216 30320
rect 146260 30280 162216 30308
rect 146260 30268 146266 30280
rect 162210 30268 162216 30280
rect 162268 30268 162274 30320
rect 168282 30268 168288 30320
rect 168340 30308 168346 30320
rect 181162 30308 181168 30320
rect 168340 30280 181168 30308
rect 168340 30268 168346 30280
rect 181162 30268 181168 30280
rect 181220 30268 181226 30320
rect 183462 30268 183468 30320
rect 183520 30308 183526 30320
rect 194870 30308 194876 30320
rect 183520 30280 194876 30308
rect 183520 30268 183526 30280
rect 194870 30268 194876 30280
rect 194928 30268 194934 30320
rect 200022 30268 200028 30320
rect 200080 30308 200086 30320
rect 209682 30308 209688 30320
rect 200080 30280 209688 30308
rect 200080 30268 200086 30280
rect 209682 30268 209688 30280
rect 209740 30268 209746 30320
rect 224862 30268 224868 30320
rect 224920 30308 224926 30320
rect 231762 30308 231768 30320
rect 224920 30280 231768 30308
rect 224920 30268 224926 30280
rect 231762 30268 231768 30280
rect 231820 30268 231826 30320
rect 244090 30268 244096 30320
rect 244148 30308 244154 30320
rect 248690 30308 248696 30320
rect 244148 30280 248696 30308
rect 244148 30268 244154 30280
rect 248690 30268 248696 30280
rect 248748 30268 248754 30320
rect 255222 30268 255228 30320
rect 255280 30308 255286 30320
rect 259178 30308 259184 30320
rect 255280 30280 259184 30308
rect 255280 30268 255286 30280
rect 259178 30268 259184 30280
rect 259236 30268 259242 30320
rect 277302 30268 277308 30320
rect 277360 30308 277366 30320
rect 278222 30308 278228 30320
rect 277360 30280 278228 30308
rect 277360 30268 277366 30280
rect 278222 30268 278228 30280
rect 278280 30268 278286 30320
rect 286962 30268 286968 30320
rect 287020 30308 287026 30320
rect 287698 30308 287704 30320
rect 287020 30280 287704 30308
rect 287020 30268 287026 30280
rect 287698 30268 287704 30280
rect 287756 30268 287762 30320
rect 315114 30268 315120 30320
rect 315172 30308 315178 30320
rect 316218 30308 316224 30320
rect 315172 30280 316224 30308
rect 315172 30268 315178 30280
rect 316218 30268 316224 30280
rect 316276 30268 316282 30320
rect 16482 30200 16488 30252
rect 16540 30240 16546 30252
rect 40954 30240 40960 30252
rect 16540 30212 40960 30240
rect 16540 30200 16546 30212
rect 40954 30200 40960 30212
rect 41012 30200 41018 30252
rect 41049 30243 41107 30249
rect 41049 30209 41061 30243
rect 41095 30240 41107 30243
rect 48222 30240 48228 30252
rect 41095 30212 48228 30240
rect 41095 30209 41107 30212
rect 41049 30203 41107 30209
rect 48222 30200 48228 30212
rect 48280 30200 48286 30252
rect 50065 30243 50123 30249
rect 50065 30209 50077 30243
rect 50111 30240 50123 30243
rect 54570 30240 54576 30252
rect 50111 30212 54576 30240
rect 50111 30209 50123 30212
rect 50065 30203 50123 30209
rect 54570 30200 54576 30212
rect 54628 30200 54634 30252
rect 56502 30200 56508 30252
rect 56560 30240 56566 30252
rect 81986 30240 81992 30252
rect 56560 30212 81992 30240
rect 56560 30200 56566 30212
rect 81986 30200 81992 30212
rect 82044 30200 82050 30252
rect 86862 30200 86868 30252
rect 86920 30240 86926 30252
rect 109402 30240 109408 30252
rect 86920 30212 109408 30240
rect 86920 30200 86926 30212
rect 109402 30200 109408 30212
rect 109460 30200 109466 30252
rect 111610 30200 111616 30252
rect 111668 30240 111674 30252
rect 130562 30240 130568 30252
rect 111668 30212 130568 30240
rect 111668 30200 111674 30212
rect 130562 30200 130568 30212
rect 130620 30200 130626 30252
rect 155770 30200 155776 30252
rect 155828 30240 155834 30252
rect 170582 30240 170588 30252
rect 155828 30212 170588 30240
rect 155828 30200 155834 30212
rect 170582 30200 170588 30212
rect 170640 30200 170646 30252
rect 179322 30200 179328 30252
rect 179380 30240 179386 30252
rect 191742 30240 191748 30252
rect 179380 30212 191748 30240
rect 179380 30200 179386 30212
rect 191742 30200 191748 30212
rect 191800 30200 191806 30252
rect 193122 30200 193128 30252
rect 193180 30240 193186 30252
rect 203334 30240 203340 30252
rect 193180 30212 203340 30240
rect 193180 30200 193186 30212
rect 203334 30200 203340 30212
rect 203392 30200 203398 30252
rect 205542 30200 205548 30252
rect 205600 30240 205606 30252
rect 214926 30240 214932 30252
rect 205600 30212 214932 30240
rect 205600 30200 205606 30212
rect 214926 30200 214932 30212
rect 214984 30200 214990 30252
rect 223482 30200 223488 30252
rect 223540 30240 223546 30252
rect 230750 30240 230756 30252
rect 223540 30212 230756 30240
rect 223540 30200 223546 30212
rect 230750 30200 230756 30212
rect 230808 30200 230814 30252
rect 253842 30200 253848 30252
rect 253900 30240 253906 30252
rect 258166 30240 258172 30252
rect 253900 30212 258172 30240
rect 253900 30200 253906 30212
rect 258166 30200 258172 30212
rect 258224 30200 258230 30252
rect 470134 30200 470140 30252
rect 470192 30240 470198 30252
rect 471330 30240 471336 30252
rect 470192 30212 471336 30240
rect 470192 30200 470198 30212
rect 471330 30200 471336 30212
rect 471388 30200 471394 30252
rect 23382 30132 23388 30184
rect 23440 30172 23446 30184
rect 52454 30172 52460 30184
rect 23440 30144 52460 30172
rect 23440 30132 23446 30144
rect 52454 30132 52460 30144
rect 52512 30132 52518 30184
rect 53650 30132 53656 30184
rect 53708 30172 53714 30184
rect 78858 30172 78864 30184
rect 53708 30144 78864 30172
rect 53708 30132 53714 30144
rect 78858 30132 78864 30144
rect 78916 30132 78922 30184
rect 88242 30132 88248 30184
rect 88300 30172 88306 30184
rect 110506 30172 110512 30184
rect 88300 30144 110512 30172
rect 88300 30132 88306 30144
rect 110506 30132 110512 30144
rect 110564 30132 110570 30184
rect 113082 30132 113088 30184
rect 113140 30172 113146 30184
rect 132678 30172 132684 30184
rect 113140 30144 132684 30172
rect 113140 30132 113146 30144
rect 132678 30132 132684 30144
rect 132736 30132 132742 30184
rect 133782 30132 133788 30184
rect 133840 30172 133846 30184
rect 150618 30172 150624 30184
rect 133840 30144 150624 30172
rect 133840 30132 133846 30144
rect 150618 30132 150624 30144
rect 150676 30132 150682 30184
rect 158622 30132 158628 30184
rect 158680 30172 158686 30184
rect 172698 30172 172704 30184
rect 158680 30144 172704 30172
rect 158680 30132 158686 30144
rect 172698 30132 172704 30144
rect 172756 30132 172762 30184
rect 175182 30132 175188 30184
rect 175240 30172 175246 30184
rect 187510 30172 187516 30184
rect 175240 30144 187516 30172
rect 175240 30132 175246 30144
rect 187510 30132 187516 30144
rect 187568 30132 187574 30184
rect 190362 30132 190368 30184
rect 190420 30172 190426 30184
rect 201218 30172 201224 30184
rect 190420 30144 201224 30172
rect 190420 30132 190426 30144
rect 201218 30132 201224 30144
rect 201276 30132 201282 30184
rect 202782 30132 202788 30184
rect 202840 30172 202846 30184
rect 211706 30172 211712 30184
rect 202840 30144 211712 30172
rect 202840 30132 202846 30144
rect 211706 30132 211712 30144
rect 211764 30132 211770 30184
rect 216582 30132 216588 30184
rect 216640 30172 216646 30184
rect 224402 30172 224408 30184
rect 216640 30144 224408 30172
rect 216640 30132 216646 30144
rect 224402 30132 224408 30144
rect 224460 30132 224466 30184
rect 244182 30132 244188 30184
rect 244240 30172 244246 30184
rect 249702 30172 249708 30184
rect 244240 30144 249708 30172
rect 244240 30132 244246 30144
rect 249702 30132 249708 30144
rect 249760 30132 249766 30184
rect 10962 30064 10968 30116
rect 11020 30104 11026 30116
rect 40770 30104 40776 30116
rect 11020 30076 40776 30104
rect 11020 30064 11026 30076
rect 40770 30064 40776 30076
rect 40828 30064 40834 30116
rect 66162 30104 66168 30116
rect 41064 30076 66168 30104
rect 31021 30039 31079 30045
rect 31021 30005 31033 30039
rect 31067 30036 31079 30039
rect 36630 30036 36636 30048
rect 31067 30008 36636 30036
rect 31067 30005 31079 30008
rect 31021 29999 31079 30005
rect 36630 29996 36636 30008
rect 36688 29996 36694 30048
rect 38562 29996 38568 30048
rect 38620 30036 38626 30048
rect 41064 30036 41092 30076
rect 66162 30064 66168 30076
rect 66220 30064 66226 30116
rect 67542 30064 67548 30116
rect 67600 30104 67606 30116
rect 91554 30104 91560 30116
rect 67600 30076 91560 30104
rect 67600 30064 67606 30076
rect 91554 30064 91560 30076
rect 91612 30064 91618 30116
rect 92382 30064 92388 30116
rect 92440 30104 92446 30116
rect 113634 30104 113640 30116
rect 92440 30076 113640 30104
rect 92440 30064 92446 30076
rect 113634 30064 113640 30076
rect 113692 30064 113698 30116
rect 124122 30064 124128 30116
rect 124180 30104 124186 30116
rect 142154 30104 142160 30116
rect 124180 30076 142160 30104
rect 124180 30064 124186 30076
rect 142154 30064 142160 30076
rect 142212 30064 142218 30116
rect 147582 30064 147588 30116
rect 147640 30104 147646 30116
rect 163222 30104 163228 30116
rect 147640 30076 163228 30104
rect 147640 30064 147646 30076
rect 163222 30064 163228 30076
rect 163280 30064 163286 30116
rect 166902 30064 166908 30116
rect 166960 30104 166966 30116
rect 180150 30104 180156 30116
rect 166960 30076 180156 30104
rect 166960 30064 166966 30076
rect 180150 30064 180156 30076
rect 180208 30064 180214 30116
rect 182082 30064 182088 30116
rect 182140 30104 182146 30116
rect 193858 30104 193864 30116
rect 182140 30076 193864 30104
rect 182140 30064 182146 30076
rect 193858 30064 193864 30076
rect 193916 30064 193922 30116
rect 195882 30064 195888 30116
rect 195940 30104 195946 30116
rect 206462 30104 206468 30116
rect 195940 30076 206468 30104
rect 195940 30064 195946 30076
rect 206462 30064 206468 30076
rect 206520 30064 206526 30116
rect 206922 30064 206928 30116
rect 206980 30104 206986 30116
rect 215938 30104 215944 30116
rect 206980 30076 215944 30104
rect 206980 30064 206986 30076
rect 215938 30064 215944 30076
rect 215996 30064 216002 30116
rect 217962 30064 217968 30116
rect 218020 30104 218026 30116
rect 225506 30104 225512 30116
rect 218020 30076 225512 30104
rect 218020 30064 218026 30076
rect 225506 30064 225512 30076
rect 225564 30064 225570 30116
rect 226242 30064 226248 30116
rect 226300 30104 226306 30116
rect 232866 30104 232872 30116
rect 226300 30076 232872 30104
rect 226300 30064 226306 30076
rect 232866 30064 232872 30076
rect 232924 30064 232930 30116
rect 233142 30064 233148 30116
rect 233200 30104 233206 30116
rect 239214 30104 239220 30116
rect 233200 30076 239220 30104
rect 233200 30064 233206 30076
rect 239214 30064 239220 30076
rect 239272 30064 239278 30116
rect 38620 30008 41092 30036
rect 41141 30039 41199 30045
rect 38620 29996 38626 30008
rect 41141 30005 41153 30039
rect 41187 30036 41199 30039
rect 63034 30036 63040 30048
rect 41187 30008 63040 30036
rect 41187 30005 41199 30008
rect 41141 29999 41199 30005
rect 63034 29996 63040 30008
rect 63092 29996 63098 30048
rect 63402 29996 63408 30048
rect 63460 30036 63466 30048
rect 88334 30036 88340 30048
rect 63460 30008 88340 30036
rect 63460 29996 63466 30008
rect 88334 29996 88340 30008
rect 88392 29996 88398 30048
rect 89622 29996 89628 30048
rect 89680 30036 89686 30048
rect 111518 30036 111524 30048
rect 89680 30008 111524 30036
rect 89680 29996 89686 30008
rect 111518 29996 111524 30008
rect 111576 29996 111582 30048
rect 111702 29996 111708 30048
rect 111760 30036 111766 30048
rect 131574 30036 131580 30048
rect 111760 30008 131580 30036
rect 111760 29996 111766 30008
rect 131574 29996 131580 30008
rect 131632 29996 131638 30048
rect 132402 29996 132408 30048
rect 132460 30036 132466 30048
rect 149514 30036 149520 30048
rect 132460 30008 149520 30036
rect 132460 29996 132466 30008
rect 149514 29996 149520 30008
rect 149572 29996 149578 30048
rect 154482 29996 154488 30048
rect 154540 30036 154546 30048
rect 169570 30036 169576 30048
rect 154540 30008 169576 30036
rect 154540 29996 154546 30008
rect 169570 29996 169576 30008
rect 169628 29996 169634 30048
rect 173710 29996 173716 30048
rect 173768 30036 173774 30048
rect 186406 30036 186412 30048
rect 173768 30008 186412 30036
rect 173768 29996 173774 30008
rect 186406 29996 186412 30008
rect 186464 29996 186470 30048
rect 197262 29996 197268 30048
rect 197320 30036 197326 30048
rect 207566 30036 207572 30048
rect 197320 30008 207572 30036
rect 197320 29996 197326 30008
rect 207566 29996 207572 30008
rect 207624 29996 207630 30048
rect 13722 29928 13728 29980
rect 13780 29968 13786 29980
rect 40037 29971 40095 29977
rect 13780 29940 39988 29968
rect 13780 29928 13786 29940
rect 15102 29860 15108 29912
rect 15160 29900 15166 29912
rect 39853 29903 39911 29909
rect 39853 29900 39865 29903
rect 15160 29872 39865 29900
rect 15160 29860 15166 29872
rect 39853 29869 39865 29872
rect 39899 29869 39911 29903
rect 39960 29900 39988 29940
rect 40037 29937 40049 29971
rect 40083 29968 40095 29971
rect 40865 29971 40923 29977
rect 40865 29968 40877 29971
rect 40083 29940 40877 29968
rect 40083 29937 40095 29940
rect 40037 29931 40095 29937
rect 40865 29937 40877 29940
rect 40911 29937 40923 29971
rect 40865 29931 40923 29937
rect 40954 29928 40960 29980
rect 41012 29968 41018 29980
rect 46198 29968 46204 29980
rect 41012 29940 46204 29968
rect 41012 29928 41018 29940
rect 46198 29928 46204 29940
rect 46256 29928 46262 29980
rect 46753 29971 46811 29977
rect 46753 29937 46765 29971
rect 46799 29968 46811 29971
rect 50065 29971 50123 29977
rect 50065 29968 50077 29971
rect 46799 29940 50077 29968
rect 46799 29937 46811 29940
rect 46753 29931 46811 29937
rect 50065 29937 50077 29940
rect 50111 29937 50123 29971
rect 50065 29931 50123 29937
rect 50249 29971 50307 29977
rect 50249 29937 50261 29971
rect 50295 29968 50307 29971
rect 71498 29968 71504 29980
rect 50295 29940 71504 29968
rect 50295 29937 50307 29940
rect 50249 29931 50307 29937
rect 71498 29928 71504 29940
rect 71556 29928 71562 29980
rect 82722 29928 82728 29980
rect 82780 29968 82786 29980
rect 105262 29968 105268 29980
rect 82780 29940 105268 29968
rect 82780 29928 82786 29940
rect 105262 29928 105268 29940
rect 105320 29928 105326 29980
rect 108942 29928 108948 29980
rect 109000 29968 109006 29980
rect 128446 29968 128452 29980
rect 109000 29940 128452 29968
rect 109000 29928 109006 29940
rect 128446 29928 128452 29940
rect 128504 29928 128510 29980
rect 131022 29928 131028 29980
rect 131080 29968 131086 29980
rect 148502 29968 148508 29980
rect 131080 29940 148508 29968
rect 131080 29928 131086 29940
rect 148502 29928 148508 29940
rect 148560 29928 148566 29980
rect 148962 29928 148968 29980
rect 149020 29968 149026 29980
rect 164326 29968 164332 29980
rect 149020 29940 164332 29968
rect 149020 29928 149026 29940
rect 164326 29928 164332 29940
rect 164384 29928 164390 29980
rect 171042 29928 171048 29980
rect 171100 29968 171106 29980
rect 184290 29968 184296 29980
rect 171100 29940 184296 29968
rect 171100 29928 171106 29940
rect 184290 29928 184296 29940
rect 184348 29928 184354 29980
rect 188982 29928 188988 29980
rect 189040 29968 189046 29980
rect 200114 29968 200120 29980
rect 189040 29940 200120 29968
rect 189040 29928 189046 29940
rect 200114 29928 200120 29940
rect 200172 29928 200178 29980
rect 204162 29928 204168 29980
rect 204220 29968 204226 29980
rect 213822 29968 213828 29980
rect 204220 29940 213828 29968
rect 204220 29928 204226 29940
rect 213822 29928 213828 29940
rect 213880 29928 213886 29980
rect 215202 29928 215208 29980
rect 215260 29968 215266 29980
rect 223390 29968 223396 29980
rect 215260 29940 223396 29968
rect 215260 29928 215266 29940
rect 223390 29928 223396 29940
rect 223448 29928 223454 29980
rect 227438 29928 227444 29980
rect 227496 29968 227502 29980
rect 233878 29968 233884 29980
rect 227496 29940 233884 29968
rect 227496 29928 227502 29940
rect 233878 29928 233884 29940
rect 233936 29928 233942 29980
rect 523954 29928 523960 29980
rect 524012 29968 524018 29980
rect 529290 29968 529296 29980
rect 524012 29940 529296 29968
rect 524012 29928 524018 29940
rect 529290 29928 529296 29940
rect 529348 29928 529354 29980
rect 44082 29900 44088 29912
rect 39960 29872 44088 29900
rect 39853 29863 39911 29869
rect 44082 29860 44088 29872
rect 44140 29860 44146 29912
rect 45462 29860 45468 29912
rect 45520 29900 45526 29912
rect 72510 29900 72516 29912
rect 45520 29872 72516 29900
rect 45520 29860 45526 29872
rect 72510 29860 72516 29872
rect 72568 29860 72574 29912
rect 75822 29860 75828 29912
rect 75880 29900 75886 29912
rect 98914 29900 98920 29912
rect 75880 29872 98920 29900
rect 75880 29860 75886 29872
rect 98914 29860 98920 29872
rect 98972 29860 98978 29912
rect 100662 29860 100668 29912
rect 100720 29900 100726 29912
rect 121086 29900 121092 29912
rect 100720 29872 121092 29900
rect 100720 29860 100726 29872
rect 121086 29860 121092 29872
rect 121144 29860 121150 29912
rect 122742 29860 122748 29912
rect 122800 29900 122806 29912
rect 141050 29900 141056 29912
rect 122800 29872 141056 29900
rect 122800 29860 122806 29872
rect 141050 29860 141056 29872
rect 141108 29860 141114 29912
rect 143442 29860 143448 29912
rect 143500 29900 143506 29912
rect 158990 29900 158996 29912
rect 143500 29872 158996 29900
rect 143500 29860 143506 29872
rect 158990 29860 158996 29872
rect 159048 29860 159054 29912
rect 164142 29860 164148 29912
rect 164200 29900 164206 29912
rect 178034 29900 178040 29912
rect 164200 29872 178040 29900
rect 164200 29860 164206 29872
rect 178034 29860 178040 29872
rect 178092 29860 178098 29912
rect 180702 29860 180708 29912
rect 180760 29900 180766 29912
rect 192754 29900 192760 29912
rect 180760 29872 192760 29900
rect 180760 29860 180766 29872
rect 192754 29860 192760 29872
rect 192812 29860 192818 29912
rect 194502 29860 194508 29912
rect 194560 29900 194566 29912
rect 205450 29900 205456 29912
rect 194560 29872 205456 29900
rect 194560 29860 194566 29872
rect 205450 29860 205456 29872
rect 205508 29860 205514 29912
rect 209682 29860 209688 29912
rect 209740 29900 209746 29912
rect 218054 29900 218060 29912
rect 209740 29872 218060 29900
rect 209740 29860 209746 29872
rect 218054 29860 218060 29872
rect 218112 29860 218118 29912
rect 219342 29860 219348 29912
rect 219400 29900 219406 29912
rect 227530 29900 227536 29912
rect 219400 29872 227536 29900
rect 219400 29860 219406 29872
rect 227530 29860 227536 29872
rect 227588 29860 227594 29912
rect 227622 29860 227628 29912
rect 227680 29900 227686 29912
rect 234982 29900 234988 29912
rect 227680 29872 234988 29900
rect 227680 29860 227686 29872
rect 234982 29860 234988 29872
rect 235040 29860 235046 29912
rect 248322 29860 248328 29912
rect 248380 29900 248386 29912
rect 252922 29900 252928 29912
rect 248380 29872 252928 29900
rect 248380 29860 248386 29872
rect 252922 29860 252928 29872
rect 252980 29860 252986 29912
rect 257982 29860 257988 29912
rect 258040 29900 258046 29912
rect 261294 29900 261300 29912
rect 258040 29872 261300 29900
rect 258040 29860 258046 29872
rect 261294 29860 261300 29872
rect 261352 29860 261358 29912
rect 546126 29860 546132 29912
rect 546184 29900 546190 29912
rect 556798 29900 556804 29912
rect 546184 29872 556804 29900
rect 546184 29860 546190 29872
rect 556798 29860 556804 29872
rect 556856 29860 556862 29912
rect 12250 29792 12256 29844
rect 12308 29832 12314 29844
rect 41966 29832 41972 29844
rect 12308 29804 41972 29832
rect 12308 29792 12314 29804
rect 41966 29792 41972 29804
rect 42024 29792 42030 29844
rect 45370 29792 45376 29844
rect 45428 29832 45434 29844
rect 50249 29835 50307 29841
rect 50249 29832 50261 29835
rect 45428 29804 50261 29832
rect 45428 29792 45434 29804
rect 50249 29801 50261 29804
rect 50295 29801 50307 29835
rect 69382 29832 69388 29844
rect 50249 29795 50307 29801
rect 50356 29804 69388 29832
rect 6822 29724 6828 29776
rect 6880 29764 6886 29776
rect 37734 29764 37740 29776
rect 6880 29736 37740 29764
rect 6880 29724 6886 29736
rect 37734 29724 37740 29736
rect 37792 29724 37798 29776
rect 39853 29767 39911 29773
rect 39853 29733 39865 29767
rect 39899 29764 39911 29767
rect 45094 29764 45100 29776
rect 39899 29736 45100 29764
rect 39899 29733 39911 29736
rect 39853 29727 39911 29733
rect 45094 29724 45100 29736
rect 45152 29724 45158 29776
rect 3970 29656 3976 29708
rect 4028 29696 4034 29708
rect 35618 29696 35624 29708
rect 4028 29668 35624 29696
rect 4028 29656 4034 29668
rect 35618 29656 35624 29668
rect 35676 29656 35682 29708
rect 35802 29656 35808 29708
rect 35860 29696 35866 29708
rect 41141 29699 41199 29705
rect 41141 29696 41153 29699
rect 35860 29668 41153 29696
rect 35860 29656 35866 29668
rect 41141 29665 41153 29668
rect 41187 29665 41199 29699
rect 41141 29659 41199 29665
rect 42702 29656 42708 29708
rect 42760 29696 42766 29708
rect 50356 29696 50384 29804
rect 69382 29792 69388 29804
rect 69440 29792 69446 29844
rect 70302 29792 70308 29844
rect 70360 29832 70366 29844
rect 94682 29832 94688 29844
rect 70360 29804 94688 29832
rect 70360 29792 70366 29804
rect 94682 29792 94688 29804
rect 94740 29792 94746 29844
rect 96522 29792 96528 29844
rect 96580 29832 96586 29844
rect 117866 29832 117872 29844
rect 96580 29804 117872 29832
rect 96580 29792 96586 29804
rect 117866 29792 117872 29804
rect 117924 29792 117930 29844
rect 118602 29792 118608 29844
rect 118660 29832 118666 29844
rect 136818 29832 136824 29844
rect 118660 29804 136824 29832
rect 118660 29792 118666 29804
rect 136818 29792 136824 29804
rect 136876 29792 136882 29844
rect 137922 29792 137928 29844
rect 137980 29832 137986 29844
rect 154758 29832 154764 29844
rect 137980 29804 154764 29832
rect 137980 29792 137986 29804
rect 154758 29792 154764 29804
rect 154816 29792 154822 29844
rect 157242 29792 157248 29844
rect 157300 29832 157306 29844
rect 171686 29832 171692 29844
rect 157300 29804 171692 29832
rect 157300 29792 157306 29804
rect 171686 29792 171692 29804
rect 171744 29792 171750 29844
rect 172422 29792 172428 29844
rect 172480 29832 172486 29844
rect 185394 29832 185400 29844
rect 172480 29804 185400 29832
rect 172480 29792 172486 29804
rect 185394 29792 185400 29804
rect 185452 29792 185458 29844
rect 187602 29792 187608 29844
rect 187660 29832 187666 29844
rect 199102 29832 199108 29844
rect 187660 29804 199108 29832
rect 187660 29792 187666 29804
rect 199102 29792 199108 29804
rect 199160 29792 199166 29844
rect 201402 29792 201408 29844
rect 201460 29832 201466 29844
rect 210694 29832 210700 29844
rect 201460 29804 210700 29832
rect 201460 29792 201466 29804
rect 210694 29792 210700 29804
rect 210752 29792 210758 29844
rect 212442 29792 212448 29844
rect 212500 29832 212506 29844
rect 221274 29832 221280 29844
rect 212500 29804 221280 29832
rect 212500 29792 212506 29804
rect 221274 29792 221280 29804
rect 221332 29792 221338 29844
rect 222102 29792 222108 29844
rect 222160 29832 222166 29844
rect 229646 29832 229652 29844
rect 222160 29804 229652 29832
rect 222160 29792 222166 29804
rect 229646 29792 229652 29804
rect 229704 29792 229710 29844
rect 530302 29792 530308 29844
rect 530360 29832 530366 29844
rect 557534 29832 557540 29844
rect 530360 29804 557540 29832
rect 530360 29792 530366 29804
rect 557534 29792 557540 29804
rect 557592 29792 557598 29844
rect 50433 29767 50491 29773
rect 50433 29733 50445 29767
rect 50479 29764 50491 29767
rect 67266 29764 67272 29776
rect 50479 29736 67272 29764
rect 50479 29733 50491 29736
rect 50433 29727 50491 29733
rect 67266 29724 67272 29736
rect 67324 29724 67330 29776
rect 68922 29724 68928 29776
rect 68980 29764 68986 29776
rect 92566 29764 92572 29776
rect 68980 29736 92572 29764
rect 68980 29724 68986 29736
rect 92566 29724 92572 29736
rect 92624 29724 92630 29776
rect 93762 29724 93768 29776
rect 93820 29764 93826 29776
rect 114738 29764 114744 29776
rect 93820 29736 114744 29764
rect 93820 29724 93826 29736
rect 114738 29724 114744 29736
rect 114796 29724 114802 29776
rect 119890 29724 119896 29776
rect 119948 29764 119954 29776
rect 138934 29764 138940 29776
rect 119948 29736 138940 29764
rect 119948 29724 119954 29736
rect 138934 29724 138940 29736
rect 138992 29724 138998 29776
rect 144730 29724 144736 29776
rect 144788 29764 144794 29776
rect 161106 29764 161112 29776
rect 144788 29736 161112 29764
rect 144788 29724 144794 29736
rect 161106 29724 161112 29736
rect 161164 29724 161170 29776
rect 162762 29724 162768 29776
rect 162820 29764 162826 29776
rect 176930 29764 176936 29776
rect 162820 29736 176936 29764
rect 162820 29724 162826 29736
rect 176930 29724 176936 29736
rect 176988 29724 176994 29776
rect 177850 29724 177856 29776
rect 177908 29764 177914 29776
rect 189626 29764 189632 29776
rect 177908 29736 189632 29764
rect 177908 29724 177914 29736
rect 189626 29724 189632 29736
rect 189684 29724 189690 29776
rect 198642 29724 198648 29776
rect 198700 29764 198706 29776
rect 208578 29764 208584 29776
rect 198700 29736 208584 29764
rect 198700 29724 198706 29736
rect 208578 29724 208584 29736
rect 208636 29724 208642 29776
rect 211062 29724 211068 29776
rect 211120 29764 211126 29776
rect 220170 29764 220176 29776
rect 211120 29736 220176 29764
rect 211120 29724 211126 29736
rect 220170 29724 220176 29736
rect 220228 29724 220234 29776
rect 238662 29724 238668 29776
rect 238720 29764 238726 29776
rect 244458 29764 244464 29776
rect 238720 29736 244464 29764
rect 238720 29724 238726 29736
rect 244458 29724 244464 29736
rect 244516 29724 244522 29776
rect 256602 29724 256608 29776
rect 256660 29764 256666 29776
rect 260282 29764 260288 29776
rect 256660 29736 260288 29764
rect 256660 29724 256666 29736
rect 260282 29724 260288 29736
rect 260340 29724 260346 29776
rect 536650 29724 536656 29776
rect 536708 29764 536714 29776
rect 564526 29764 564532 29776
rect 536708 29736 564532 29764
rect 536708 29724 536714 29736
rect 564526 29724 564532 29736
rect 564584 29724 564590 29776
rect 42760 29668 50384 29696
rect 50525 29699 50583 29705
rect 42760 29656 42766 29668
rect 50525 29665 50537 29699
rect 50571 29696 50583 29699
rect 73614 29696 73620 29708
rect 50571 29668 73620 29696
rect 50571 29665 50583 29668
rect 50525 29659 50583 29665
rect 73614 29656 73620 29668
rect 73672 29656 73678 29708
rect 78490 29656 78496 29708
rect 78548 29696 78554 29708
rect 102042 29696 102048 29708
rect 78548 29668 102048 29696
rect 78548 29656 78554 29668
rect 102042 29656 102048 29668
rect 102100 29656 102106 29708
rect 105265 29699 105323 29705
rect 105265 29665 105277 29699
rect 105311 29696 105323 29699
rect 107473 29699 107531 29705
rect 107473 29696 107485 29699
rect 105311 29668 107485 29696
rect 105311 29665 105323 29668
rect 105265 29659 105323 29665
rect 107473 29665 107485 29668
rect 107519 29665 107531 29699
rect 107473 29659 107531 29665
rect 107562 29656 107568 29708
rect 107620 29696 107626 29708
rect 127342 29696 127348 29708
rect 107620 29668 127348 29696
rect 107620 29656 107626 29668
rect 127342 29656 127348 29668
rect 127400 29656 127406 29708
rect 136450 29656 136456 29708
rect 136508 29696 136514 29708
rect 153746 29696 153752 29708
rect 136508 29668 153752 29696
rect 136508 29656 136514 29668
rect 153746 29656 153752 29668
rect 153804 29656 153810 29708
rect 161290 29656 161296 29708
rect 161348 29696 161354 29708
rect 175918 29696 175924 29708
rect 161348 29668 175924 29696
rect 161348 29656 161354 29668
rect 175918 29656 175924 29668
rect 175976 29656 175982 29708
rect 177942 29656 177948 29708
rect 178000 29696 178006 29708
rect 190638 29696 190644 29708
rect 178000 29668 190644 29696
rect 178000 29656 178006 29668
rect 190638 29656 190644 29668
rect 190696 29656 190702 29708
rect 194410 29656 194416 29708
rect 194468 29696 194474 29708
rect 204346 29696 204352 29708
rect 194468 29668 204352 29696
rect 194468 29656 194474 29668
rect 204346 29656 204352 29668
rect 204404 29656 204410 29708
rect 208302 29656 208308 29708
rect 208360 29696 208366 29708
rect 217042 29696 217048 29708
rect 208360 29668 217048 29696
rect 208360 29656 208366 29668
rect 217042 29656 217048 29668
rect 217100 29656 217106 29708
rect 219250 29656 219256 29708
rect 219308 29696 219314 29708
rect 226518 29696 226524 29708
rect 219308 29668 226524 29696
rect 219308 29656 219314 29668
rect 226518 29656 226524 29668
rect 226576 29656 226582 29708
rect 229002 29656 229008 29708
rect 229060 29696 229066 29708
rect 235994 29696 236000 29708
rect 229060 29668 236000 29696
rect 229060 29656 229066 29668
rect 235994 29656 236000 29668
rect 236052 29656 236058 29708
rect 237282 29656 237288 29708
rect 237340 29696 237346 29708
rect 243354 29696 243360 29708
rect 237340 29668 243360 29696
rect 237340 29656 237346 29668
rect 243354 29656 243360 29668
rect 243412 29656 243418 29708
rect 246942 29656 246948 29708
rect 247000 29696 247006 29708
rect 251818 29696 251824 29708
rect 247000 29668 251824 29696
rect 247000 29656 247006 29668
rect 251818 29656 251824 29668
rect 251876 29656 251882 29708
rect 508130 29656 508136 29708
rect 508188 29696 508194 29708
rect 511350 29696 511356 29708
rect 508188 29668 511356 29696
rect 508188 29656 508194 29668
rect 511350 29656 511356 29668
rect 511408 29656 511414 29708
rect 514478 29656 514484 29708
rect 514536 29696 514542 29708
rect 525058 29696 525064 29708
rect 514536 29668 525064 29696
rect 514536 29656 514542 29668
rect 525058 29656 525064 29668
rect 525116 29656 525122 29708
rect 539778 29656 539784 29708
rect 539836 29696 539842 29708
rect 568574 29696 568580 29708
rect 539836 29668 568580 29696
rect 539836 29656 539842 29668
rect 568574 29656 568580 29668
rect 568632 29656 568638 29708
rect 5442 29588 5448 29640
rect 5500 29628 5506 29640
rect 31021 29631 31079 29637
rect 31021 29628 31033 29631
rect 5500 29600 31033 29628
rect 5500 29588 5506 29600
rect 31021 29597 31033 29600
rect 31067 29597 31079 29631
rect 31021 29591 31079 29597
rect 33042 29588 33048 29640
rect 33100 29628 33106 29640
rect 40681 29631 40739 29637
rect 40681 29628 40693 29631
rect 33100 29600 40693 29628
rect 33100 29588 33106 29600
rect 40681 29597 40693 29600
rect 40727 29597 40739 29631
rect 40681 29591 40739 29597
rect 44082 29588 44088 29640
rect 44140 29628 44146 29640
rect 70394 29628 70400 29640
rect 44140 29600 70400 29628
rect 44140 29588 44146 29600
rect 70394 29588 70400 29600
rect 70452 29588 70458 29640
rect 71682 29588 71688 29640
rect 71740 29628 71746 29640
rect 95694 29628 95700 29640
rect 71740 29600 95700 29628
rect 71740 29588 71746 29600
rect 95694 29588 95700 29600
rect 95752 29588 95758 29640
rect 100754 29588 100760 29640
rect 100812 29628 100818 29640
rect 103146 29628 103152 29640
rect 100812 29600 103152 29628
rect 100812 29588 100818 29600
rect 103146 29588 103152 29600
rect 103204 29588 103210 29640
rect 103330 29588 103336 29640
rect 103388 29628 103394 29640
rect 124214 29628 124220 29640
rect 103388 29600 124220 29628
rect 103388 29588 103394 29600
rect 124214 29588 124220 29600
rect 124272 29588 124278 29640
rect 128170 29588 128176 29640
rect 128228 29628 128234 29640
rect 146386 29628 146392 29640
rect 128228 29600 146392 29628
rect 128228 29588 128234 29600
rect 146386 29588 146392 29600
rect 146444 29588 146450 29640
rect 153010 29588 153016 29640
rect 153068 29628 153074 29640
rect 168466 29628 168472 29640
rect 153068 29600 168472 29628
rect 153068 29588 153074 29600
rect 168466 29588 168472 29600
rect 168524 29588 168530 29640
rect 169570 29588 169576 29640
rect 169628 29628 169634 29640
rect 182174 29628 182180 29640
rect 169628 29600 182180 29628
rect 169628 29588 169634 29600
rect 182174 29588 182180 29600
rect 182232 29588 182238 29640
rect 186130 29588 186136 29640
rect 186188 29628 186194 29640
rect 197998 29628 198004 29640
rect 186188 29600 198004 29628
rect 186188 29588 186194 29600
rect 197998 29588 198004 29600
rect 198056 29588 198062 29640
rect 202690 29588 202696 29640
rect 202748 29628 202754 29640
rect 212810 29628 212816 29640
rect 202748 29600 212816 29628
rect 202748 29588 202754 29600
rect 212810 29588 212816 29600
rect 212868 29588 212874 29640
rect 213822 29588 213828 29640
rect 213880 29628 213886 29640
rect 222286 29628 222292 29640
rect 213880 29600 222292 29628
rect 213880 29588 213886 29600
rect 222286 29588 222292 29600
rect 222344 29588 222350 29640
rect 235810 29588 235816 29640
rect 235868 29628 235874 29640
rect 242342 29628 242348 29640
rect 235868 29600 242348 29628
rect 235868 29588 235874 29600
rect 242342 29588 242348 29600
rect 242400 29588 242406 29640
rect 498654 29588 498660 29640
rect 498712 29628 498718 29640
rect 520918 29628 520924 29640
rect 498712 29600 520924 29628
rect 498712 29588 498718 29600
rect 520918 29588 520924 29600
rect 520976 29588 520982 29640
rect 572806 29628 572812 29640
rect 547846 29600 572812 29628
rect 20530 29520 20536 29572
rect 20588 29560 20594 29572
rect 49326 29560 49332 29572
rect 20588 29532 49332 29560
rect 20588 29520 20594 29532
rect 49326 29520 49332 29532
rect 49384 29520 49390 29572
rect 49602 29520 49608 29572
rect 49660 29560 49666 29572
rect 75730 29560 75736 29572
rect 49660 29532 75736 29560
rect 49660 29520 49666 29532
rect 75730 29520 75736 29532
rect 75788 29520 75794 29572
rect 81342 29520 81348 29572
rect 81400 29560 81406 29572
rect 104158 29560 104164 29572
rect 81400 29532 104164 29560
rect 81400 29520 81406 29532
rect 104158 29520 104164 29532
rect 104216 29520 104222 29572
rect 104802 29520 104808 29572
rect 104860 29560 104866 29572
rect 125226 29560 125232 29572
rect 104860 29532 125232 29560
rect 104860 29520 104866 29532
rect 125226 29520 125232 29532
rect 125284 29520 125290 29572
rect 125502 29520 125508 29572
rect 125560 29560 125566 29572
rect 143166 29560 143172 29572
rect 125560 29532 143172 29560
rect 125560 29520 125566 29532
rect 143166 29520 143172 29532
rect 143224 29520 143230 29572
rect 144822 29520 144828 29572
rect 144880 29560 144886 29572
rect 160094 29560 160100 29572
rect 144880 29532 160100 29560
rect 144880 29520 144886 29532
rect 160094 29520 160100 29532
rect 160152 29520 160158 29572
rect 165522 29520 165528 29572
rect 165580 29560 165586 29572
rect 179046 29560 179052 29572
rect 165580 29532 179052 29560
rect 165580 29520 165586 29532
rect 179046 29520 179052 29532
rect 179104 29520 179110 29572
rect 186222 29520 186228 29572
rect 186280 29560 186286 29572
rect 196986 29560 196992 29572
rect 186280 29532 196992 29560
rect 186280 29520 186286 29532
rect 196986 29520 196992 29532
rect 197044 29520 197050 29572
rect 235902 29520 235908 29572
rect 235960 29560 235966 29572
rect 241238 29560 241244 29572
rect 235960 29532 241244 29560
rect 235960 29520 235966 29532
rect 241238 29520 241244 29532
rect 241296 29520 241302 29572
rect 542906 29520 542912 29572
rect 542964 29560 542970 29572
rect 547846 29560 547874 29600
rect 572806 29588 572812 29600
rect 572864 29588 572870 29640
rect 542964 29532 547874 29560
rect 542964 29520 542970 29532
rect 28810 29452 28816 29504
rect 28868 29492 28874 29504
rect 57790 29492 57796 29504
rect 28868 29464 57796 29492
rect 28868 29452 28874 29464
rect 57790 29452 57796 29464
rect 57848 29452 57854 29504
rect 57882 29452 57888 29504
rect 57940 29492 57946 29504
rect 83090 29492 83096 29504
rect 57940 29464 83096 29492
rect 57940 29452 57946 29464
rect 83090 29452 83096 29464
rect 83148 29452 83154 29504
rect 86770 29452 86776 29504
rect 86828 29492 86834 29504
rect 108390 29492 108396 29504
rect 86828 29464 108396 29492
rect 86828 29452 86834 29464
rect 108390 29452 108396 29464
rect 108448 29452 108454 29504
rect 112622 29492 112628 29504
rect 108500 29464 112628 29492
rect 31662 29384 31668 29436
rect 31720 29424 31726 29436
rect 40589 29427 40647 29433
rect 40589 29424 40601 29427
rect 31720 29396 40601 29424
rect 31720 29384 31726 29396
rect 40589 29393 40601 29396
rect 40635 29393 40647 29427
rect 40589 29387 40647 29393
rect 40681 29427 40739 29433
rect 40681 29393 40693 29427
rect 40727 29424 40739 29427
rect 60918 29424 60924 29436
rect 40727 29396 60924 29424
rect 40727 29393 40739 29396
rect 40681 29387 40739 29393
rect 60918 29384 60924 29396
rect 60976 29384 60982 29436
rect 64782 29384 64788 29436
rect 64840 29424 64846 29436
rect 89438 29424 89444 29436
rect 64840 29396 89444 29424
rect 64840 29384 64846 29396
rect 89438 29384 89444 29396
rect 89496 29384 89502 29436
rect 91002 29384 91008 29436
rect 91060 29424 91066 29436
rect 105265 29427 105323 29433
rect 105265 29424 105277 29427
rect 91060 29396 105277 29424
rect 91060 29384 91066 29396
rect 105265 29393 105277 29396
rect 105311 29393 105323 29427
rect 107286 29424 107292 29436
rect 105265 29387 105323 29393
rect 105372 29396 107292 29424
rect 24762 29316 24768 29368
rect 24820 29356 24826 29368
rect 53558 29356 53564 29368
rect 24820 29328 53564 29356
rect 24820 29316 24826 29328
rect 53558 29316 53564 29328
rect 53616 29316 53622 29368
rect 53742 29316 53748 29368
rect 53800 29356 53806 29368
rect 79870 29356 79876 29368
rect 53800 29328 79876 29356
rect 53800 29316 53806 29328
rect 79870 29316 79876 29328
rect 79928 29316 79934 29368
rect 85482 29316 85488 29368
rect 85540 29356 85546 29368
rect 105372 29356 105400 29396
rect 107286 29384 107292 29396
rect 107344 29384 107350 29436
rect 107473 29427 107531 29433
rect 107473 29393 107485 29427
rect 107519 29424 107531 29427
rect 108500 29424 108528 29464
rect 112622 29452 112628 29464
rect 112680 29452 112686 29504
rect 114462 29452 114468 29504
rect 114520 29492 114526 29504
rect 133690 29492 133696 29504
rect 114520 29464 133696 29492
rect 114520 29452 114526 29464
rect 133690 29452 133696 29464
rect 133748 29452 133754 29504
rect 140682 29452 140688 29504
rect 140740 29492 140746 29504
rect 156874 29492 156880 29504
rect 140740 29464 156880 29492
rect 140740 29452 140746 29464
rect 156874 29452 156880 29464
rect 156932 29452 156938 29504
rect 160002 29452 160008 29504
rect 160060 29492 160066 29504
rect 173802 29492 173808 29504
rect 160060 29464 173808 29492
rect 160060 29452 160066 29464
rect 173802 29452 173808 29464
rect 173860 29452 173866 29504
rect 176562 29452 176568 29504
rect 176620 29492 176626 29504
rect 188522 29492 188528 29504
rect 176620 29464 188528 29492
rect 176620 29452 176626 29464
rect 188522 29452 188528 29464
rect 188580 29452 188586 29504
rect 191742 29452 191748 29504
rect 191800 29492 191806 29504
rect 202230 29492 202236 29504
rect 191800 29464 202236 29492
rect 191800 29452 191806 29464
rect 202230 29452 202236 29464
rect 202288 29452 202294 29504
rect 266262 29452 266268 29504
rect 266320 29492 266326 29504
rect 268746 29492 268752 29504
rect 266320 29464 268752 29492
rect 266320 29452 266326 29464
rect 268746 29452 268752 29464
rect 268804 29452 268810 29504
rect 107519 29396 108528 29424
rect 107519 29393 107531 29396
rect 107473 29387 107531 29393
rect 110322 29384 110328 29436
rect 110380 29424 110386 29436
rect 129458 29424 129464 29436
rect 110380 29396 129464 29424
rect 110380 29384 110386 29396
rect 129458 29384 129464 29396
rect 129516 29384 129522 29436
rect 129642 29384 129648 29436
rect 129700 29424 129706 29436
rect 147398 29424 147404 29436
rect 129700 29396 147404 29424
rect 129700 29384 129706 29396
rect 147398 29384 147404 29396
rect 147456 29384 147462 29436
rect 153102 29384 153108 29436
rect 153160 29424 153166 29436
rect 167454 29424 167460 29436
rect 153160 29396 167460 29424
rect 153160 29384 153166 29396
rect 167454 29384 167460 29396
rect 167512 29384 167518 29436
rect 169662 29384 169668 29436
rect 169720 29424 169726 29436
rect 183278 29424 183284 29436
rect 169720 29396 183284 29424
rect 169720 29384 169726 29396
rect 183278 29384 183284 29396
rect 183336 29384 183342 29436
rect 184842 29384 184848 29436
rect 184900 29424 184906 29436
rect 195790 29424 195796 29436
rect 184900 29396 195796 29424
rect 184900 29384 184906 29396
rect 195790 29384 195796 29396
rect 195848 29384 195854 29436
rect 85540 29328 105400 29356
rect 85540 29316 85546 29328
rect 106182 29316 106188 29368
rect 106240 29356 106246 29368
rect 126330 29356 126336 29368
rect 106240 29328 126336 29356
rect 106240 29316 106246 29328
rect 126330 29316 126336 29328
rect 126388 29316 126394 29368
rect 126882 29316 126888 29368
rect 126940 29356 126946 29368
rect 144270 29356 144276 29368
rect 126940 29328 144276 29356
rect 126940 29316 126946 29328
rect 144270 29316 144276 29328
rect 144328 29316 144334 29368
rect 150342 29316 150348 29368
rect 150400 29356 150406 29368
rect 165338 29356 165344 29368
rect 150400 29328 165344 29356
rect 150400 29316 150406 29328
rect 165338 29316 165344 29328
rect 165396 29316 165402 29368
rect 19242 29248 19248 29300
rect 19300 29288 19306 29300
rect 39853 29291 39911 29297
rect 39853 29288 39865 29291
rect 19300 29260 39865 29288
rect 19300 29248 19306 29260
rect 39853 29257 39865 29260
rect 39899 29257 39911 29291
rect 39853 29251 39911 29257
rect 39942 29248 39948 29300
rect 40000 29288 40006 29300
rect 50433 29291 50491 29297
rect 50433 29288 50445 29291
rect 40000 29260 50445 29288
rect 40000 29248 40006 29260
rect 50433 29257 50445 29260
rect 50479 29257 50491 29291
rect 50433 29251 50491 29257
rect 61930 29248 61936 29300
rect 61988 29288 61994 29300
rect 86218 29288 86224 29300
rect 61988 29260 86224 29288
rect 61988 29248 61994 29260
rect 86218 29248 86224 29260
rect 86276 29248 86282 29300
rect 95142 29248 95148 29300
rect 95200 29288 95206 29300
rect 116854 29288 116860 29300
rect 95200 29260 116860 29288
rect 95200 29248 95206 29260
rect 116854 29248 116860 29260
rect 116912 29248 116918 29300
rect 118970 29288 118976 29300
rect 116964 29260 118976 29288
rect 28902 29180 28908 29232
rect 28960 29220 28966 29232
rect 56686 29220 56692 29232
rect 28960 29192 56692 29220
rect 28960 29180 28966 29192
rect 56686 29180 56692 29192
rect 56744 29180 56750 29232
rect 60642 29180 60648 29232
rect 60700 29220 60706 29232
rect 85206 29220 85212 29232
rect 60700 29192 85212 29220
rect 60700 29180 60706 29192
rect 85206 29180 85212 29192
rect 85264 29180 85270 29232
rect 97902 29180 97908 29232
rect 97960 29220 97966 29232
rect 116964 29220 116992 29260
rect 118970 29248 118976 29260
rect 119028 29248 119034 29300
rect 121362 29248 121368 29300
rect 121420 29288 121426 29300
rect 140038 29288 140044 29300
rect 121420 29260 140044 29288
rect 121420 29248 121426 29260
rect 140038 29248 140044 29260
rect 140096 29248 140102 29300
rect 142062 29248 142068 29300
rect 142120 29288 142126 29300
rect 157978 29288 157984 29300
rect 142120 29260 157984 29288
rect 142120 29248 142126 29260
rect 157978 29248 157984 29260
rect 158036 29248 158042 29300
rect 161382 29248 161388 29300
rect 161440 29288 161446 29300
rect 174814 29288 174820 29300
rect 161440 29260 174820 29288
rect 161440 29248 161446 29260
rect 174814 29248 174820 29260
rect 174872 29248 174878 29300
rect 234522 29248 234528 29300
rect 234580 29288 234586 29300
rect 240226 29288 240232 29300
rect 234580 29260 240232 29288
rect 234580 29248 234586 29260
rect 240226 29248 240232 29260
rect 240284 29248 240290 29300
rect 267550 29248 267556 29300
rect 267608 29288 267614 29300
rect 269758 29288 269764 29300
rect 267608 29260 269764 29288
rect 267608 29248 267614 29260
rect 269758 29248 269764 29260
rect 269816 29248 269822 29300
rect 97960 29192 116992 29220
rect 97960 29180 97966 29192
rect 117222 29180 117228 29232
rect 117280 29220 117286 29232
rect 135806 29220 135812 29232
rect 117280 29192 135812 29220
rect 117280 29180 117286 29192
rect 135806 29180 135812 29192
rect 135864 29180 135870 29232
rect 136542 29180 136548 29232
rect 136600 29220 136606 29232
rect 152642 29220 152648 29232
rect 136600 29192 152648 29220
rect 136600 29180 136606 29192
rect 152642 29180 152648 29192
rect 152700 29180 152706 29232
rect 241422 29180 241428 29232
rect 241480 29220 241486 29232
rect 246574 29220 246580 29232
rect 241480 29192 246580 29220
rect 241480 29180 241486 29192
rect 246574 29180 246580 29192
rect 246632 29180 246638 29232
rect 249702 29180 249708 29232
rect 249760 29220 249766 29232
rect 253934 29220 253940 29232
rect 249760 29192 253940 29220
rect 249760 29180 249766 29192
rect 253934 29180 253940 29192
rect 253992 29180 253998 29232
rect 262122 29180 262128 29232
rect 262180 29220 262186 29232
rect 265526 29220 265532 29232
rect 262180 29192 265532 29220
rect 262180 29180 262186 29192
rect 265526 29180 265532 29192
rect 265584 29180 265590 29232
rect 270402 29180 270408 29232
rect 270460 29220 270466 29232
rect 272886 29220 272892 29232
rect 270460 29192 272892 29220
rect 270460 29180 270466 29192
rect 272886 29180 272892 29192
rect 272944 29180 272950 29232
rect 26142 29112 26148 29164
rect 26200 29152 26206 29164
rect 46753 29155 46811 29161
rect 46753 29152 46765 29155
rect 26200 29124 46765 29152
rect 26200 29112 26206 29124
rect 46753 29121 46765 29124
rect 46799 29121 46811 29155
rect 46753 29115 46811 29121
rect 46842 29112 46848 29164
rect 46900 29152 46906 29164
rect 50525 29155 50583 29161
rect 50525 29152 50537 29155
rect 46900 29124 50537 29152
rect 46900 29112 46906 29124
rect 50525 29121 50537 29124
rect 50571 29121 50583 29155
rect 50525 29115 50583 29121
rect 74442 29112 74448 29164
rect 74500 29152 74506 29164
rect 97810 29152 97816 29164
rect 74500 29124 97816 29152
rect 74500 29112 74506 29124
rect 97810 29112 97816 29124
rect 97868 29112 97874 29164
rect 103422 29112 103428 29164
rect 103480 29152 103486 29164
rect 123110 29152 123116 29164
rect 103480 29124 123116 29152
rect 103480 29112 103486 29124
rect 123110 29112 123116 29124
rect 123168 29112 123174 29164
rect 135162 29112 135168 29164
rect 135220 29152 135226 29164
rect 151630 29152 151636 29164
rect 135220 29124 151636 29152
rect 135220 29112 135226 29124
rect 151630 29112 151636 29124
rect 151688 29112 151694 29164
rect 151722 29112 151728 29164
rect 151780 29152 151786 29164
rect 166350 29152 166356 29164
rect 151780 29124 166356 29152
rect 151780 29112 151786 29124
rect 166350 29112 166356 29124
rect 166408 29112 166414 29164
rect 210970 29112 210976 29164
rect 211028 29152 211034 29164
rect 219158 29152 219164 29164
rect 211028 29124 219164 29152
rect 211028 29112 211034 29124
rect 219158 29112 219164 29124
rect 219216 29112 219222 29164
rect 230382 29112 230388 29164
rect 230440 29152 230446 29164
rect 237098 29152 237104 29164
rect 230440 29124 237104 29152
rect 230440 29112 230446 29124
rect 237098 29112 237104 29124
rect 237156 29112 237162 29164
rect 240042 29112 240048 29164
rect 240100 29152 240106 29164
rect 245470 29152 245476 29164
rect 240100 29124 245476 29152
rect 240100 29112 240106 29124
rect 245470 29112 245476 29124
rect 245528 29112 245534 29164
rect 245562 29112 245568 29164
rect 245620 29152 245626 29164
rect 250806 29152 250812 29164
rect 245620 29124 250812 29152
rect 245620 29112 245626 29124
rect 250806 29112 250812 29124
rect 250864 29112 250870 29164
rect 252462 29112 252468 29164
rect 252520 29152 252526 29164
rect 256050 29152 256056 29164
rect 252520 29124 256056 29152
rect 252520 29112 252526 29124
rect 256050 29112 256056 29124
rect 256108 29112 256114 29164
rect 260650 29112 260656 29164
rect 260708 29152 260714 29164
rect 263410 29152 263416 29164
rect 260708 29124 263416 29152
rect 260708 29112 260714 29124
rect 263410 29112 263416 29124
rect 263468 29112 263474 29164
rect 264882 29112 264888 29164
rect 264940 29152 264946 29164
rect 267642 29152 267648 29164
rect 264940 29124 267648 29152
rect 264940 29112 264946 29124
rect 267642 29112 267648 29124
rect 267700 29112 267706 29164
rect 271782 29112 271788 29164
rect 271840 29152 271846 29164
rect 273990 29152 273996 29164
rect 271840 29124 273996 29152
rect 271840 29112 271846 29124
rect 273990 29112 273996 29124
rect 274048 29112 274054 29164
rect 274542 29112 274548 29164
rect 274600 29152 274606 29164
rect 276106 29152 276112 29164
rect 274600 29124 276112 29152
rect 274600 29112 274606 29124
rect 276106 29112 276112 29124
rect 276164 29112 276170 29164
rect 277210 29112 277216 29164
rect 277268 29152 277274 29164
rect 279234 29152 279240 29164
rect 277268 29124 279240 29152
rect 277268 29112 277274 29124
rect 279234 29112 279240 29124
rect 279292 29112 279298 29164
rect 281442 29112 281448 29164
rect 281500 29152 281506 29164
rect 282454 29152 282460 29164
rect 281500 29124 282460 29152
rect 281500 29112 281506 29124
rect 282454 29112 282460 29124
rect 282512 29112 282518 29164
rect 289906 29112 289912 29164
rect 289964 29152 289970 29164
rect 290826 29152 290832 29164
rect 289964 29124 290832 29152
rect 289964 29112 289970 29124
rect 290826 29112 290832 29124
rect 290884 29112 290890 29164
rect 296714 29112 296720 29164
rect 296772 29152 296778 29164
rect 297174 29152 297180 29164
rect 296772 29124 297180 29152
rect 296772 29112 296778 29124
rect 297174 29112 297180 29124
rect 297232 29112 297238 29164
rect 299566 29112 299572 29164
rect 299624 29152 299630 29164
rect 300302 29152 300308 29164
rect 299624 29124 300308 29152
rect 299624 29112 299630 29124
rect 300302 29112 300308 29124
rect 300360 29112 300366 29164
rect 305638 29112 305644 29164
rect 305696 29152 305702 29164
rect 306282 29152 306288 29164
rect 305696 29124 306288 29152
rect 305696 29112 305702 29124
rect 306282 29112 306288 29124
rect 306340 29112 306346 29164
rect 306650 29112 306656 29164
rect 306708 29152 306714 29164
rect 307662 29152 307668 29164
rect 306708 29124 307668 29152
rect 306708 29112 306714 29124
rect 307662 29112 307668 29124
rect 307720 29112 307726 29164
rect 309870 29112 309876 29164
rect 309928 29152 309934 29164
rect 310422 29152 310428 29164
rect 309928 29124 310428 29152
rect 309928 29112 309934 29124
rect 310422 29112 310428 29124
rect 310480 29112 310486 29164
rect 310882 29112 310888 29164
rect 310940 29152 310946 29164
rect 311802 29152 311808 29164
rect 310940 29124 311808 29152
rect 310940 29112 310946 29124
rect 311802 29112 311808 29124
rect 311860 29112 311866 29164
rect 316126 29112 316132 29164
rect 316184 29152 316190 29164
rect 317322 29152 317328 29164
rect 316184 29124 317328 29152
rect 316184 29112 316190 29124
rect 317322 29112 317328 29124
rect 317380 29112 317386 29164
rect 318242 29112 318248 29164
rect 318300 29152 318306 29164
rect 318702 29152 318708 29164
rect 318300 29124 318708 29152
rect 318300 29112 318306 29124
rect 318702 29112 318708 29124
rect 318760 29112 318766 29164
rect 320358 29112 320364 29164
rect 320416 29152 320422 29164
rect 321278 29152 321284 29164
rect 320416 29124 321284 29152
rect 320416 29112 320422 29124
rect 321278 29112 321284 29124
rect 321336 29112 321342 29164
rect 323578 29112 323584 29164
rect 323636 29152 323642 29164
rect 324222 29152 324228 29164
rect 323636 29124 324228 29152
rect 323636 29112 323642 29124
rect 324222 29112 324228 29124
rect 324280 29112 324286 29164
rect 327810 29112 327816 29164
rect 327868 29152 327874 29164
rect 328362 29152 328368 29164
rect 327868 29124 328368 29152
rect 327868 29112 327874 29124
rect 328362 29112 328368 29124
rect 328420 29112 328426 29164
rect 328822 29112 328828 29164
rect 328880 29152 328886 29164
rect 329742 29152 329748 29164
rect 328880 29124 329748 29152
rect 328880 29112 328886 29124
rect 329742 29112 329748 29124
rect 329800 29112 329806 29164
rect 329834 29112 329840 29164
rect 329892 29152 329898 29164
rect 331122 29152 331128 29164
rect 329892 29124 331128 29152
rect 329892 29112 329898 29124
rect 331122 29112 331128 29124
rect 331180 29112 331186 29164
rect 331950 29112 331956 29164
rect 332008 29152 332014 29164
rect 332502 29152 332508 29164
rect 332008 29124 332508 29152
rect 332008 29112 332014 29124
rect 332502 29112 332508 29124
rect 332560 29112 332566 29164
rect 333054 29112 333060 29164
rect 333112 29152 333118 29164
rect 333882 29152 333888 29164
rect 333112 29124 333888 29152
rect 333112 29112 333118 29124
rect 333882 29112 333888 29124
rect 333940 29112 333946 29164
rect 334066 29112 334072 29164
rect 334124 29152 334130 29164
rect 335078 29152 335084 29164
rect 334124 29124 335084 29152
rect 334124 29112 334130 29124
rect 335078 29112 335084 29124
rect 335136 29112 335142 29164
rect 336182 29112 336188 29164
rect 336240 29152 336246 29164
rect 336642 29152 336648 29164
rect 336240 29124 336648 29152
rect 336240 29112 336246 29124
rect 336642 29112 336648 29124
rect 336700 29112 336706 29164
rect 337286 29112 337292 29164
rect 337344 29152 337350 29164
rect 338022 29152 338028 29164
rect 337344 29124 338028 29152
rect 337344 29112 337350 29124
rect 338022 29112 338028 29124
rect 338080 29112 338086 29164
rect 338298 29112 338304 29164
rect 338356 29152 338362 29164
rect 339310 29152 339316 29164
rect 338356 29124 339316 29152
rect 338356 29112 338362 29124
rect 339310 29112 339316 29124
rect 339368 29112 339374 29164
rect 341518 29112 341524 29164
rect 341576 29152 341582 29164
rect 342162 29152 342168 29164
rect 341576 29124 342168 29152
rect 341576 29112 341582 29124
rect 342162 29112 342168 29124
rect 342220 29112 342226 29164
rect 342530 29112 342536 29164
rect 342588 29152 342594 29164
rect 343542 29152 343548 29164
rect 342588 29124 343548 29152
rect 342588 29112 342594 29124
rect 343542 29112 343548 29124
rect 343600 29112 343606 29164
rect 345658 29112 345664 29164
rect 345716 29152 345722 29164
rect 346302 29152 346308 29164
rect 345716 29124 346308 29152
rect 345716 29112 345722 29124
rect 346302 29112 346308 29124
rect 346360 29112 346366 29164
rect 346762 29112 346768 29164
rect 346820 29152 346826 29164
rect 347682 29152 347688 29164
rect 346820 29124 347688 29152
rect 346820 29112 346826 29124
rect 347682 29112 347688 29124
rect 347740 29112 347746 29164
rect 350994 29112 351000 29164
rect 351052 29152 351058 29164
rect 351822 29152 351828 29164
rect 351052 29124 351828 29152
rect 351052 29112 351058 29124
rect 351822 29112 351828 29124
rect 351880 29112 351886 29164
rect 352006 29112 352012 29164
rect 352064 29152 352070 29164
rect 353202 29152 353208 29164
rect 352064 29124 353208 29152
rect 352064 29112 352070 29124
rect 353202 29112 353208 29124
rect 353260 29112 353266 29164
rect 354122 29112 354128 29164
rect 354180 29152 354186 29164
rect 354582 29152 354588 29164
rect 354180 29124 354588 29152
rect 354180 29112 354186 29124
rect 354582 29112 354588 29124
rect 354640 29112 354646 29164
rect 356238 29112 356244 29164
rect 356296 29152 356302 29164
rect 357250 29152 357256 29164
rect 356296 29124 357256 29152
rect 356296 29112 356302 29124
rect 357250 29112 357256 29124
rect 357308 29112 357314 29164
rect 359366 29112 359372 29164
rect 359424 29152 359430 29164
rect 360102 29152 360108 29164
rect 359424 29124 360108 29152
rect 359424 29112 359430 29124
rect 360102 29112 360108 29124
rect 360160 29112 360166 29164
rect 360470 29112 360476 29164
rect 360528 29152 360534 29164
rect 361390 29152 361396 29164
rect 360528 29124 361396 29152
rect 360528 29112 360534 29124
rect 361390 29112 361396 29124
rect 361448 29112 361454 29164
rect 363598 29112 363604 29164
rect 363656 29152 363662 29164
rect 364242 29152 364248 29164
rect 363656 29124 364248 29152
rect 363656 29112 363662 29124
rect 364242 29112 364248 29124
rect 364300 29112 364306 29164
rect 364702 29112 364708 29164
rect 364760 29152 364766 29164
rect 365622 29152 365628 29164
rect 364760 29124 365628 29152
rect 364760 29112 364766 29124
rect 365622 29112 365628 29124
rect 365680 29112 365686 29164
rect 365714 29112 365720 29164
rect 365772 29152 365778 29164
rect 367002 29152 367008 29164
rect 365772 29124 367008 29152
rect 365772 29112 365778 29124
rect 367002 29112 367008 29124
rect 367060 29112 367066 29164
rect 367830 29112 367836 29164
rect 367888 29152 367894 29164
rect 368382 29152 368388 29164
rect 367888 29124 368388 29152
rect 367888 29112 367894 29124
rect 368382 29112 368388 29124
rect 368440 29112 368446 29164
rect 368934 29112 368940 29164
rect 368992 29152 368998 29164
rect 369762 29152 369768 29164
rect 368992 29124 369768 29152
rect 368992 29112 368998 29124
rect 369762 29112 369768 29124
rect 369820 29112 369826 29164
rect 369946 29112 369952 29164
rect 370004 29152 370010 29164
rect 370958 29152 370964 29164
rect 370004 29124 370964 29152
rect 370004 29112 370010 29124
rect 370958 29112 370964 29124
rect 371016 29112 371022 29164
rect 372062 29112 372068 29164
rect 372120 29152 372126 29164
rect 372522 29152 372528 29164
rect 372120 29124 372528 29152
rect 372120 29112 372126 29124
rect 372522 29112 372528 29124
rect 372580 29112 372586 29164
rect 373166 29112 373172 29164
rect 373224 29152 373230 29164
rect 373902 29152 373908 29164
rect 373224 29124 373908 29152
rect 373224 29112 373230 29124
rect 373902 29112 373908 29124
rect 373960 29112 373966 29164
rect 374178 29112 374184 29164
rect 374236 29152 374242 29164
rect 375282 29152 375288 29164
rect 374236 29124 375288 29152
rect 374236 29112 374242 29124
rect 375282 29112 375288 29124
rect 375340 29112 375346 29164
rect 377306 29112 377312 29164
rect 377364 29152 377370 29164
rect 378042 29152 378048 29164
rect 377364 29124 378048 29152
rect 377364 29112 377370 29124
rect 378042 29112 378048 29124
rect 378100 29112 378106 29164
rect 378410 29112 378416 29164
rect 378468 29152 378474 29164
rect 379238 29152 379244 29164
rect 378468 29124 379244 29152
rect 378468 29112 378474 29124
rect 379238 29112 379244 29124
rect 379296 29112 379302 29164
rect 381538 29112 381544 29164
rect 381596 29152 381602 29164
rect 382182 29152 382188 29164
rect 381596 29124 382188 29152
rect 381596 29112 381602 29124
rect 382182 29112 382188 29124
rect 382240 29112 382246 29164
rect 382642 29112 382648 29164
rect 382700 29152 382706 29164
rect 383562 29152 383568 29164
rect 382700 29124 383568 29152
rect 382700 29112 382706 29124
rect 383562 29112 383568 29124
rect 383620 29112 383626 29164
rect 386874 29112 386880 29164
rect 386932 29152 386938 29164
rect 387702 29152 387708 29164
rect 386932 29124 387708 29152
rect 386932 29112 386938 29124
rect 387702 29112 387708 29124
rect 387760 29112 387766 29164
rect 387886 29112 387892 29164
rect 387944 29152 387950 29164
rect 388898 29152 388904 29164
rect 387944 29124 388904 29152
rect 387944 29112 387950 29124
rect 388898 29112 388904 29124
rect 388956 29112 388962 29164
rect 390002 29112 390008 29164
rect 390060 29152 390066 29164
rect 390462 29152 390468 29164
rect 390060 29124 390468 29152
rect 390060 29112 390066 29124
rect 390462 29112 390468 29124
rect 390520 29112 390526 29164
rect 391014 29112 391020 29164
rect 391072 29152 391078 29164
rect 391842 29152 391848 29164
rect 391072 29124 391848 29152
rect 391072 29112 391078 29124
rect 391842 29112 391848 29124
rect 391900 29112 391906 29164
rect 392118 29112 392124 29164
rect 392176 29152 392182 29164
rect 393038 29152 393044 29164
rect 392176 29124 393044 29152
rect 392176 29112 392182 29124
rect 393038 29112 393044 29124
rect 393096 29112 393102 29164
rect 395246 29112 395252 29164
rect 395304 29152 395310 29164
rect 395982 29152 395988 29164
rect 395304 29124 395988 29152
rect 395304 29112 395310 29124
rect 395982 29112 395988 29124
rect 396040 29112 396046 29164
rect 396350 29112 396356 29164
rect 396408 29152 396414 29164
rect 397270 29152 397276 29164
rect 396408 29124 397276 29152
rect 396408 29112 396414 29124
rect 397270 29112 397276 29124
rect 397328 29112 397334 29164
rect 399478 29112 399484 29164
rect 399536 29152 399542 29164
rect 400122 29152 400128 29164
rect 399536 29124 400128 29152
rect 399536 29112 399542 29124
rect 400122 29112 400128 29124
rect 400180 29112 400186 29164
rect 400582 29112 400588 29164
rect 400640 29152 400646 29164
rect 401502 29152 401508 29164
rect 400640 29124 401508 29152
rect 400640 29112 400646 29124
rect 401502 29112 401508 29124
rect 401560 29112 401566 29164
rect 403710 29112 403716 29164
rect 403768 29152 403774 29164
rect 404262 29152 404268 29164
rect 403768 29124 404268 29152
rect 403768 29112 403774 29124
rect 404262 29112 404268 29124
rect 404320 29112 404326 29164
rect 404722 29112 404728 29164
rect 404780 29152 404786 29164
rect 405642 29152 405648 29164
rect 404780 29124 405648 29152
rect 404780 29112 404786 29124
rect 405642 29112 405648 29124
rect 405700 29112 405706 29164
rect 407942 29112 407948 29164
rect 408000 29152 408006 29164
rect 408402 29152 408408 29164
rect 408000 29124 408408 29152
rect 408000 29112 408006 29124
rect 408402 29112 408408 29124
rect 408460 29112 408466 29164
rect 408954 29112 408960 29164
rect 409012 29152 409018 29164
rect 409782 29152 409788 29164
rect 409012 29124 409788 29152
rect 409012 29112 409018 29124
rect 409782 29112 409788 29124
rect 409840 29112 409846 29164
rect 410058 29112 410064 29164
rect 410116 29152 410122 29164
rect 411162 29152 411168 29164
rect 410116 29124 411168 29152
rect 410116 29112 410122 29124
rect 411162 29112 411168 29124
rect 411220 29112 411226 29164
rect 414290 29112 414296 29164
rect 414348 29152 414354 29164
rect 415118 29152 415124 29164
rect 414348 29124 415124 29152
rect 414348 29112 414354 29124
rect 415118 29112 415124 29124
rect 415176 29112 415182 29164
rect 417418 29112 417424 29164
rect 417476 29152 417482 29164
rect 418062 29152 418068 29164
rect 417476 29124 418068 29152
rect 417476 29112 417482 29124
rect 418062 29112 418068 29124
rect 418120 29112 418126 29164
rect 418522 29112 418528 29164
rect 418580 29152 418586 29164
rect 419442 29152 419448 29164
rect 418580 29124 419448 29152
rect 418580 29112 418586 29124
rect 419442 29112 419448 29124
rect 419500 29112 419506 29164
rect 419534 29112 419540 29164
rect 419592 29152 419598 29164
rect 420822 29152 420828 29164
rect 419592 29124 420828 29152
rect 419592 29112 419598 29124
rect 420822 29112 420828 29124
rect 420880 29112 420886 29164
rect 421650 29112 421656 29164
rect 421708 29152 421714 29164
rect 422202 29152 422208 29164
rect 421708 29124 422208 29152
rect 421708 29112 421714 29124
rect 422202 29112 422208 29124
rect 422260 29112 422266 29164
rect 422662 29112 422668 29164
rect 422720 29152 422726 29164
rect 423582 29152 423588 29164
rect 422720 29124 423588 29152
rect 422720 29112 422726 29124
rect 423582 29112 423588 29124
rect 423640 29112 423646 29164
rect 423766 29112 423772 29164
rect 423824 29152 423830 29164
rect 424962 29152 424968 29164
rect 423824 29124 424968 29152
rect 423824 29112 423830 29124
rect 424962 29112 424968 29124
rect 425020 29112 425026 29164
rect 425882 29112 425888 29164
rect 425940 29152 425946 29164
rect 426342 29152 426348 29164
rect 425940 29124 426348 29152
rect 425940 29112 425946 29124
rect 426342 29112 426348 29124
rect 426400 29112 426406 29164
rect 426894 29112 426900 29164
rect 426952 29152 426958 29164
rect 427722 29152 427728 29164
rect 426952 29124 427728 29152
rect 426952 29112 426958 29124
rect 427722 29112 427728 29124
rect 427780 29112 427786 29164
rect 427998 29112 428004 29164
rect 428056 29152 428062 29164
rect 428918 29152 428924 29164
rect 428056 29124 428924 29152
rect 428056 29112 428062 29124
rect 428918 29112 428924 29124
rect 428976 29112 428982 29164
rect 435358 29112 435364 29164
rect 435416 29152 435422 29164
rect 436002 29152 436008 29164
rect 435416 29124 436008 29152
rect 435416 29112 435422 29124
rect 436002 29112 436008 29124
rect 436060 29112 436066 29164
rect 436370 29112 436376 29164
rect 436428 29152 436434 29164
rect 437382 29152 437388 29164
rect 436428 29124 437388 29152
rect 436428 29112 436434 29124
rect 437382 29112 437388 29124
rect 437440 29112 437446 29164
rect 437474 29112 437480 29164
rect 437532 29152 437538 29164
rect 438762 29152 438768 29164
rect 437532 29124 438768 29152
rect 437532 29112 437538 29124
rect 438762 29112 438768 29124
rect 438820 29112 438826 29164
rect 439590 29112 439596 29164
rect 439648 29152 439654 29164
rect 440142 29152 440148 29164
rect 439648 29124 440148 29152
rect 439648 29112 439654 29124
rect 440142 29112 440148 29124
rect 440200 29112 440206 29164
rect 440602 29112 440608 29164
rect 440660 29152 440666 29164
rect 441522 29152 441528 29164
rect 440660 29124 441528 29152
rect 440660 29112 440666 29124
rect 441522 29112 441528 29124
rect 441580 29112 441586 29164
rect 441706 29112 441712 29164
rect 441764 29152 441770 29164
rect 442902 29152 442908 29164
rect 441764 29124 442908 29152
rect 441764 29112 441770 29124
rect 442902 29112 442908 29124
rect 442960 29112 442966 29164
rect 443822 29112 443828 29164
rect 443880 29152 443886 29164
rect 444282 29152 444288 29164
rect 443880 29124 444288 29152
rect 443880 29112 443886 29124
rect 444282 29112 444288 29124
rect 444340 29112 444346 29164
rect 444834 29112 444840 29164
rect 444892 29152 444898 29164
rect 445662 29152 445668 29164
rect 444892 29124 445668 29152
rect 444892 29112 444898 29124
rect 445662 29112 445668 29124
rect 445720 29112 445726 29164
rect 445938 29112 445944 29164
rect 445996 29152 446002 29164
rect 446858 29152 446864 29164
rect 445996 29124 446864 29152
rect 445996 29112 446002 29124
rect 446858 29112 446864 29124
rect 446916 29112 446922 29164
rect 449066 29112 449072 29164
rect 449124 29152 449130 29164
rect 449802 29152 449808 29164
rect 449124 29124 449808 29152
rect 449124 29112 449130 29124
rect 449802 29112 449808 29124
rect 449860 29112 449866 29164
rect 450078 29112 450084 29164
rect 450136 29152 450142 29164
rect 451090 29152 451096 29164
rect 450136 29124 451096 29152
rect 450136 29112 450142 29124
rect 451090 29112 451096 29124
rect 451148 29112 451154 29164
rect 453298 29112 453304 29164
rect 453356 29152 453362 29164
rect 453942 29152 453948 29164
rect 453356 29124 453948 29152
rect 453356 29112 453362 29124
rect 453942 29112 453948 29124
rect 454000 29112 454006 29164
rect 454310 29112 454316 29164
rect 454368 29152 454374 29164
rect 455322 29152 455328 29164
rect 454368 29124 455328 29152
rect 454368 29112 454374 29124
rect 455322 29112 455328 29124
rect 455380 29112 455386 29164
rect 455414 29112 455420 29164
rect 455472 29152 455478 29164
rect 456702 29152 456708 29164
rect 455472 29124 456708 29152
rect 455472 29112 455478 29124
rect 456702 29112 456708 29124
rect 456760 29112 456766 29164
rect 457530 29112 457536 29164
rect 457588 29152 457594 29164
rect 458082 29152 458088 29164
rect 457588 29124 458088 29152
rect 457588 29112 457594 29124
rect 458082 29112 458088 29124
rect 458140 29112 458146 29164
rect 458542 29112 458548 29164
rect 458600 29152 458606 29164
rect 459462 29152 459468 29164
rect 458600 29124 459468 29152
rect 458600 29112 458606 29124
rect 459462 29112 459468 29124
rect 459520 29112 459526 29164
rect 461762 29112 461768 29164
rect 461820 29152 461826 29164
rect 462222 29152 462228 29164
rect 461820 29124 462228 29152
rect 461820 29112 461826 29124
rect 462222 29112 462228 29124
rect 462280 29112 462286 29164
rect 462774 29112 462780 29164
rect 462832 29152 462838 29164
rect 463602 29152 463608 29164
rect 462832 29124 463608 29152
rect 462832 29112 462838 29124
rect 463602 29112 463608 29124
rect 463660 29112 463666 29164
rect 463786 29112 463792 29164
rect 463844 29152 463850 29164
rect 464982 29152 464988 29164
rect 463844 29124 464988 29152
rect 463844 29112 463850 29124
rect 464982 29112 464988 29124
rect 465040 29112 465046 29164
rect 465902 29112 465908 29164
rect 465960 29152 465966 29164
rect 466362 29152 466368 29164
rect 465960 29124 466368 29152
rect 465960 29112 465966 29124
rect 466362 29112 466368 29124
rect 466420 29112 466426 29164
rect 467006 29112 467012 29164
rect 467064 29152 467070 29164
rect 467742 29152 467748 29164
rect 467064 29124 467748 29152
rect 467064 29112 467070 29124
rect 467742 29112 467748 29124
rect 467800 29112 467806 29164
rect 468018 29112 468024 29164
rect 468076 29152 468082 29164
rect 469030 29152 469036 29164
rect 468076 29124 469036 29152
rect 468076 29112 468082 29124
rect 469030 29112 469036 29124
rect 469088 29112 469094 29164
rect 471238 29112 471244 29164
rect 471296 29152 471302 29164
rect 471882 29152 471888 29164
rect 471296 29124 471888 29152
rect 471296 29112 471302 29124
rect 471882 29112 471888 29124
rect 471940 29112 471946 29164
rect 472250 29112 472256 29164
rect 472308 29152 472314 29164
rect 473262 29152 473268 29164
rect 472308 29124 473268 29152
rect 472308 29112 472314 29124
rect 473262 29112 473268 29124
rect 473320 29112 473326 29164
rect 473354 29112 473360 29164
rect 473412 29152 473418 29164
rect 475378 29152 475384 29164
rect 473412 29124 475384 29152
rect 473412 29112 473418 29124
rect 475378 29112 475384 29124
rect 475436 29112 475442 29164
rect 475470 29112 475476 29164
rect 475528 29152 475534 29164
rect 476022 29152 476028 29164
rect 475528 29124 476028 29152
rect 475528 29112 475534 29124
rect 476022 29112 476028 29124
rect 476080 29112 476086 29164
rect 476482 29112 476488 29164
rect 476540 29152 476546 29164
rect 477402 29152 477408 29164
rect 476540 29124 477408 29152
rect 476540 29112 476546 29124
rect 477402 29112 477408 29124
rect 477460 29112 477466 29164
rect 477586 29112 477592 29164
rect 477644 29152 477650 29164
rect 478782 29152 478788 29164
rect 477644 29124 478788 29152
rect 477644 29112 477650 29124
rect 478782 29112 478788 29124
rect 478840 29112 478846 29164
rect 479610 29112 479616 29164
rect 479668 29152 479674 29164
rect 480162 29152 480168 29164
rect 479668 29124 480168 29152
rect 479668 29112 479674 29124
rect 480162 29112 480168 29124
rect 480220 29112 480226 29164
rect 480714 29112 480720 29164
rect 480772 29152 480778 29164
rect 481542 29152 481548 29164
rect 480772 29124 481548 29152
rect 480772 29112 480778 29124
rect 481542 29112 481548 29124
rect 481600 29112 481606 29164
rect 481726 29112 481732 29164
rect 481784 29152 481790 29164
rect 482922 29152 482928 29164
rect 481784 29124 482928 29152
rect 481784 29112 481790 29124
rect 482922 29112 482928 29124
rect 482980 29112 482986 29164
rect 483842 29112 483848 29164
rect 483900 29152 483906 29164
rect 484302 29152 484308 29164
rect 483900 29124 484308 29152
rect 483900 29112 483906 29124
rect 484302 29112 484308 29124
rect 484360 29112 484366 29164
rect 484946 29112 484952 29164
rect 485004 29152 485010 29164
rect 485682 29152 485688 29164
rect 485004 29124 485688 29152
rect 485004 29112 485010 29124
rect 485682 29112 485688 29124
rect 485740 29112 485746 29164
rect 485958 29112 485964 29164
rect 486016 29152 486022 29164
rect 486970 29152 486976 29164
rect 486016 29124 486976 29152
rect 486016 29112 486022 29124
rect 486970 29112 486976 29124
rect 487028 29112 487034 29164
rect 489178 29112 489184 29164
rect 489236 29152 489242 29164
rect 489822 29152 489828 29164
rect 489236 29124 489828 29152
rect 489236 29112 489242 29124
rect 489822 29112 489828 29124
rect 489880 29112 489886 29164
rect 490190 29112 490196 29164
rect 490248 29152 490254 29164
rect 491202 29152 491208 29164
rect 490248 29124 491208 29152
rect 490248 29112 490254 29124
rect 491202 29112 491208 29124
rect 491260 29112 491266 29164
rect 491294 29112 491300 29164
rect 491352 29152 491358 29164
rect 492582 29152 492588 29164
rect 491352 29124 492588 29152
rect 491352 29112 491358 29124
rect 492582 29112 492588 29124
rect 492640 29112 492646 29164
rect 493318 29112 493324 29164
rect 493376 29152 493382 29164
rect 493962 29152 493968 29164
rect 493376 29124 493968 29152
rect 493376 29112 493382 29124
rect 493962 29112 493968 29124
rect 494020 29112 494026 29164
rect 494422 29112 494428 29164
rect 494480 29152 494486 29164
rect 495342 29152 495348 29164
rect 494480 29124 495348 29152
rect 494480 29112 494486 29124
rect 495342 29112 495348 29124
rect 495400 29112 495406 29164
rect 495434 29112 495440 29164
rect 495492 29152 495498 29164
rect 497458 29152 497464 29164
rect 495492 29124 497464 29152
rect 495492 29112 495498 29124
rect 497458 29112 497464 29124
rect 497516 29112 497522 29164
rect 497550 29112 497556 29164
rect 497608 29152 497614 29164
rect 498102 29152 498108 29164
rect 497608 29124 498108 29152
rect 497608 29112 497614 29124
rect 498102 29112 498108 29124
rect 498160 29112 498166 29164
rect 499666 29112 499672 29164
rect 499724 29152 499730 29164
rect 500678 29152 500684 29164
rect 499724 29124 500684 29152
rect 499724 29112 499730 29124
rect 500678 29112 500684 29124
rect 500736 29112 500742 29164
rect 501782 29112 501788 29164
rect 501840 29152 501846 29164
rect 502242 29152 502248 29164
rect 501840 29124 502248 29152
rect 501840 29112 501846 29124
rect 502242 29112 502248 29124
rect 502300 29112 502306 29164
rect 502886 29112 502892 29164
rect 502944 29152 502950 29164
rect 503622 29152 503628 29164
rect 502944 29124 503628 29152
rect 502944 29112 502950 29124
rect 503622 29112 503628 29124
rect 503680 29112 503686 29164
rect 503898 29112 503904 29164
rect 503956 29152 503962 29164
rect 504818 29152 504824 29164
rect 503956 29124 504824 29152
rect 503956 29112 503962 29124
rect 504818 29112 504824 29124
rect 504876 29112 504882 29164
rect 507118 29112 507124 29164
rect 507176 29152 507182 29164
rect 507762 29152 507768 29164
rect 507176 29124 507768 29152
rect 507176 29112 507182 29124
rect 507762 29112 507768 29124
rect 507820 29112 507826 29164
rect 511258 29112 511264 29164
rect 511316 29152 511322 29164
rect 511902 29152 511908 29164
rect 511316 29124 511908 29152
rect 511316 29112 511322 29124
rect 511902 29112 511908 29124
rect 511960 29112 511966 29164
rect 512362 29112 512368 29164
rect 512420 29152 512426 29164
rect 513282 29152 513288 29164
rect 512420 29124 513288 29152
rect 512420 29112 512426 29124
rect 513282 29112 513288 29124
rect 513340 29112 513346 29164
rect 513374 29112 513380 29164
rect 513432 29152 513438 29164
rect 514662 29152 514668 29164
rect 513432 29124 514668 29152
rect 513432 29112 513438 29124
rect 514662 29112 514668 29124
rect 514720 29112 514726 29164
rect 515490 29112 515496 29164
rect 515548 29152 515554 29164
rect 516042 29152 516048 29164
rect 515548 29124 516048 29152
rect 515548 29112 515554 29124
rect 516042 29112 516048 29124
rect 516100 29112 516106 29164
rect 516594 29112 516600 29164
rect 516652 29152 516658 29164
rect 517422 29152 517428 29164
rect 516652 29124 517428 29152
rect 516652 29112 516658 29124
rect 517422 29112 517428 29124
rect 517480 29112 517486 29164
rect 517606 29112 517612 29164
rect 517664 29152 517670 29164
rect 518618 29152 518624 29164
rect 517664 29124 518624 29152
rect 517664 29112 517670 29124
rect 518618 29112 518624 29124
rect 518676 29112 518682 29164
rect 519722 29112 519728 29164
rect 519780 29152 519786 29164
rect 520182 29152 520188 29164
rect 519780 29124 520188 29152
rect 519780 29112 519786 29124
rect 520182 29112 520188 29124
rect 520240 29112 520246 29164
rect 520826 29112 520832 29164
rect 520884 29152 520890 29164
rect 521562 29152 521568 29164
rect 520884 29124 521568 29152
rect 520884 29112 520890 29124
rect 521562 29112 521568 29124
rect 521620 29112 521626 29164
rect 521838 29112 521844 29164
rect 521896 29152 521902 29164
rect 522942 29152 522948 29164
rect 521896 29124 522948 29152
rect 521896 29112 521902 29124
rect 522942 29112 522948 29124
rect 523000 29112 523006 29164
rect 524966 29112 524972 29164
rect 525024 29152 525030 29164
rect 525702 29152 525708 29164
rect 525024 29124 525708 29152
rect 525024 29112 525030 29124
rect 525702 29112 525708 29124
rect 525760 29112 525766 29164
rect 531314 29112 531320 29164
rect 531372 29152 531378 29164
rect 532602 29152 532608 29164
rect 531372 29124 532608 29152
rect 531372 29112 531378 29124
rect 532602 29112 532608 29124
rect 532660 29112 532666 29164
rect 533430 29112 533436 29164
rect 533488 29152 533494 29164
rect 533982 29152 533988 29164
rect 533488 29124 533988 29152
rect 533488 29112 533494 29124
rect 533982 29112 533988 29124
rect 534040 29112 534046 29164
rect 534534 29112 534540 29164
rect 534592 29152 534598 29164
rect 535362 29152 535368 29164
rect 534592 29124 535368 29152
rect 534592 29112 534598 29124
rect 535362 29112 535368 29124
rect 535420 29112 535426 29164
rect 535546 29112 535552 29164
rect 535604 29152 535610 29164
rect 536742 29152 536748 29164
rect 535604 29124 536748 29152
rect 535604 29112 535610 29124
rect 536742 29112 536748 29124
rect 536800 29112 536806 29164
rect 537662 29112 537668 29164
rect 537720 29152 537726 29164
rect 538122 29152 538128 29164
rect 537720 29124 538128 29152
rect 537720 29112 537726 29124
rect 538122 29112 538128 29124
rect 538180 29112 538186 29164
rect 538674 29112 538680 29164
rect 538732 29152 538738 29164
rect 539502 29152 539508 29164
rect 538732 29124 539508 29152
rect 538732 29112 538738 29124
rect 539502 29112 539508 29124
rect 539560 29112 539566 29164
rect 544010 29112 544016 29164
rect 544068 29152 544074 29164
rect 544930 29152 544936 29164
rect 544068 29124 544936 29152
rect 544068 29112 544074 29124
rect 544930 29112 544936 29124
rect 544988 29112 544994 29164
rect 548242 29112 548248 29164
rect 548300 29152 548306 29164
rect 549162 29152 549168 29164
rect 548300 29124 549168 29152
rect 548300 29112 548306 29124
rect 549162 29112 549168 29124
rect 549220 29112 549226 29164
rect 39850 29084 39856 29096
rect 26206 29056 39856 29084
rect 9582 28976 9588 29028
rect 9640 29016 9646 29028
rect 26206 29016 26234 29056
rect 39850 29044 39856 29056
rect 39908 29044 39914 29096
rect 40589 29087 40647 29093
rect 40589 29053 40601 29087
rect 40635 29084 40647 29087
rect 59906 29084 59912 29096
rect 40635 29056 59912 29084
rect 40635 29053 40647 29056
rect 40589 29047 40647 29053
rect 59906 29044 59912 29056
rect 59964 29044 59970 29096
rect 95050 29044 95056 29096
rect 95108 29084 95114 29096
rect 115750 29084 115756 29096
rect 95108 29056 115756 29084
rect 95108 29044 95114 29056
rect 115750 29044 115756 29056
rect 115808 29044 115814 29096
rect 115842 29044 115848 29096
rect 115900 29084 115906 29096
rect 134794 29084 134800 29096
rect 115900 29056 134800 29084
rect 115900 29044 115906 29056
rect 134794 29044 134800 29056
rect 134852 29044 134858 29096
rect 139302 29044 139308 29096
rect 139360 29084 139366 29096
rect 155862 29084 155868 29096
rect 139360 29056 155868 29084
rect 139360 29044 139366 29056
rect 155862 29044 155868 29056
rect 155920 29044 155926 29096
rect 220722 29044 220728 29096
rect 220780 29084 220786 29096
rect 228634 29084 228640 29096
rect 220780 29056 228640 29084
rect 220780 29044 220786 29056
rect 228634 29044 228640 29056
rect 228692 29044 228698 29096
rect 242802 29044 242808 29096
rect 242860 29084 242866 29096
rect 247586 29084 247592 29096
rect 242860 29056 247592 29084
rect 242860 29044 242866 29056
rect 247586 29044 247592 29056
rect 247644 29044 247650 29096
rect 251082 29044 251088 29096
rect 251140 29084 251146 29096
rect 255038 29084 255044 29096
rect 251140 29056 255044 29084
rect 251140 29044 251146 29056
rect 255038 29044 255044 29056
rect 255096 29044 255102 29096
rect 259362 29044 259368 29096
rect 259420 29084 259426 29096
rect 262398 29084 262404 29096
rect 259420 29056 262404 29084
rect 259420 29044 259426 29056
rect 262398 29044 262404 29056
rect 262456 29044 262462 29096
rect 263502 29044 263508 29096
rect 263560 29084 263566 29096
rect 266630 29084 266636 29096
rect 263560 29056 266636 29084
rect 263560 29044 263566 29056
rect 266630 29044 266636 29056
rect 266688 29044 266694 29096
rect 269022 29044 269028 29096
rect 269080 29084 269086 29096
rect 270770 29084 270776 29096
rect 269080 29056 270776 29084
rect 269080 29044 269086 29056
rect 270770 29044 270776 29056
rect 270828 29044 270834 29096
rect 273898 29044 273904 29096
rect 273956 29084 273962 29096
rect 275002 29084 275008 29096
rect 273956 29056 275008 29084
rect 273956 29044 273962 29056
rect 275002 29044 275008 29056
rect 275060 29044 275066 29096
rect 278682 29044 278688 29096
rect 278740 29084 278746 29096
rect 280338 29084 280344 29096
rect 278740 29056 280344 29084
rect 278740 29044 278746 29056
rect 280338 29044 280344 29056
rect 280396 29044 280402 29096
rect 311986 29044 311992 29096
rect 312044 29084 312050 29096
rect 313274 29084 313280 29096
rect 312044 29056 313280 29084
rect 312044 29044 312050 29056
rect 313274 29044 313280 29056
rect 313332 29044 313338 29096
rect 319346 29044 319352 29096
rect 319404 29084 319410 29096
rect 321554 29084 321560 29096
rect 319404 29056 321560 29084
rect 319404 29044 319410 29056
rect 321554 29044 321560 29056
rect 321612 29044 321618 29096
rect 324590 29044 324596 29096
rect 324648 29084 324654 29096
rect 325602 29084 325608 29096
rect 324648 29056 325608 29084
rect 324648 29044 324654 29056
rect 325602 29044 325608 29056
rect 325660 29044 325666 29096
rect 347774 29044 347780 29096
rect 347832 29084 347838 29096
rect 348970 29084 348976 29096
rect 347832 29056 348976 29084
rect 347832 29044 347838 29056
rect 348970 29044 348976 29056
rect 349028 29044 349034 29096
rect 355226 29044 355232 29096
rect 355284 29084 355290 29096
rect 355962 29084 355968 29096
rect 355284 29056 355968 29084
rect 355284 29044 355290 29056
rect 355962 29044 355968 29056
rect 356020 29044 356026 29096
rect 383654 29044 383660 29096
rect 383712 29084 383718 29096
rect 384850 29084 384856 29096
rect 383712 29056 384856 29084
rect 383712 29044 383718 29056
rect 384850 29044 384856 29056
rect 384908 29044 384914 29096
rect 405826 29044 405832 29096
rect 405884 29084 405890 29096
rect 406930 29084 406936 29096
rect 405884 29056 406936 29084
rect 405884 29044 405890 29056
rect 406930 29044 406936 29056
rect 406988 29044 406994 29096
rect 413186 29044 413192 29096
rect 413244 29084 413250 29096
rect 413922 29084 413928 29096
rect 413244 29056 413928 29084
rect 413244 29044 413250 29056
rect 413922 29044 413928 29056
rect 413980 29044 413986 29096
rect 431126 29044 431132 29096
rect 431184 29084 431190 29096
rect 431862 29084 431868 29096
rect 431184 29056 431868 29084
rect 431184 29044 431190 29056
rect 431862 29044 431868 29056
rect 431920 29044 431926 29096
rect 432230 29044 432236 29096
rect 432288 29084 432294 29096
rect 433058 29084 433064 29096
rect 432288 29056 433064 29084
rect 432288 29044 432294 29056
rect 433058 29044 433064 29056
rect 433116 29044 433122 29096
rect 492306 29044 492312 29096
rect 492364 29084 492370 29096
rect 493410 29084 493416 29096
rect 492364 29056 493416 29084
rect 492364 29044 492370 29056
rect 493410 29044 493416 29056
rect 493468 29044 493474 29096
rect 526070 29044 526076 29096
rect 526128 29084 526134 29096
rect 526898 29084 526904 29096
rect 526128 29056 526904 29084
rect 526128 29044 526134 29056
rect 526898 29044 526904 29056
rect 526956 29044 526962 29096
rect 547138 29044 547144 29096
rect 547196 29084 547202 29096
rect 547782 29084 547788 29096
rect 547196 29056 547788 29084
rect 547196 29044 547202 29056
rect 547782 29044 547788 29056
rect 547840 29044 547846 29096
rect 549254 29044 549260 29096
rect 549312 29084 549318 29096
rect 550450 29084 550456 29096
rect 549312 29056 550456 29084
rect 549312 29044 549318 29056
rect 550450 29044 550456 29056
rect 550508 29044 550514 29096
rect 9640 28988 26234 29016
rect 9640 28976 9646 28988
rect 37182 28976 37188 29028
rect 37240 29016 37246 29028
rect 64046 29016 64052 29028
rect 37240 28988 64052 29016
rect 37240 28976 37246 28988
rect 64046 28976 64052 28988
rect 64104 28976 64110 29028
rect 99282 28976 99288 29028
rect 99340 29016 99346 29028
rect 119706 29016 119712 29028
rect 99340 28988 119712 29016
rect 99340 28976 99346 28988
rect 119706 28976 119712 28988
rect 119764 28976 119770 29028
rect 119798 28976 119804 29028
rect 119856 29016 119862 29028
rect 137830 29016 137836 29028
rect 119856 28988 137836 29016
rect 119856 28976 119862 28988
rect 137830 28976 137836 28988
rect 137888 28976 137894 29028
rect 231762 28976 231768 29028
rect 231820 29016 231826 29028
rect 238110 29016 238116 29028
rect 231820 28988 238116 29016
rect 231820 28976 231826 28988
rect 238110 28976 238116 28988
rect 238168 28976 238174 29028
rect 252370 28976 252376 29028
rect 252428 29016 252434 29028
rect 257062 29016 257068 29028
rect 252428 28988 257068 29016
rect 252428 28976 252434 28988
rect 257062 28976 257068 28988
rect 257120 28976 257126 29028
rect 260742 28976 260748 29028
rect 260800 29016 260806 29028
rect 264514 29016 264520 29028
rect 260800 28988 264520 29016
rect 260800 28976 260806 28988
rect 264514 28976 264520 28988
rect 264572 28976 264578 29028
rect 268930 28976 268936 29028
rect 268988 29016 268994 29028
rect 271874 29016 271880 29028
rect 268988 28988 271880 29016
rect 268988 28976 268994 28988
rect 271874 28976 271880 28988
rect 271932 28976 271938 29028
rect 282822 28976 282828 29028
rect 282880 29016 282886 29028
rect 283466 29016 283472 29028
rect 282880 28988 283472 29016
rect 282880 28976 282886 28988
rect 283466 28976 283472 28988
rect 283524 28976 283530 29028
rect 314102 28976 314108 29028
rect 314160 29016 314166 29028
rect 314562 29016 314568 29028
rect 314160 28988 314568 29016
rect 314160 28976 314166 28988
rect 314562 28976 314568 28988
rect 314620 28976 314626 29028
rect 325694 28976 325700 29028
rect 325752 29016 325758 29028
rect 327718 29016 327724 29028
rect 325752 28988 327724 29016
rect 325752 28976 325758 28988
rect 327718 28976 327724 28988
rect 327776 28976 327782 29028
rect 343634 28976 343640 29028
rect 343692 29016 343698 29028
rect 344830 29016 344836 29028
rect 343692 28988 344836 29016
rect 343692 28976 343698 28988
rect 344830 28976 344836 28988
rect 344888 28976 344894 29028
rect 349890 28976 349896 29028
rect 349948 29016 349954 29028
rect 350442 29016 350448 29028
rect 349948 28988 350448 29016
rect 349948 28976 349954 28988
rect 350442 28976 350448 28988
rect 350500 28976 350506 29028
rect 385770 28976 385776 29028
rect 385828 29016 385834 29028
rect 386322 29016 386328 29028
rect 385828 28988 386328 29016
rect 385828 28976 385834 28988
rect 386322 28976 386328 28988
rect 386380 28976 386386 29028
rect 401594 28976 401600 29028
rect 401652 29016 401658 29028
rect 402790 29016 402796 29028
rect 401652 28988 402796 29016
rect 401652 28976 401658 28988
rect 402790 28976 402796 28988
rect 402848 28976 402854 29028
rect 459646 28976 459652 29028
rect 459704 29016 459710 29028
rect 460750 29016 460756 29028
rect 459704 28988 460756 29016
rect 459704 28976 459710 28988
rect 460750 28976 460756 28988
rect 460808 28976 460814 29028
rect 529198 28976 529204 29028
rect 529256 29016 529262 29028
rect 529842 29016 529848 29028
rect 529256 28988 529848 29016
rect 529256 28976 529262 28988
rect 529842 28976 529848 28988
rect 529900 28976 529906 29028
rect 66162 28568 66168 28620
rect 66220 28608 66226 28620
rect 90450 28608 90456 28620
rect 66220 28580 90456 28608
rect 66220 28568 66226 28580
rect 90450 28568 90456 28580
rect 90508 28568 90514 28620
rect 52362 28500 52368 28552
rect 52420 28540 52426 28552
rect 77754 28540 77760 28552
rect 52420 28512 77760 28540
rect 52420 28500 52426 28512
rect 77754 28500 77760 28512
rect 77812 28500 77818 28552
rect 79962 28500 79968 28552
rect 80020 28540 80026 28552
rect 100754 28540 100760 28552
rect 80020 28512 100760 28540
rect 80020 28500 80026 28512
rect 100754 28500 100760 28512
rect 100812 28500 100818 28552
rect 30282 28432 30288 28484
rect 30340 28472 30346 28484
rect 58802 28472 58808 28484
rect 30340 28444 58808 28472
rect 30340 28432 30346 28444
rect 58802 28432 58808 28444
rect 58860 28432 58866 28484
rect 59262 28432 59268 28484
rect 59320 28472 59326 28484
rect 84102 28472 84108 28484
rect 59320 28444 84108 28472
rect 59320 28432 59326 28444
rect 84102 28432 84108 28444
rect 84160 28432 84166 28484
rect 17862 28364 17868 28416
rect 17920 28404 17926 28416
rect 47210 28404 47216 28416
rect 17920 28376 47216 28404
rect 17920 28364 17926 28376
rect 47210 28364 47216 28376
rect 47268 28364 47274 28416
rect 48222 28364 48228 28416
rect 48280 28404 48286 28416
rect 74626 28404 74632 28416
rect 48280 28376 74632 28404
rect 48280 28364 48286 28376
rect 74626 28364 74632 28376
rect 74684 28364 74690 28416
rect 77202 28364 77208 28416
rect 77260 28404 77266 28416
rect 99926 28404 99932 28416
rect 77260 28376 99932 28404
rect 77260 28364 77266 28376
rect 99926 28364 99932 28376
rect 99984 28364 99990 28416
rect 22002 28296 22008 28348
rect 22060 28336 22066 28348
rect 51442 28336 51448 28348
rect 22060 28308 51448 28336
rect 22060 28296 22066 28308
rect 51442 28296 51448 28308
rect 51500 28296 51506 28348
rect 55122 28296 55128 28348
rect 55180 28336 55186 28348
rect 80974 28336 80980 28348
rect 55180 28308 80980 28336
rect 55180 28296 55186 28308
rect 80974 28296 80980 28308
rect 81032 28296 81038 28348
rect 84102 28296 84108 28348
rect 84160 28336 84166 28348
rect 106274 28336 106280 28348
rect 84160 28308 106280 28336
rect 84160 28296 84166 28308
rect 106274 28296 106280 28308
rect 106332 28296 106338 28348
rect 8202 28228 8208 28280
rect 8260 28268 8266 28280
rect 38746 28268 38752 28280
rect 8260 28240 38752 28268
rect 8260 28228 8266 28240
rect 38746 28228 38752 28240
rect 38804 28228 38810 28280
rect 41322 28228 41328 28280
rect 41380 28268 41386 28280
rect 68278 28268 68284 28280
rect 41380 28240 68284 28268
rect 41380 28228 41386 28240
rect 68278 28228 68284 28240
rect 68336 28228 68342 28280
rect 73062 28228 73068 28280
rect 73120 28268 73126 28280
rect 96798 28268 96804 28280
rect 73120 28240 96804 28268
rect 73120 28228 73126 28240
rect 96798 28228 96804 28240
rect 96856 28228 96862 28280
rect 51718 27616 51724 27668
rect 51776 27656 51782 27668
rect 55674 27656 55680 27668
rect 51776 27628 55680 27656
rect 51776 27616 51782 27628
rect 55674 27616 55680 27628
rect 55732 27616 55738 27668
rect 60826 26732 60832 26784
rect 60884 26772 60890 26784
rect 62022 26772 62028 26784
rect 60884 26744 62028 26772
rect 60884 26732 60890 26744
rect 62022 26732 62028 26744
rect 62080 26732 62086 26784
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 18598 20652 18604 20664
rect 3476 20624 18604 20652
rect 3476 20612 3482 20624
rect 18598 20612 18604 20624
rect 18656 20612 18662 20664
rect 552658 20612 552664 20664
rect 552716 20652 552722 20664
rect 579982 20652 579988 20664
rect 552716 20624 579988 20652
rect 552716 20612 552722 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 299566 11704 299572 11756
rect 299624 11744 299630 11756
rect 300762 11744 300768 11756
rect 299624 11716 300768 11744
rect 299624 11704 299630 11716
rect 300762 11704 300768 11716
rect 300820 11704 300826 11756
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 15838 6848 15844 6860
rect 3476 6820 15844 6848
rect 3476 6808 3482 6820
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 555418 6808 555424 6860
rect 555476 6848 555482 6860
rect 580166 6848 580172 6860
rect 555476 6820 580172 6848
rect 555476 6808 555482 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 69106 6128 69112 6180
rect 69164 6168 69170 6180
rect 93578 6168 93584 6180
rect 69164 6140 93584 6168
rect 69164 6128 69170 6140
rect 93578 6128 93584 6140
rect 93636 6128 93642 6180
rect 526990 6128 526996 6180
rect 527048 6168 527054 6180
rect 554958 6168 554964 6180
rect 527048 6140 554964 6168
rect 527048 6128 527054 6140
rect 554958 6128 554964 6140
rect 555016 6128 555022 6180
rect 62206 5244 62212 5296
rect 62264 5284 62270 5296
rect 65150 5284 65156 5296
rect 62264 5256 65156 5284
rect 62264 5244 62270 5256
rect 65150 5244 65156 5256
rect 65208 5244 65214 5296
rect 475378 5244 475384 5296
rect 475436 5284 475442 5296
rect 494698 5284 494704 5296
rect 475436 5256 494704 5284
rect 475436 5244 475442 5256
rect 494698 5244 494704 5256
rect 494756 5244 494762 5296
rect 511350 5244 511356 5296
rect 511408 5284 511414 5296
rect 533706 5284 533712 5296
rect 511408 5256 533712 5284
rect 511408 5244 511414 5256
rect 533706 5244 533712 5256
rect 533764 5244 533770 5296
rect 493410 5176 493416 5228
rect 493468 5216 493474 5228
rect 515950 5216 515956 5228
rect 493468 5188 515956 5216
rect 493468 5176 493474 5188
rect 515950 5176 515956 5188
rect 516008 5176 516014 5228
rect 471330 5108 471336 5160
rect 471388 5148 471394 5160
rect 491110 5148 491116 5160
rect 471388 5120 491116 5148
rect 471388 5108 471394 5120
rect 491110 5108 491116 5120
rect 491168 5108 491174 5160
rect 497458 5108 497464 5160
rect 497516 5148 497522 5160
rect 519538 5148 519544 5160
rect 497516 5120 519544 5148
rect 497516 5108 497522 5120
rect 519538 5108 519544 5120
rect 519596 5108 519602 5160
rect 525058 5108 525064 5160
rect 525116 5148 525122 5160
rect 540790 5148 540796 5160
rect 525116 5120 540796 5148
rect 525116 5108 525122 5120
rect 540790 5108 540796 5120
rect 540848 5108 540854 5160
rect 477402 5040 477408 5092
rect 477460 5080 477466 5092
rect 498194 5080 498200 5092
rect 477460 5052 498200 5080
rect 477460 5040 477466 5052
rect 498194 5040 498200 5052
rect 498252 5040 498258 5092
rect 502242 5040 502248 5092
rect 502300 5080 502306 5092
rect 526622 5080 526628 5092
rect 502300 5052 526628 5080
rect 502300 5040 502306 5052
rect 526622 5040 526628 5052
rect 526680 5040 526686 5092
rect 529290 5040 529296 5092
rect 529348 5080 529354 5092
rect 551462 5080 551468 5092
rect 529348 5052 551468 5080
rect 529348 5040 529354 5052
rect 551462 5040 551468 5052
rect 551520 5040 551526 5092
rect 8110 4972 8116 5024
rect 8168 5012 8174 5024
rect 31754 5012 31760 5024
rect 8168 4984 31760 5012
rect 8168 4972 8174 4984
rect 31754 4972 31760 4984
rect 31812 4972 31818 5024
rect 486970 4972 486976 5024
rect 487028 5012 487034 5024
rect 508866 5012 508872 5024
rect 487028 4984 508872 5012
rect 487028 4972 487034 4984
rect 508866 4972 508872 4984
rect 508924 4972 508930 5024
rect 511902 4972 511908 5024
rect 511960 5012 511966 5024
rect 537202 5012 537208 5024
rect 511960 4984 537208 5012
rect 511960 4972 511966 4984
rect 537202 4972 537208 4984
rect 537260 4972 537266 5024
rect 8018 4904 8024 4956
rect 8076 4944 8082 4956
rect 33502 4944 33508 4956
rect 8076 4916 33508 4944
rect 8076 4904 8082 4916
rect 33502 4904 33508 4916
rect 33560 4904 33566 4956
rect 33594 4904 33600 4956
rect 33652 4944 33658 4956
rect 60826 4944 60832 4956
rect 33652 4916 60832 4944
rect 33652 4904 33658 4916
rect 60826 4904 60832 4916
rect 60884 4904 60890 4956
rect 467742 4904 467748 4956
rect 467800 4944 467806 4956
rect 487614 4944 487620 4956
rect 467800 4916 487620 4944
rect 467800 4904 467806 4916
rect 487614 4904 487620 4916
rect 487672 4904 487678 4956
rect 489822 4904 489828 4956
rect 489880 4944 489886 4956
rect 512454 4944 512460 4956
rect 489880 4916 512460 4944
rect 489880 4904 489886 4916
rect 512454 4904 512460 4916
rect 512512 4904 512518 4956
rect 518618 4904 518624 4956
rect 518676 4944 518682 4956
rect 544378 4944 544384 4956
rect 518676 4916 544384 4944
rect 518676 4904 518682 4916
rect 544378 4904 544384 4916
rect 544436 4904 544442 4956
rect 12342 4836 12348 4888
rect 12400 4876 12406 4888
rect 42978 4876 42984 4888
rect 12400 4848 42984 4876
rect 12400 4836 12406 4848
rect 42978 4836 42984 4848
rect 43036 4836 43042 4888
rect 482830 4836 482836 4888
rect 482888 4876 482894 4888
rect 505370 4876 505376 4888
rect 482888 4848 505376 4876
rect 482888 4836 482894 4848
rect 505370 4836 505376 4848
rect 505428 4836 505434 4888
rect 521562 4836 521568 4888
rect 521620 4876 521626 4888
rect 547874 4876 547880 4888
rect 521620 4848 547880 4876
rect 521620 4836 521626 4848
rect 547874 4836 547880 4848
rect 547932 4836 547938 4888
rect 556798 4836 556804 4888
rect 556856 4876 556862 4888
rect 576302 4876 576308 4888
rect 556856 4848 576308 4876
rect 556856 4836 556862 4848
rect 576302 4836 576308 4848
rect 576360 4836 576366 4888
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 34514 4808 34520 4820
rect 2924 4780 34520 4808
rect 2924 4768 2930 4780
rect 34514 4768 34520 4780
rect 34572 4768 34578 4820
rect 62114 4768 62120 4820
rect 62172 4808 62178 4820
rect 87322 4808 87328 4820
rect 62172 4780 87328 4808
rect 62172 4768 62178 4780
rect 87322 4768 87328 4780
rect 87380 4768 87386 4820
rect 480162 4768 480168 4820
rect 480220 4808 480226 4820
rect 501782 4808 501788 4820
rect 480220 4780 501788 4808
rect 480220 4768 480226 4780
rect 501782 4768 501788 4780
rect 501840 4768 501846 4820
rect 504910 4768 504916 4820
rect 504968 4808 504974 4820
rect 530118 4808 530124 4820
rect 504968 4780 530124 4808
rect 504968 4768 504974 4780
rect 530118 4768 530124 4780
rect 530176 4768 530182 4820
rect 533982 4768 533988 4820
rect 534040 4808 534046 4820
rect 562042 4808 562048 4820
rect 534040 4780 562048 4808
rect 534040 4768 534046 4780
rect 562042 4768 562048 4780
rect 562100 4768 562106 4820
rect 520918 4156 520924 4208
rect 520976 4196 520982 4208
rect 523034 4196 523040 4208
rect 520976 4168 523040 4196
rect 520976 4156 520982 4168
rect 523034 4156 523040 4168
rect 523092 4156 523098 4208
rect 314562 4088 314568 4140
rect 314620 4128 314626 4140
rect 316218 4128 316224 4140
rect 314620 4100 316224 4128
rect 314620 4088 314626 4100
rect 316218 4088 316224 4100
rect 316276 4088 316282 4140
rect 325602 4088 325608 4140
rect 325660 4128 325666 4140
rect 327994 4128 328000 4140
rect 325660 4100 328000 4128
rect 325660 4088 325666 4100
rect 327994 4088 328000 4100
rect 328052 4088 328058 4140
rect 342162 4088 342168 4140
rect 342220 4128 342226 4140
rect 346946 4128 346952 4140
rect 342220 4100 346952 4128
rect 342220 4088 342226 4100
rect 346946 4088 346952 4100
rect 347004 4088 347010 4140
rect 350442 4088 350448 4140
rect 350500 4128 350506 4140
rect 356330 4128 356336 4140
rect 350500 4100 356336 4128
rect 350500 4088 350506 4100
rect 356330 4088 356336 4100
rect 356388 4088 356394 4140
rect 358722 4088 358728 4140
rect 358780 4128 358786 4140
rect 365806 4128 365812 4140
rect 358780 4100 365812 4128
rect 358780 4088 358786 4100
rect 365806 4088 365812 4100
rect 365864 4088 365870 4140
rect 382182 4088 382188 4140
rect 382240 4128 382246 4140
rect 391842 4128 391848 4140
rect 382240 4100 391848 4128
rect 382240 4088 382246 4100
rect 391842 4088 391848 4100
rect 391900 4088 391906 4140
rect 397270 4088 397276 4140
rect 397328 4128 397334 4140
rect 408402 4128 408408 4140
rect 397328 4100 408408 4128
rect 397328 4088 397334 4100
rect 408402 4088 408408 4100
rect 408460 4088 408466 4140
rect 413922 4088 413928 4140
rect 413980 4128 413986 4140
rect 427262 4128 427268 4140
rect 413980 4100 427268 4128
rect 413980 4088 413986 4100
rect 427262 4088 427268 4100
rect 427320 4088 427326 4140
rect 430482 4088 430488 4140
rect 430540 4128 430546 4140
rect 446214 4128 446220 4140
rect 430540 4100 446220 4128
rect 430540 4088 430546 4100
rect 446214 4088 446220 4100
rect 446272 4088 446278 4140
rect 455322 4088 455328 4140
rect 455380 4128 455386 4140
rect 473446 4128 473452 4140
rect 455380 4100 473452 4128
rect 455380 4088 455386 4100
rect 473446 4088 473452 4100
rect 473504 4088 473510 4140
rect 481542 4088 481548 4140
rect 481600 4128 481606 4140
rect 502978 4128 502984 4140
rect 481600 4100 502984 4128
rect 481600 4088 481606 4100
rect 502978 4088 502984 4100
rect 503036 4088 503042 4140
rect 503622 4088 503628 4140
rect 503680 4128 503686 4140
rect 527818 4128 527824 4140
rect 503680 4100 527824 4128
rect 503680 4088 503686 4100
rect 527818 4088 527824 4100
rect 527876 4088 527882 4140
rect 538122 4088 538128 4140
rect 538180 4128 538186 4140
rect 566826 4128 566832 4140
rect 538180 4100 566832 4128
rect 538180 4088 538186 4100
rect 566826 4088 566832 4100
rect 566884 4088 566890 4140
rect 340782 4020 340788 4072
rect 340840 4060 340846 4072
rect 345750 4060 345756 4072
rect 340840 4032 345756 4060
rect 340840 4020 340846 4032
rect 345750 4020 345756 4032
rect 345808 4020 345814 4072
rect 375282 4020 375288 4072
rect 375340 4060 375346 4072
rect 383470 4060 383476 4072
rect 375340 4032 383476 4060
rect 375340 4020 375346 4032
rect 383470 4020 383476 4032
rect 383528 4020 383534 4072
rect 384850 4020 384856 4072
rect 384908 4060 384914 4072
rect 394234 4060 394240 4072
rect 384908 4032 394240 4060
rect 384908 4020 384914 4032
rect 394234 4020 394240 4032
rect 394292 4020 394298 4072
rect 394602 4020 394608 4072
rect 394660 4060 394666 4072
rect 406010 4060 406016 4072
rect 394660 4032 406016 4060
rect 394660 4020 394666 4032
rect 406010 4020 406016 4032
rect 406068 4020 406074 4072
rect 411162 4020 411168 4072
rect 411220 4060 411226 4072
rect 423766 4060 423772 4072
rect 411220 4032 423772 4060
rect 411220 4020 411226 4032
rect 423766 4020 423772 4032
rect 423824 4020 423830 4072
rect 424962 4020 424968 4072
rect 425020 4060 425026 4072
rect 439130 4060 439136 4072
rect 425020 4032 439136 4060
rect 425020 4020 425026 4032
rect 439130 4020 439136 4032
rect 439188 4020 439194 4072
rect 440142 4020 440148 4072
rect 440200 4060 440206 4072
rect 456886 4060 456892 4072
rect 440200 4032 456892 4060
rect 440200 4020 440206 4032
rect 456886 4020 456892 4032
rect 456944 4020 456950 4072
rect 460750 4020 460756 4072
rect 460808 4060 460814 4072
rect 479334 4060 479340 4072
rect 460808 4032 479340 4060
rect 460808 4020 460814 4032
rect 479334 4020 479340 4032
rect 479392 4020 479398 4072
rect 487062 4020 487068 4072
rect 487120 4060 487126 4072
rect 510062 4060 510068 4072
rect 487120 4032 510068 4060
rect 487120 4020 487126 4032
rect 510062 4020 510068 4032
rect 510120 4020 510126 4072
rect 513282 4020 513288 4072
rect 513340 4060 513346 4072
rect 538398 4060 538404 4072
rect 513340 4032 538404 4060
rect 513340 4020 513346 4032
rect 538398 4020 538404 4032
rect 538456 4020 538462 4072
rect 544930 4020 544936 4072
rect 544988 4060 544994 4072
rect 573910 4060 573916 4072
rect 544988 4032 573916 4060
rect 544988 4020 544994 4032
rect 573910 4020 573916 4032
rect 573968 4020 573974 4072
rect 333882 3952 333888 4004
rect 333940 3992 333946 4004
rect 337470 3992 337476 4004
rect 333940 3964 337476 3992
rect 333940 3952 333946 3964
rect 337470 3952 337476 3964
rect 337528 3952 337534 4004
rect 353202 3952 353208 4004
rect 353260 3992 353266 4004
rect 358722 3992 358728 4004
rect 353260 3964 358728 3992
rect 353260 3952 353266 3964
rect 358722 3952 358728 3964
rect 358780 3952 358786 4004
rect 369762 3952 369768 4004
rect 369820 3992 369826 4004
rect 377674 3992 377680 4004
rect 369820 3964 377680 3992
rect 369820 3952 369826 3964
rect 377674 3952 377680 3964
rect 377732 3952 377738 4004
rect 383562 3952 383568 4004
rect 383620 3992 383626 4004
rect 392946 3992 392952 4004
rect 383620 3964 392952 3992
rect 383620 3952 383626 3964
rect 392946 3952 392952 3964
rect 393004 3952 393010 4004
rect 393038 3952 393044 4004
rect 393096 3992 393102 4004
rect 403618 3992 403624 4004
rect 393096 3964 403624 3992
rect 393096 3952 393102 3964
rect 403618 3952 403624 3964
rect 403676 3952 403682 4004
rect 404262 3952 404268 4004
rect 404320 3992 404326 4004
rect 416682 3992 416688 4004
rect 404320 3964 416688 3992
rect 404320 3952 404326 3964
rect 416682 3952 416688 3964
rect 416740 3952 416746 4004
rect 418062 3952 418068 4004
rect 418120 3992 418126 4004
rect 432046 3992 432052 4004
rect 418120 3964 432052 3992
rect 418120 3952 418126 3964
rect 432046 3952 432052 3964
rect 432104 3952 432110 4004
rect 433058 3952 433064 4004
rect 433116 3992 433122 4004
rect 448606 3992 448612 4004
rect 433116 3964 448612 3992
rect 433116 3952 433122 3964
rect 448606 3952 448612 3964
rect 448664 3952 448670 4004
rect 451182 3952 451188 4004
rect 451240 3992 451246 4004
rect 469858 3992 469864 4004
rect 451240 3964 469864 3992
rect 451240 3952 451246 3964
rect 469858 3952 469864 3964
rect 469916 3952 469922 4004
rect 476022 3952 476028 4004
rect 476080 3992 476086 4004
rect 497090 3992 497096 4004
rect 476080 3964 497096 3992
rect 476080 3952 476086 3964
rect 497090 3952 497096 3964
rect 497148 3952 497154 4004
rect 506382 3952 506388 4004
rect 506440 3992 506446 4004
rect 531314 3992 531320 4004
rect 506440 3964 531320 3992
rect 506440 3952 506446 3964
rect 531314 3952 531320 3964
rect 531372 3952 531378 4004
rect 532510 3952 532516 4004
rect 532568 3992 532574 4004
rect 560846 3992 560852 4004
rect 532568 3964 560852 3992
rect 532568 3952 532574 3964
rect 560846 3952 560852 3964
rect 560904 3952 560910 4004
rect 373902 3884 373908 3936
rect 373960 3924 373966 3936
rect 382366 3924 382372 3936
rect 373960 3896 382372 3924
rect 373960 3884 373966 3896
rect 382366 3884 382372 3896
rect 382424 3884 382430 3936
rect 387702 3884 387708 3936
rect 387760 3924 387766 3936
rect 397730 3924 397736 3936
rect 387760 3896 397736 3924
rect 387760 3884 387766 3896
rect 397730 3884 397736 3896
rect 397788 3884 397794 3936
rect 398742 3884 398748 3936
rect 398800 3924 398806 3936
rect 410794 3924 410800 3936
rect 398800 3896 410800 3924
rect 398800 3884 398806 3896
rect 410794 3884 410800 3896
rect 410852 3884 410858 3936
rect 416590 3884 416596 3936
rect 416648 3924 416654 3936
rect 430850 3924 430856 3936
rect 416648 3896 430856 3924
rect 416648 3884 416654 3896
rect 430850 3884 430856 3896
rect 430908 3884 430914 3936
rect 436002 3884 436008 3936
rect 436060 3924 436066 3936
rect 452102 3924 452108 3936
rect 436060 3896 452108 3924
rect 436060 3884 436066 3896
rect 452102 3884 452108 3896
rect 452160 3884 452166 3936
rect 452562 3884 452568 3936
rect 452620 3924 452626 3936
rect 471054 3924 471060 3936
rect 452620 3896 471060 3924
rect 452620 3884 452626 3896
rect 471054 3884 471060 3896
rect 471112 3884 471118 3936
rect 478690 3884 478696 3936
rect 478748 3924 478754 3936
rect 500586 3924 500592 3936
rect 478748 3896 500592 3924
rect 478748 3884 478754 3896
rect 500586 3884 500592 3896
rect 500644 3884 500650 3936
rect 509142 3884 509148 3936
rect 509200 3924 509206 3936
rect 534902 3924 534908 3936
rect 509200 3896 534908 3924
rect 509200 3884 509206 3896
rect 534902 3884 534908 3896
rect 534960 3884 534966 3936
rect 542262 3884 542268 3936
rect 542320 3924 542326 3936
rect 571518 3924 571524 3936
rect 542320 3896 571524 3924
rect 542320 3884 542326 3896
rect 571518 3884 571524 3896
rect 571576 3884 571582 3936
rect 367002 3816 367008 3868
rect 367060 3856 367066 3868
rect 374086 3856 374092 3868
rect 367060 3828 374092 3856
rect 367060 3816 367066 3828
rect 374086 3816 374092 3828
rect 374144 3816 374150 3868
rect 376662 3816 376668 3868
rect 376720 3856 376726 3868
rect 385954 3856 385960 3868
rect 376720 3828 385960 3856
rect 376720 3816 376726 3828
rect 385954 3816 385960 3828
rect 386012 3816 386018 3868
rect 386322 3816 386328 3868
rect 386380 3856 386386 3868
rect 396534 3856 396540 3868
rect 386380 3828 396540 3856
rect 386380 3816 386386 3828
rect 396534 3816 396540 3828
rect 396592 3816 396598 3868
rect 397362 3816 397368 3868
rect 397420 3856 397426 3868
rect 397420 3828 400260 3856
rect 397420 3816 397426 3828
rect 344922 3748 344928 3800
rect 344980 3788 344986 3800
rect 350442 3788 350448 3800
rect 344980 3760 350448 3788
rect 344980 3748 344986 3760
rect 350442 3748 350448 3760
rect 350500 3748 350506 3800
rect 351822 3748 351828 3800
rect 351880 3788 351886 3800
rect 357526 3788 357532 3800
rect 351880 3760 357532 3788
rect 351880 3748 351886 3760
rect 357526 3748 357532 3760
rect 357584 3748 357590 3800
rect 361390 3748 361396 3800
rect 361448 3788 361454 3800
rect 368198 3788 368204 3800
rect 361448 3760 368204 3788
rect 361448 3748 361454 3760
rect 368198 3748 368204 3760
rect 368256 3748 368262 3800
rect 378042 3748 378048 3800
rect 378100 3788 378106 3800
rect 387150 3788 387156 3800
rect 378100 3760 387156 3788
rect 378100 3748 378106 3760
rect 387150 3748 387156 3760
rect 387208 3748 387214 3800
rect 389082 3748 389088 3800
rect 389140 3788 389146 3800
rect 389140 3760 399984 3788
rect 389140 3748 389146 3760
rect 354582 3680 354588 3732
rect 354640 3720 354646 3732
rect 361114 3720 361120 3732
rect 354640 3692 361120 3720
rect 354640 3680 354646 3692
rect 361114 3680 361120 3692
rect 361172 3680 361178 3732
rect 361482 3680 361488 3732
rect 361540 3720 361546 3732
rect 369394 3720 369400 3732
rect 361540 3692 369400 3720
rect 361540 3680 361546 3692
rect 369394 3680 369400 3692
rect 369452 3680 369458 3732
rect 372522 3680 372528 3732
rect 372580 3720 372586 3732
rect 381170 3720 381176 3732
rect 372580 3692 381176 3720
rect 372580 3680 372586 3692
rect 381170 3680 381176 3692
rect 381228 3680 381234 3732
rect 384942 3680 384948 3732
rect 385000 3720 385006 3732
rect 395338 3720 395344 3732
rect 385000 3692 395344 3720
rect 385000 3680 385006 3692
rect 395338 3680 395344 3692
rect 395396 3680 395402 3732
rect 399956 3720 399984 3760
rect 400122 3720 400128 3732
rect 399956 3692 400128 3720
rect 400122 3680 400128 3692
rect 400180 3680 400186 3732
rect 400232 3720 400260 3828
rect 402882 3816 402888 3868
rect 402940 3856 402946 3868
rect 415486 3856 415492 3868
rect 402940 3828 415492 3856
rect 402940 3816 402946 3828
rect 415486 3816 415492 3828
rect 415544 3816 415550 3868
rect 422202 3816 422208 3868
rect 422260 3856 422266 3868
rect 436738 3856 436744 3868
rect 422260 3828 436744 3856
rect 422260 3816 422266 3828
rect 436738 3816 436744 3828
rect 436796 3816 436802 3868
rect 437382 3816 437388 3868
rect 437440 3856 437446 3868
rect 453298 3856 453304 3868
rect 437440 3828 453304 3856
rect 437440 3816 437446 3828
rect 453298 3816 453304 3828
rect 453356 3816 453362 3868
rect 456610 3816 456616 3868
rect 456668 3856 456674 3868
rect 475746 3856 475752 3868
rect 456668 3828 475752 3856
rect 456668 3816 456674 3828
rect 475746 3816 475752 3828
rect 475804 3816 475810 3868
rect 491202 3816 491208 3868
rect 491260 3856 491266 3868
rect 513558 3856 513564 3868
rect 491260 3828 513564 3856
rect 491260 3816 491266 3828
rect 513558 3816 513564 3828
rect 513616 3816 513622 3868
rect 517422 3816 517428 3868
rect 517480 3856 517486 3868
rect 543182 3856 543188 3868
rect 517480 3828 543188 3856
rect 517480 3816 517486 3828
rect 543182 3816 543188 3828
rect 543240 3816 543246 3868
rect 545022 3816 545028 3868
rect 545080 3856 545086 3868
rect 575106 3856 575112 3868
rect 545080 3828 575112 3856
rect 545080 3816 545086 3828
rect 575106 3816 575112 3828
rect 575164 3816 575170 3868
rect 400306 3748 400312 3800
rect 400364 3788 400370 3800
rect 411898 3788 411904 3800
rect 400364 3760 411904 3788
rect 400364 3748 400370 3760
rect 411898 3748 411904 3760
rect 411956 3748 411962 3800
rect 412542 3748 412548 3800
rect 412600 3788 412606 3800
rect 426158 3788 426164 3800
rect 412600 3760 426164 3788
rect 412600 3748 412606 3760
rect 426158 3748 426164 3760
rect 426216 3748 426222 3800
rect 428918 3748 428924 3800
rect 428976 3788 428982 3800
rect 443822 3788 443828 3800
rect 428976 3760 443828 3788
rect 428976 3748 428982 3760
rect 443822 3748 443828 3760
rect 443880 3748 443886 3800
rect 444282 3748 444288 3800
rect 444340 3788 444346 3800
rect 461578 3788 461584 3800
rect 444340 3760 461584 3788
rect 444340 3748 444346 3760
rect 461578 3748 461584 3760
rect 461636 3748 461642 3800
rect 462222 3748 462228 3800
rect 462280 3788 462286 3800
rect 481726 3788 481732 3800
rect 462280 3760 481732 3788
rect 462280 3748 462286 3760
rect 481726 3748 481732 3760
rect 481784 3748 481790 3800
rect 492582 3748 492588 3800
rect 492640 3788 492646 3800
rect 514754 3788 514760 3800
rect 492640 3760 514760 3788
rect 492640 3748 492646 3760
rect 514754 3748 514760 3760
rect 514812 3748 514818 3800
rect 516042 3748 516048 3800
rect 516100 3788 516106 3800
rect 541986 3788 541992 3800
rect 516100 3760 541992 3788
rect 516100 3748 516106 3760
rect 541986 3748 541992 3760
rect 542044 3748 542050 3800
rect 549162 3748 549168 3800
rect 549220 3788 549226 3800
rect 578602 3788 578608 3800
rect 549220 3760 578608 3788
rect 549220 3748 549226 3760
rect 578602 3748 578608 3760
rect 578660 3748 578666 3800
rect 409598 3720 409604 3732
rect 400232 3692 409604 3720
rect 409598 3680 409604 3692
rect 409656 3680 409662 3732
rect 409782 3680 409788 3732
rect 409840 3720 409846 3732
rect 422570 3720 422576 3732
rect 409840 3692 422576 3720
rect 409840 3680 409846 3692
rect 422570 3680 422576 3692
rect 422628 3680 422634 3732
rect 423582 3680 423588 3732
rect 423640 3720 423646 3732
rect 437934 3720 437940 3732
rect 423640 3692 437940 3720
rect 423640 3680 423646 3692
rect 437934 3680 437940 3692
rect 437992 3680 437998 3732
rect 442810 3680 442816 3732
rect 442868 3720 442874 3732
rect 460382 3720 460388 3732
rect 442868 3692 460388 3720
rect 442868 3680 442874 3692
rect 460382 3680 460388 3692
rect 460440 3680 460446 3732
rect 466362 3680 466368 3732
rect 466420 3720 466426 3732
rect 486418 3720 486424 3732
rect 466420 3692 486424 3720
rect 466420 3680 466426 3692
rect 486418 3680 486424 3692
rect 486476 3680 486482 3732
rect 488442 3680 488448 3732
rect 488500 3720 488506 3732
rect 511258 3720 511264 3732
rect 488500 3692 511264 3720
rect 488500 3680 488506 3692
rect 511258 3680 511264 3692
rect 511316 3680 511322 3732
rect 514662 3680 514668 3732
rect 514720 3720 514726 3732
rect 539594 3720 539600 3732
rect 514720 3692 539600 3720
rect 514720 3680 514726 3692
rect 539594 3680 539600 3692
rect 539652 3680 539658 3732
rect 547782 3680 547788 3732
rect 547840 3720 547846 3732
rect 577406 3720 577412 3732
rect 547840 3692 577412 3720
rect 547840 3680 547846 3692
rect 577406 3680 577412 3692
rect 577464 3680 577470 3732
rect 324222 3612 324228 3664
rect 324280 3652 324286 3664
rect 326798 3652 326804 3664
rect 324280 3624 326804 3652
rect 324280 3612 324286 3624
rect 326798 3612 326804 3624
rect 326856 3612 326862 3664
rect 332502 3612 332508 3664
rect 332560 3652 332566 3664
rect 336274 3652 336280 3664
rect 332560 3624 336280 3652
rect 332560 3612 332566 3624
rect 336274 3612 336280 3624
rect 336332 3612 336338 3664
rect 357342 3612 357348 3664
rect 357400 3652 357406 3664
rect 364610 3652 364616 3664
rect 357400 3624 364616 3652
rect 357400 3612 357406 3624
rect 364610 3612 364616 3624
rect 364668 3612 364674 3664
rect 370958 3612 370964 3664
rect 371016 3652 371022 3664
rect 378870 3652 378876 3664
rect 371016 3624 378876 3652
rect 371016 3612 371022 3624
rect 378870 3612 378876 3624
rect 378928 3612 378934 3664
rect 379238 3612 379244 3664
rect 379296 3652 379302 3664
rect 388254 3652 388260 3664
rect 379296 3624 388260 3652
rect 379296 3612 379302 3624
rect 388254 3612 388260 3624
rect 388312 3612 388318 3664
rect 393222 3612 393228 3664
rect 393280 3652 393286 3664
rect 404814 3652 404820 3664
rect 393280 3624 404820 3652
rect 393280 3612 393286 3624
rect 404814 3612 404820 3624
rect 404872 3612 404878 3664
rect 407022 3612 407028 3664
rect 407080 3652 407086 3664
rect 420178 3652 420184 3664
rect 407080 3624 420184 3652
rect 407080 3612 407086 3624
rect 420178 3612 420184 3624
rect 420236 3612 420242 3664
rect 420730 3612 420736 3664
rect 420788 3652 420794 3664
rect 435542 3652 435548 3664
rect 420788 3624 435548 3652
rect 420788 3612 420794 3624
rect 435542 3612 435548 3624
rect 435600 3612 435606 3664
rect 438670 3612 438676 3664
rect 438728 3652 438734 3664
rect 455690 3652 455696 3664
rect 438728 3624 455696 3652
rect 438728 3612 438734 3624
rect 455690 3612 455696 3624
rect 455748 3612 455754 3664
rect 460842 3612 460848 3664
rect 460900 3652 460906 3664
rect 480530 3652 480536 3664
rect 460900 3624 480536 3652
rect 460900 3612 460906 3624
rect 480530 3612 480536 3624
rect 480588 3612 480594 3664
rect 484302 3612 484308 3664
rect 484360 3652 484366 3664
rect 506474 3652 506480 3664
rect 484360 3624 506480 3652
rect 484360 3612 484366 3624
rect 506474 3612 506480 3624
rect 506532 3612 506538 3664
rect 510522 3612 510528 3664
rect 510580 3652 510586 3664
rect 536098 3652 536104 3664
rect 510580 3624 536104 3652
rect 510580 3612 510586 3624
rect 536098 3612 536104 3624
rect 536156 3612 536162 3664
rect 540882 3612 540888 3664
rect 540940 3652 540946 3664
rect 570322 3652 570328 3664
rect 540940 3624 570328 3652
rect 540940 3612 540946 3624
rect 570322 3612 570328 3624
rect 570380 3612 570386 3664
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28810 3584 28816 3596
rect 27764 3556 28816 3584
rect 27764 3544 27770 3556
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 51718 3584 51724 3596
rect 45526 3556 51724 3584
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12250 3516 12256 3528
rect 11204 3488 12256 3516
rect 11204 3476 11210 3488
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 26142 3516 26148 3528
rect 25372 3488 26148 3516
rect 25372 3476 25378 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 45526 3516 45554 3556
rect 51718 3544 51724 3556
rect 51776 3544 51782 3596
rect 62206 3584 62212 3596
rect 55186 3556 62212 3584
rect 33152 3488 45554 3516
rect 26510 3408 26516 3460
rect 26568 3448 26574 3460
rect 33152 3448 33180 3488
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 52362 3516 52368 3528
rect 51408 3488 52368 3516
rect 51408 3476 51414 3488
rect 52362 3476 52368 3488
rect 52420 3476 52426 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 53650 3516 53656 3528
rect 52604 3488 53656 3516
rect 52604 3476 52610 3488
rect 53650 3476 53656 3488
rect 53708 3476 53714 3528
rect 26568 3420 33180 3448
rect 26568 3408 26574 3420
rect 34790 3408 34796 3460
rect 34848 3448 34854 3460
rect 35802 3448 35808 3460
rect 34848 3420 35808 3448
rect 34848 3408 34854 3420
rect 35802 3408 35808 3420
rect 35860 3408 35866 3460
rect 35986 3408 35992 3460
rect 36044 3448 36050 3460
rect 37182 3448 37188 3460
rect 36044 3420 37188 3448
rect 36044 3408 36050 3420
rect 37182 3408 37188 3420
rect 37240 3408 37246 3460
rect 40678 3408 40684 3460
rect 40736 3448 40742 3460
rect 41322 3448 41328 3460
rect 40736 3420 41328 3448
rect 40736 3408 40742 3420
rect 41322 3408 41328 3420
rect 41380 3408 41386 3460
rect 41874 3408 41880 3460
rect 41932 3448 41938 3460
rect 42702 3448 42708 3460
rect 41932 3420 42708 3448
rect 41932 3408 41938 3420
rect 42702 3408 42708 3420
rect 42760 3408 42766 3460
rect 43070 3408 43076 3460
rect 43128 3448 43134 3460
rect 44082 3448 44088 3460
rect 43128 3420 44088 3448
rect 43128 3408 43134 3420
rect 44082 3408 44088 3420
rect 44140 3408 44146 3460
rect 44266 3408 44272 3460
rect 44324 3448 44330 3460
rect 45370 3448 45376 3460
rect 44324 3420 45376 3448
rect 44324 3408 44330 3420
rect 45370 3408 45376 3420
rect 45428 3408 45434 3460
rect 48958 3408 48964 3460
rect 49016 3448 49022 3460
rect 49602 3448 49608 3460
rect 49016 3420 49608 3448
rect 49016 3408 49022 3420
rect 49602 3408 49608 3420
rect 49660 3408 49666 3460
rect 19426 3272 19432 3324
rect 19484 3312 19490 3324
rect 20530 3312 20536 3324
rect 19484 3284 20536 3312
rect 19484 3272 19490 3284
rect 20530 3272 20536 3284
rect 20588 3272 20594 3324
rect 37182 3272 37188 3324
rect 37240 3312 37246 3324
rect 55186 3312 55214 3556
rect 62206 3544 62212 3556
rect 62264 3544 62270 3596
rect 77386 3544 77392 3596
rect 77444 3584 77450 3596
rect 78490 3584 78496 3596
rect 77444 3556 78496 3584
rect 77444 3544 77450 3556
rect 78490 3544 78496 3556
rect 78548 3544 78554 3596
rect 307754 3544 307760 3596
rect 307812 3584 307818 3596
rect 309042 3584 309048 3596
rect 307812 3556 309048 3584
rect 307812 3544 307818 3556
rect 309042 3544 309048 3556
rect 309100 3544 309106 3596
rect 326982 3544 326988 3596
rect 327040 3584 327046 3596
rect 330386 3584 330392 3596
rect 327040 3556 330392 3584
rect 327040 3544 327046 3556
rect 330386 3544 330392 3556
rect 330444 3544 330450 3596
rect 335262 3544 335268 3596
rect 335320 3584 335326 3596
rect 339862 3584 339868 3596
rect 335320 3556 339868 3584
rect 335320 3544 335326 3556
rect 339862 3544 339868 3556
rect 339920 3544 339926 3596
rect 353110 3544 353116 3596
rect 353168 3584 353174 3596
rect 359918 3584 359924 3596
rect 353168 3556 359924 3584
rect 353168 3544 353174 3556
rect 359918 3544 359924 3556
rect 359976 3544 359982 3596
rect 362862 3544 362868 3596
rect 362920 3584 362926 3596
rect 370590 3584 370596 3596
rect 362920 3556 370596 3584
rect 362920 3544 362926 3556
rect 370590 3544 370596 3556
rect 370648 3544 370654 3596
rect 371142 3544 371148 3596
rect 371200 3584 371206 3596
rect 379974 3584 379980 3596
rect 371200 3556 379980 3584
rect 371200 3544 371206 3556
rect 379974 3544 379980 3556
rect 380032 3544 380038 3596
rect 380802 3544 380808 3596
rect 380860 3584 380866 3596
rect 390646 3584 390652 3596
rect 380860 3556 390652 3584
rect 380860 3544 380866 3556
rect 390646 3544 390652 3556
rect 390704 3544 390710 3596
rect 401502 3544 401508 3596
rect 401560 3584 401566 3596
rect 413094 3584 413100 3596
rect 401560 3556 413100 3584
rect 401560 3544 401566 3556
rect 413094 3544 413100 3556
rect 413152 3544 413158 3596
rect 415210 3544 415216 3596
rect 415268 3584 415274 3596
rect 429654 3584 429660 3596
rect 415268 3556 429660 3584
rect 415268 3544 415274 3556
rect 429654 3544 429660 3556
rect 429712 3544 429718 3596
rect 433150 3544 433156 3596
rect 433208 3584 433214 3596
rect 449802 3584 449808 3596
rect 433208 3556 449808 3584
rect 433208 3544 433214 3556
rect 449802 3544 449808 3556
rect 449860 3544 449866 3596
rect 451090 3544 451096 3596
rect 451148 3584 451154 3596
rect 468662 3584 468668 3596
rect 451148 3556 468668 3584
rect 451148 3544 451154 3556
rect 468662 3544 468668 3556
rect 468720 3544 468726 3596
rect 469030 3544 469036 3596
rect 469088 3584 469094 3596
rect 488810 3584 488816 3596
rect 469088 3556 488816 3584
rect 469088 3544 469094 3556
rect 488810 3544 488816 3556
rect 488868 3544 488874 3596
rect 495342 3544 495348 3596
rect 495400 3584 495406 3596
rect 518342 3584 518348 3596
rect 495400 3556 518348 3584
rect 495400 3544 495406 3556
rect 518342 3544 518348 3556
rect 518400 3544 518406 3596
rect 518802 3544 518808 3596
rect 518860 3584 518866 3596
rect 545482 3584 545488 3596
rect 518860 3556 545488 3584
rect 518860 3544 518866 3556
rect 545482 3544 545488 3556
rect 545540 3544 545546 3596
rect 550542 3544 550548 3596
rect 550600 3584 550606 3596
rect 582190 3584 582196 3596
rect 550600 3556 582196 3584
rect 550600 3544 550606 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 56502 3516 56508 3528
rect 56100 3488 56508 3516
rect 56100 3476 56106 3488
rect 56502 3476 56508 3488
rect 56560 3476 56566 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 60826 3476 60832 3528
rect 60884 3516 60890 3528
rect 62022 3516 62028 3528
rect 60884 3488 62028 3516
rect 60884 3476 60890 3488
rect 62022 3476 62028 3488
rect 62080 3476 62086 3528
rect 64322 3476 64328 3528
rect 64380 3516 64386 3528
rect 64782 3516 64788 3528
rect 64380 3488 64788 3516
rect 64380 3476 64386 3488
rect 64782 3476 64788 3488
rect 64840 3476 64846 3528
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 66714 3476 66720 3528
rect 66772 3516 66778 3528
rect 67542 3516 67548 3528
rect 66772 3488 67548 3516
rect 66772 3476 66778 3488
rect 67542 3476 67548 3488
rect 67600 3476 67606 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 82078 3476 82084 3528
rect 82136 3516 82142 3528
rect 82722 3516 82728 3528
rect 82136 3488 82728 3516
rect 82136 3476 82142 3488
rect 82722 3476 82728 3488
rect 82780 3476 82786 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 84102 3516 84108 3528
rect 83332 3488 84108 3516
rect 83332 3476 83338 3488
rect 84102 3476 84108 3488
rect 84160 3476 84166 3528
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 85482 3516 85488 3528
rect 84528 3488 85488 3516
rect 84528 3476 84534 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 92382 3516 92388 3528
rect 91612 3488 92388 3516
rect 91612 3476 91618 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 106182 3516 106188 3528
rect 105780 3488 106188 3516
rect 105780 3476 105786 3488
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 110322 3516 110328 3528
rect 109368 3488 110328 3516
rect 109368 3476 109374 3488
rect 110322 3476 110328 3488
rect 110380 3476 110386 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111518 3516 111524 3528
rect 110564 3488 111524 3516
rect 110564 3476 110570 3488
rect 111518 3476 111524 3488
rect 111576 3476 111582 3528
rect 114002 3476 114008 3528
rect 114060 3516 114066 3528
rect 114462 3516 114468 3528
rect 114060 3488 114468 3516
rect 114060 3476 114066 3488
rect 114462 3476 114468 3488
rect 114520 3476 114526 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 116394 3476 116400 3528
rect 116452 3516 116458 3528
rect 117222 3516 117228 3528
rect 116452 3488 117228 3516
rect 116452 3476 116458 3488
rect 117222 3476 117228 3488
rect 117280 3476 117286 3528
rect 117590 3476 117596 3528
rect 117648 3516 117654 3528
rect 118602 3516 118608 3528
rect 117648 3488 118608 3516
rect 117648 3476 117654 3488
rect 118602 3476 118608 3488
rect 118660 3476 118666 3528
rect 122282 3476 122288 3528
rect 122340 3516 122346 3528
rect 122742 3516 122748 3528
rect 122340 3488 122748 3516
rect 122340 3476 122346 3488
rect 122742 3476 122748 3488
rect 122800 3476 122806 3528
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126882 3516 126888 3528
rect 125928 3488 126888 3516
rect 125928 3476 125934 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128262 3516 128268 3528
rect 127032 3488 128268 3516
rect 127032 3476 127038 3488
rect 128262 3476 128268 3488
rect 128320 3476 128326 3528
rect 130562 3476 130568 3528
rect 130620 3516 130626 3528
rect 131022 3516 131028 3528
rect 130620 3488 131028 3516
rect 130620 3476 130626 3488
rect 131022 3476 131028 3488
rect 131080 3476 131086 3528
rect 132954 3476 132960 3528
rect 133012 3516 133018 3528
rect 133782 3516 133788 3528
rect 133012 3488 133788 3516
rect 133012 3476 133018 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
rect 134150 3476 134156 3528
rect 134208 3516 134214 3528
rect 135162 3516 135168 3528
rect 134208 3488 135168 3516
rect 134208 3476 134214 3488
rect 135162 3476 135168 3488
rect 135220 3476 135226 3528
rect 138842 3476 138848 3528
rect 138900 3516 138906 3528
rect 139302 3516 139308 3528
rect 138900 3488 139308 3516
rect 138900 3476 138906 3488
rect 139302 3476 139308 3488
rect 139360 3476 139366 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 140682 3516 140688 3528
rect 140096 3488 140688 3516
rect 140096 3476 140102 3488
rect 140682 3476 140688 3488
rect 140740 3476 140746 3528
rect 141234 3476 141240 3528
rect 141292 3516 141298 3528
rect 142062 3516 142068 3528
rect 141292 3488 142068 3516
rect 141292 3476 141298 3488
rect 142062 3476 142068 3488
rect 142120 3476 142126 3528
rect 142430 3476 142436 3528
rect 142488 3516 142494 3528
rect 143442 3516 143448 3528
rect 142488 3488 143448 3516
rect 142488 3476 142494 3488
rect 143442 3476 143448 3488
rect 143500 3476 143506 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
rect 150342 3516 150348 3528
rect 149572 3488 150348 3516
rect 149572 3476 149578 3488
rect 150342 3476 150348 3488
rect 150400 3476 150406 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 153102 3516 153108 3528
rect 151872 3488 153108 3516
rect 151872 3476 151878 3488
rect 153102 3476 153108 3488
rect 153160 3476 153166 3528
rect 156598 3476 156604 3528
rect 156656 3516 156662 3528
rect 157242 3516 157248 3528
rect 156656 3488 157248 3516
rect 156656 3476 156662 3488
rect 157242 3476 157248 3488
rect 157300 3476 157306 3528
rect 157794 3476 157800 3528
rect 157852 3516 157858 3528
rect 158622 3516 158628 3528
rect 157852 3488 158628 3516
rect 157852 3476 157858 3488
rect 158622 3476 158628 3488
rect 158680 3476 158686 3528
rect 158898 3476 158904 3528
rect 158956 3516 158962 3528
rect 160002 3516 160008 3528
rect 158956 3488 160008 3516
rect 158956 3476 158962 3488
rect 160002 3476 160008 3488
rect 160060 3476 160066 3528
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161382 3516 161388 3528
rect 160152 3488 161388 3516
rect 160152 3476 160158 3488
rect 161382 3476 161388 3488
rect 161440 3476 161446 3528
rect 163682 3476 163688 3528
rect 163740 3516 163746 3528
rect 164142 3516 164148 3528
rect 163740 3488 164148 3516
rect 163740 3476 163746 3488
rect 164142 3476 164148 3488
rect 164200 3476 164206 3528
rect 164878 3476 164884 3528
rect 164936 3516 164942 3528
rect 165522 3516 165528 3528
rect 164936 3488 165528 3516
rect 164936 3476 164942 3488
rect 165522 3476 165528 3488
rect 165580 3476 165586 3528
rect 166074 3476 166080 3528
rect 166132 3516 166138 3528
rect 166902 3516 166908 3528
rect 166132 3488 166908 3516
rect 166132 3476 166138 3488
rect 166902 3476 166908 3488
rect 166960 3476 166966 3528
rect 167178 3476 167184 3528
rect 167236 3516 167242 3528
rect 168282 3516 168288 3528
rect 167236 3488 168288 3516
rect 167236 3476 167242 3488
rect 168282 3476 168288 3488
rect 168340 3476 168346 3528
rect 171962 3476 171968 3528
rect 172020 3516 172026 3528
rect 172422 3516 172428 3528
rect 172020 3488 172428 3516
rect 172020 3476 172026 3488
rect 172422 3476 172428 3488
rect 172480 3476 172486 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173802 3516 173808 3528
rect 173216 3488 173808 3516
rect 173216 3476 173222 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 174262 3476 174268 3528
rect 174320 3516 174326 3528
rect 175182 3516 175188 3528
rect 174320 3488 175188 3516
rect 174320 3476 174326 3488
rect 175182 3476 175188 3488
rect 175240 3476 175246 3528
rect 175458 3476 175464 3528
rect 175516 3516 175522 3528
rect 176562 3516 176568 3528
rect 175516 3488 176568 3516
rect 175516 3476 175522 3488
rect 176562 3476 176568 3488
rect 176620 3476 176626 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177758 3516 177764 3528
rect 176712 3488 177764 3516
rect 176712 3476 176718 3488
rect 177758 3476 177764 3488
rect 177816 3476 177822 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180702 3516 180708 3528
rect 180300 3488 180708 3516
rect 180300 3476 180306 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 181438 3476 181444 3528
rect 181496 3516 181502 3528
rect 182082 3516 182088 3528
rect 181496 3488 182088 3516
rect 181496 3476 181502 3488
rect 182082 3476 182088 3488
rect 182140 3476 182146 3528
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 184934 3476 184940 3528
rect 184992 3516 184998 3528
rect 186222 3516 186228 3528
rect 184992 3488 186228 3516
rect 184992 3476 184998 3488
rect 186222 3476 186228 3488
rect 186280 3476 186286 3528
rect 188522 3476 188528 3528
rect 188580 3516 188586 3528
rect 188982 3516 188988 3528
rect 188580 3488 188988 3516
rect 188580 3476 188586 3488
rect 188982 3476 188988 3488
rect 189040 3476 189046 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 191742 3516 191748 3528
rect 190880 3488 191748 3516
rect 190880 3476 190886 3488
rect 191742 3476 191748 3488
rect 191800 3476 191806 3528
rect 192018 3476 192024 3528
rect 192076 3516 192082 3528
rect 193122 3516 193128 3528
rect 192076 3488 193128 3516
rect 192076 3476 192082 3488
rect 193122 3476 193128 3488
rect 193180 3476 193186 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194318 3516 194324 3528
rect 193272 3488 194324 3516
rect 193272 3476 193278 3488
rect 194318 3476 194324 3488
rect 194376 3476 194382 3528
rect 197906 3476 197912 3528
rect 197964 3516 197970 3528
rect 198642 3516 198648 3528
rect 197964 3488 198648 3516
rect 197964 3476 197970 3488
rect 198642 3476 198648 3488
rect 198700 3476 198706 3528
rect 199102 3476 199108 3528
rect 199160 3516 199166 3528
rect 200022 3516 200028 3528
rect 199160 3488 200028 3516
rect 199160 3476 199166 3488
rect 200022 3476 200028 3488
rect 200080 3476 200086 3528
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 202782 3516 202788 3528
rect 201552 3488 202788 3516
rect 201552 3476 201558 3488
rect 202782 3476 202788 3488
rect 202840 3476 202846 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 205542 3516 205548 3528
rect 205140 3488 205548 3516
rect 205140 3476 205146 3488
rect 205542 3476 205548 3488
rect 205600 3476 205606 3528
rect 206186 3476 206192 3528
rect 206244 3516 206250 3528
rect 206922 3516 206928 3528
rect 206244 3488 206928 3516
rect 206244 3476 206250 3488
rect 206922 3476 206928 3488
rect 206980 3476 206986 3528
rect 207382 3476 207388 3528
rect 207440 3516 207446 3528
rect 208302 3516 208308 3528
rect 207440 3488 208308 3516
rect 207440 3476 207446 3488
rect 208302 3476 208308 3488
rect 208360 3476 208366 3528
rect 209774 3476 209780 3528
rect 209832 3516 209838 3528
rect 210878 3516 210884 3528
rect 209832 3488 210884 3516
rect 209832 3476 209838 3488
rect 210878 3476 210884 3488
rect 210936 3476 210942 3528
rect 213362 3476 213368 3528
rect 213420 3516 213426 3528
rect 213822 3516 213828 3528
rect 213420 3488 213828 3516
rect 213420 3476 213426 3488
rect 213822 3476 213828 3488
rect 213880 3476 213886 3528
rect 214466 3476 214472 3528
rect 214524 3516 214530 3528
rect 215202 3516 215208 3528
rect 214524 3488 215208 3516
rect 214524 3476 214530 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 216582 3516 216588 3528
rect 215720 3488 216588 3516
rect 215720 3476 215726 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 216858 3476 216864 3528
rect 216916 3516 216922 3528
rect 217962 3516 217968 3528
rect 216916 3488 217968 3516
rect 216916 3476 216922 3488
rect 217962 3476 217968 3488
rect 218020 3476 218026 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 219158 3516 219164 3528
rect 218112 3488 219164 3516
rect 218112 3476 218118 3488
rect 219158 3476 219164 3488
rect 219216 3476 219222 3528
rect 222746 3476 222752 3528
rect 222804 3516 222810 3528
rect 223482 3516 223488 3528
rect 222804 3488 223488 3516
rect 222804 3476 222810 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 224862 3516 224868 3528
rect 224000 3488 224868 3516
rect 224000 3476 224006 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 229830 3476 229836 3528
rect 229888 3516 229894 3528
rect 230382 3516 230388 3528
rect 229888 3488 230388 3516
rect 229888 3476 229894 3488
rect 230382 3476 230388 3488
rect 230440 3476 230446 3528
rect 231026 3476 231032 3528
rect 231084 3516 231090 3528
rect 231762 3516 231768 3528
rect 231084 3488 231768 3516
rect 231084 3476 231090 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 234614 3476 234620 3528
rect 234672 3516 234678 3528
rect 235902 3516 235908 3528
rect 234672 3488 235908 3516
rect 234672 3476 234678 3488
rect 235902 3476 235908 3488
rect 235960 3476 235966 3528
rect 238110 3476 238116 3528
rect 238168 3516 238174 3528
rect 238662 3516 238668 3528
rect 238168 3488 238668 3516
rect 238168 3476 238174 3488
rect 238662 3476 238668 3488
rect 238720 3476 238726 3528
rect 239306 3476 239312 3528
rect 239364 3516 239370 3528
rect 240042 3516 240048 3528
rect 239364 3488 240048 3516
rect 239364 3476 239370 3488
rect 240042 3476 240048 3488
rect 240100 3476 240106 3528
rect 240502 3476 240508 3528
rect 240560 3516 240566 3528
rect 241422 3516 241428 3528
rect 240560 3488 241428 3516
rect 240560 3476 240566 3488
rect 241422 3476 241428 3488
rect 241480 3476 241486 3528
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 243998 3516 244004 3528
rect 242952 3488 244004 3516
rect 242952 3476 242958 3488
rect 243998 3476 244004 3488
rect 244056 3476 244062 3528
rect 247586 3476 247592 3528
rect 247644 3516 247650 3528
rect 248322 3516 248328 3528
rect 247644 3488 248328 3516
rect 247644 3476 247650 3488
rect 248322 3476 248328 3488
rect 248380 3476 248386 3528
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 251082 3516 251088 3528
rect 250036 3488 251088 3516
rect 250036 3476 250042 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 251174 3476 251180 3528
rect 251232 3516 251238 3528
rect 252462 3516 252468 3528
rect 251232 3488 252468 3516
rect 251232 3476 251238 3488
rect 252462 3476 252468 3488
rect 252520 3476 252526 3528
rect 254670 3476 254676 3528
rect 254728 3516 254734 3528
rect 255222 3516 255228 3528
rect 254728 3488 255228 3516
rect 254728 3476 254734 3488
rect 255222 3476 255228 3488
rect 255280 3476 255286 3528
rect 255866 3476 255872 3528
rect 255924 3516 255930 3528
rect 256602 3516 256608 3528
rect 255924 3488 256608 3516
rect 255924 3476 255930 3488
rect 256602 3476 256608 3488
rect 256660 3476 256666 3528
rect 257062 3476 257068 3528
rect 257120 3516 257126 3528
rect 257982 3516 257988 3528
rect 257120 3488 257988 3516
rect 257120 3476 257126 3488
rect 257982 3476 257988 3488
rect 258040 3476 258046 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 264882 3516 264888 3528
rect 264204 3488 264888 3516
rect 264204 3476 264210 3488
rect 264882 3476 264888 3488
rect 264940 3476 264946 3528
rect 265342 3476 265348 3528
rect 265400 3516 265406 3528
rect 266262 3516 266268 3528
rect 265400 3488 266268 3516
rect 265400 3476 265406 3488
rect 266262 3476 266268 3488
rect 266320 3476 266326 3528
rect 266538 3476 266544 3528
rect 266596 3516 266602 3528
rect 267550 3516 267556 3528
rect 266596 3488 267556 3516
rect 266596 3476 266602 3488
rect 267550 3476 267556 3488
rect 267608 3476 267614 3528
rect 267734 3476 267740 3528
rect 267792 3516 267798 3528
rect 269022 3516 269028 3528
rect 267792 3488 269028 3516
rect 267792 3476 267798 3488
rect 269022 3476 269028 3488
rect 269080 3476 269086 3528
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 274542 3516 274548 3528
rect 273680 3488 274548 3516
rect 273680 3476 273686 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 276014 3476 276020 3528
rect 276072 3516 276078 3528
rect 277302 3516 277308 3528
rect 276072 3488 277308 3516
rect 276072 3476 276078 3488
rect 277302 3476 277308 3488
rect 277360 3476 277366 3528
rect 280706 3476 280712 3528
rect 280764 3516 280770 3528
rect 281442 3516 281448 3528
rect 280764 3488 281448 3516
rect 280764 3476 280770 3488
rect 281442 3476 281448 3488
rect 281500 3476 281506 3528
rect 281902 3476 281908 3528
rect 281960 3516 281966 3528
rect 282822 3516 282828 3528
rect 281960 3488 282828 3516
rect 281960 3476 281966 3488
rect 282822 3476 282828 3488
rect 282880 3476 282886 3528
rect 283098 3476 283104 3528
rect 283156 3516 283162 3528
rect 284570 3516 284576 3528
rect 283156 3488 284576 3516
rect 283156 3476 283162 3488
rect 284570 3476 284576 3488
rect 284628 3476 284634 3528
rect 285398 3476 285404 3528
rect 285456 3516 285462 3528
rect 286594 3516 286600 3528
rect 285456 3488 286600 3516
rect 285456 3476 285462 3488
rect 286594 3476 286600 3488
rect 286652 3476 286658 3528
rect 288986 3476 288992 3528
rect 289044 3516 289050 3528
rect 289722 3516 289728 3528
rect 289044 3488 289728 3516
rect 289044 3476 289050 3488
rect 289722 3476 289728 3488
rect 289780 3476 289786 3528
rect 291378 3476 291384 3528
rect 291436 3516 291442 3528
rect 291930 3516 291936 3528
rect 291436 3488 291936 3516
rect 291436 3476 291442 3488
rect 291930 3476 291936 3488
rect 291988 3476 291994 3528
rect 301406 3476 301412 3528
rect 301464 3516 301470 3528
rect 301958 3516 301964 3528
rect 301464 3488 301964 3516
rect 301464 3476 301470 3488
rect 301958 3476 301964 3488
rect 302016 3476 302022 3528
rect 303522 3476 303528 3528
rect 303580 3516 303586 3528
rect 304350 3516 304356 3528
rect 303580 3488 304356 3516
rect 303580 3476 303586 3488
rect 304350 3476 304356 3488
rect 304408 3476 304414 3528
rect 304902 3476 304908 3528
rect 304960 3516 304966 3528
rect 305546 3516 305552 3528
rect 304960 3488 305552 3516
rect 304960 3476 304966 3488
rect 305546 3476 305552 3488
rect 305604 3476 305610 3528
rect 310422 3476 310428 3528
rect 310480 3516 310486 3528
rect 311434 3516 311440 3528
rect 310480 3488 311440 3516
rect 310480 3476 310486 3488
rect 311434 3476 311440 3488
rect 311492 3476 311498 3528
rect 311802 3476 311808 3528
rect 311860 3516 311866 3528
rect 312630 3516 312636 3528
rect 311860 3488 312636 3516
rect 311860 3476 311866 3488
rect 312630 3476 312636 3488
rect 312688 3476 312694 3528
rect 318702 3476 318708 3528
rect 318760 3516 318766 3528
rect 320910 3516 320916 3528
rect 318760 3488 320916 3516
rect 318760 3476 318766 3488
rect 320910 3476 320916 3488
rect 320968 3476 320974 3528
rect 321278 3476 321284 3528
rect 321336 3516 321342 3528
rect 323302 3516 323308 3528
rect 321336 3488 323308 3516
rect 321336 3476 321342 3488
rect 323302 3476 323308 3488
rect 323360 3476 323366 3528
rect 327718 3476 327724 3528
rect 327776 3516 327782 3528
rect 329190 3516 329196 3528
rect 327776 3488 329196 3516
rect 327776 3476 327782 3488
rect 329190 3476 329196 3488
rect 329248 3476 329254 3528
rect 331122 3476 331128 3528
rect 331180 3516 331186 3528
rect 333882 3516 333888 3528
rect 331180 3488 333888 3516
rect 331180 3476 331186 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 335078 3476 335084 3528
rect 335136 3516 335142 3528
rect 338666 3516 338672 3528
rect 335136 3488 338672 3516
rect 335136 3476 335142 3488
rect 338666 3476 338672 3488
rect 338724 3476 338730 3528
rect 339402 3476 339408 3528
rect 339460 3516 339466 3528
rect 344554 3516 344560 3528
rect 339460 3488 344560 3516
rect 339460 3476 339466 3488
rect 344554 3476 344560 3488
rect 344612 3476 344618 3528
rect 344830 3476 344836 3528
rect 344888 3516 344894 3528
rect 349246 3516 349252 3528
rect 344888 3488 349252 3516
rect 344888 3476 344894 3488
rect 349246 3476 349252 3488
rect 349304 3476 349310 3528
rect 357250 3476 357256 3528
rect 357308 3516 357314 3528
rect 363506 3516 363512 3528
rect 357308 3488 363512 3516
rect 357308 3476 357314 3488
rect 363506 3476 363512 3488
rect 363564 3476 363570 3528
rect 364242 3476 364248 3528
rect 364300 3516 364306 3528
rect 371694 3516 371700 3528
rect 364300 3488 371700 3516
rect 364300 3476 364306 3488
rect 371694 3476 371700 3488
rect 371752 3476 371758 3528
rect 375190 3476 375196 3528
rect 375248 3516 375254 3528
rect 384758 3516 384764 3528
rect 375248 3488 384764 3516
rect 375248 3476 375254 3488
rect 384758 3476 384764 3488
rect 384816 3476 384822 3528
rect 388898 3476 388904 3528
rect 388956 3516 388962 3528
rect 398926 3516 398932 3528
rect 388956 3488 398932 3516
rect 388956 3476 388962 3488
rect 398926 3476 398932 3488
rect 398984 3476 398990 3528
rect 402790 3476 402796 3528
rect 402848 3516 402854 3528
rect 414290 3516 414296 3528
rect 402848 3488 414296 3516
rect 402848 3476 402854 3488
rect 414290 3476 414296 3488
rect 414348 3476 414354 3528
rect 415118 3476 415124 3528
rect 415176 3516 415182 3528
rect 428458 3516 428464 3528
rect 415176 3488 428464 3516
rect 415176 3476 415182 3488
rect 428458 3476 428464 3488
rect 428516 3476 428522 3528
rect 429102 3476 429108 3528
rect 429160 3516 429166 3528
rect 445018 3516 445024 3528
rect 429160 3488 445024 3516
rect 429160 3476 429166 3488
rect 445018 3476 445024 3488
rect 445076 3476 445082 3528
rect 446858 3476 446864 3528
rect 446916 3516 446922 3528
rect 463970 3516 463976 3528
rect 446916 3488 463976 3516
rect 446916 3476 446922 3488
rect 463970 3476 463976 3488
rect 464028 3476 464034 3528
rect 464890 3476 464896 3528
rect 464948 3516 464954 3528
rect 485222 3516 485228 3528
rect 464948 3488 485228 3516
rect 464948 3476 464954 3488
rect 485222 3476 485228 3488
rect 485280 3476 485286 3528
rect 493962 3476 493968 3528
rect 494020 3516 494026 3528
rect 517146 3516 517152 3528
rect 494020 3488 517152 3516
rect 494020 3476 494026 3488
rect 517146 3476 517152 3488
rect 517204 3476 517210 3528
rect 520182 3476 520188 3528
rect 520240 3516 520246 3528
rect 546678 3516 546684 3528
rect 520240 3488 546684 3516
rect 520240 3476 520246 3488
rect 546678 3476 546684 3488
rect 546736 3476 546742 3528
rect 551922 3476 551928 3528
rect 551980 3516 551986 3528
rect 583386 3516 583392 3528
rect 551980 3488 583392 3516
rect 551980 3476 551986 3488
rect 583386 3476 583392 3488
rect 583444 3476 583450 3528
rect 57238 3408 57244 3460
rect 57296 3448 57302 3460
rect 57882 3448 57888 3460
rect 57296 3420 57888 3448
rect 57296 3408 57302 3420
rect 57882 3408 57888 3420
rect 57940 3408 57946 3460
rect 102226 3408 102232 3460
rect 102284 3448 102290 3460
rect 103422 3448 103428 3460
rect 102284 3420 103428 3448
rect 102284 3408 102290 3420
rect 103422 3408 103428 3420
rect 103480 3408 103486 3460
rect 106918 3408 106924 3460
rect 106976 3448 106982 3460
rect 107562 3448 107568 3460
rect 106976 3420 107568 3448
rect 106976 3408 106982 3420
rect 107562 3408 107568 3420
rect 107620 3408 107626 3460
rect 131758 3408 131764 3460
rect 131816 3448 131822 3460
rect 132402 3448 132408 3460
rect 131816 3420 132408 3448
rect 131816 3408 131822 3420
rect 132402 3408 132408 3420
rect 132460 3408 132466 3460
rect 189718 3408 189724 3460
rect 189776 3448 189782 3460
rect 190362 3448 190368 3460
rect 189776 3420 190368 3448
rect 189776 3408 189782 3420
rect 190362 3408 190368 3420
rect 190420 3408 190426 3460
rect 272426 3408 272432 3460
rect 272484 3448 272490 3460
rect 273898 3448 273904 3460
rect 272484 3420 273904 3448
rect 272484 3408 272490 3420
rect 273898 3408 273904 3420
rect 273956 3408 273962 3460
rect 279510 3408 279516 3460
rect 279568 3448 279574 3460
rect 281350 3448 281356 3460
rect 279568 3420 281356 3448
rect 279568 3408 279574 3420
rect 281350 3408 281356 3420
rect 281408 3408 281414 3460
rect 328362 3408 328368 3460
rect 328420 3448 328426 3460
rect 331582 3448 331588 3460
rect 328420 3420 331588 3448
rect 328420 3408 328426 3420
rect 331582 3408 331588 3420
rect 331640 3408 331646 3460
rect 338022 3408 338028 3460
rect 338080 3448 338086 3460
rect 342162 3448 342168 3460
rect 338080 3420 342168 3448
rect 338080 3408 338086 3420
rect 342162 3408 342168 3420
rect 342220 3408 342226 3460
rect 343542 3408 343548 3460
rect 343600 3448 343606 3460
rect 348050 3448 348056 3460
rect 343600 3420 348056 3448
rect 343600 3408 343606 3420
rect 348050 3408 348056 3420
rect 348108 3408 348114 3460
rect 348970 3408 348976 3460
rect 349028 3448 349034 3460
rect 354030 3448 354036 3460
rect 349028 3420 354036 3448
rect 349028 3408 349034 3420
rect 354030 3408 354036 3420
rect 354088 3408 354094 3460
rect 366910 3408 366916 3460
rect 366968 3448 366974 3460
rect 375282 3448 375288 3460
rect 366968 3420 375288 3448
rect 366968 3408 366974 3420
rect 375282 3408 375288 3420
rect 375340 3408 375346 3460
rect 379330 3408 379336 3460
rect 379388 3448 379394 3460
rect 389450 3448 389456 3460
rect 379388 3420 389456 3448
rect 379388 3408 379394 3420
rect 389450 3408 389456 3420
rect 389508 3408 389514 3460
rect 395982 3408 395988 3460
rect 396040 3448 396046 3460
rect 407206 3448 407212 3460
rect 396040 3420 407212 3448
rect 396040 3408 396046 3420
rect 407206 3408 407212 3420
rect 407264 3408 407270 3460
rect 411070 3408 411076 3460
rect 411128 3448 411134 3460
rect 424962 3448 424968 3460
rect 411128 3420 424968 3448
rect 411128 3408 411134 3420
rect 424962 3408 424968 3420
rect 425020 3408 425026 3460
rect 434622 3408 434628 3460
rect 434680 3448 434686 3460
rect 434680 3420 441614 3448
rect 434680 3408 434686 3420
rect 331030 3340 331036 3392
rect 331088 3380 331094 3392
rect 335078 3380 335084 3392
rect 331088 3352 335084 3380
rect 331088 3340 331094 3352
rect 335078 3340 335084 3352
rect 335136 3340 335142 3392
rect 390462 3340 390468 3392
rect 390520 3380 390526 3392
rect 401318 3380 401324 3392
rect 390520 3352 401324 3380
rect 390520 3340 390526 3352
rect 401318 3340 401324 3352
rect 401376 3340 401382 3392
rect 408310 3340 408316 3392
rect 408368 3380 408374 3392
rect 421374 3380 421380 3392
rect 408368 3352 421380 3380
rect 408368 3340 408374 3352
rect 421374 3340 421380 3352
rect 421432 3340 421438 3392
rect 424870 3340 424876 3392
rect 424928 3380 424934 3392
rect 440326 3380 440332 3392
rect 424928 3352 440332 3380
rect 424928 3340 424934 3352
rect 440326 3340 440332 3352
rect 440384 3340 440390 3392
rect 441586 3380 441614 3420
rect 447042 3408 447048 3460
rect 447100 3448 447106 3460
rect 465166 3448 465172 3460
rect 447100 3420 465172 3448
rect 447100 3408 447106 3420
rect 465166 3408 465172 3420
rect 465224 3408 465230 3460
rect 469122 3408 469128 3460
rect 469180 3448 469186 3460
rect 489914 3448 489920 3460
rect 469180 3420 489920 3448
rect 469180 3408 469186 3420
rect 489914 3408 489920 3420
rect 489972 3408 489978 3460
rect 498102 3408 498108 3460
rect 498160 3448 498166 3460
rect 521838 3448 521844 3460
rect 498160 3420 521844 3448
rect 498160 3408 498166 3420
rect 521838 3408 521844 3420
rect 521896 3408 521902 3460
rect 522850 3408 522856 3460
rect 522908 3448 522914 3460
rect 550266 3448 550272 3460
rect 522908 3420 550272 3448
rect 522908 3408 522914 3420
rect 550266 3408 550272 3420
rect 550324 3408 550330 3460
rect 550450 3408 550456 3460
rect 550508 3448 550514 3460
rect 580994 3448 581000 3460
rect 550508 3420 581000 3448
rect 550508 3408 550514 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 450906 3380 450912 3392
rect 441586 3352 450912 3380
rect 450906 3340 450912 3352
rect 450964 3340 450970 3392
rect 453942 3340 453948 3392
rect 454000 3380 454006 3392
rect 472250 3380 472256 3392
rect 454000 3352 472256 3380
rect 454000 3340 454006 3352
rect 472250 3340 472256 3352
rect 472308 3340 472314 3392
rect 474642 3340 474648 3392
rect 474700 3380 474706 3392
rect 495894 3380 495900 3392
rect 474700 3352 495900 3380
rect 474700 3340 474706 3352
rect 495894 3340 495900 3352
rect 495952 3340 495958 3392
rect 496722 3340 496728 3392
rect 496780 3380 496786 3392
rect 520734 3380 520740 3392
rect 496780 3352 520740 3380
rect 496780 3340 496786 3352
rect 520734 3340 520740 3352
rect 520792 3340 520798 3392
rect 535362 3340 535368 3392
rect 535420 3380 535426 3392
rect 563238 3380 563244 3392
rect 535420 3352 563244 3380
rect 535420 3340 535426 3352
rect 563238 3340 563244 3352
rect 563296 3340 563302 3392
rect 37240 3284 55214 3312
rect 37240 3272 37246 3284
rect 80882 3272 80888 3324
rect 80940 3312 80946 3324
rect 81342 3312 81348 3324
rect 80940 3284 81348 3312
rect 80940 3272 80946 3284
rect 81342 3272 81348 3284
rect 81400 3272 81406 3324
rect 85666 3272 85672 3324
rect 85724 3312 85730 3324
rect 86770 3312 86776 3324
rect 85724 3284 86776 3312
rect 85724 3272 85730 3284
rect 86770 3272 86776 3284
rect 86828 3272 86834 3324
rect 89162 3272 89168 3324
rect 89220 3312 89226 3324
rect 89622 3312 89628 3324
rect 89220 3284 89628 3312
rect 89220 3272 89226 3284
rect 89622 3272 89628 3284
rect 89680 3272 89686 3324
rect 93946 3272 93952 3324
rect 94004 3312 94010 3324
rect 95050 3312 95056 3324
rect 94004 3284 95056 3312
rect 94004 3272 94010 3284
rect 95050 3272 95056 3284
rect 95108 3272 95114 3324
rect 97442 3272 97448 3324
rect 97500 3312 97506 3324
rect 97902 3312 97908 3324
rect 97500 3284 97908 3312
rect 97500 3272 97506 3284
rect 97902 3272 97908 3284
rect 97960 3272 97966 3324
rect 196802 3272 196808 3324
rect 196860 3312 196866 3324
rect 197262 3312 197268 3324
rect 196860 3284 197268 3312
rect 196860 3272 196866 3284
rect 197262 3272 197268 3284
rect 197320 3272 197326 3324
rect 221550 3272 221556 3324
rect 221608 3312 221614 3324
rect 222102 3312 222108 3324
rect 221608 3284 222108 3312
rect 221608 3272 221614 3284
rect 222102 3272 222108 3284
rect 222160 3272 222166 3324
rect 262950 3272 262956 3324
rect 263008 3312 263014 3324
rect 263502 3312 263508 3324
rect 263008 3284 263508 3312
rect 263008 3272 263014 3284
rect 263502 3272 263508 3284
rect 263560 3272 263566 3324
rect 271230 3272 271236 3324
rect 271288 3312 271294 3324
rect 271782 3312 271788 3324
rect 271288 3284 271788 3312
rect 271288 3272 271294 3284
rect 271782 3272 271788 3284
rect 271840 3272 271846 3324
rect 287790 3272 287796 3324
rect 287848 3312 287854 3324
rect 288342 3312 288348 3324
rect 287848 3284 288348 3312
rect 287848 3272 287854 3284
rect 288342 3272 288348 3284
rect 288400 3272 288406 3324
rect 317322 3272 317328 3324
rect 317380 3312 317386 3324
rect 318518 3312 318524 3324
rect 317380 3284 318524 3312
rect 317380 3272 317386 3284
rect 318518 3272 318524 3284
rect 318576 3272 318582 3324
rect 339310 3272 339316 3324
rect 339368 3312 339374 3324
rect 343358 3312 343364 3324
rect 339368 3284 343364 3312
rect 339368 3272 339374 3284
rect 343358 3272 343364 3284
rect 343416 3272 343422 3324
rect 347682 3272 347688 3324
rect 347740 3312 347746 3324
rect 352834 3312 352840 3324
rect 347740 3284 352840 3312
rect 347740 3272 347746 3284
rect 352834 3272 352840 3284
rect 352892 3272 352898 3324
rect 355962 3272 355968 3324
rect 356020 3312 356026 3324
rect 362310 3312 362316 3324
rect 356020 3284 362316 3312
rect 356020 3272 356026 3284
rect 362310 3272 362316 3284
rect 362368 3272 362374 3324
rect 391750 3272 391756 3324
rect 391808 3312 391814 3324
rect 402514 3312 402520 3324
rect 391808 3284 402520 3312
rect 391808 3272 391814 3284
rect 402514 3272 402520 3284
rect 402572 3272 402578 3324
rect 406930 3272 406936 3324
rect 406988 3312 406994 3324
rect 418982 3312 418988 3324
rect 406988 3284 418988 3312
rect 406988 3272 406994 3284
rect 418982 3272 418988 3284
rect 419040 3272 419046 3324
rect 426342 3272 426348 3324
rect 426400 3312 426406 3324
rect 441522 3312 441528 3324
rect 426400 3284 441528 3312
rect 426400 3272 426406 3284
rect 441522 3272 441528 3284
rect 441580 3272 441586 3324
rect 445662 3272 445668 3324
rect 445720 3312 445726 3324
rect 462774 3312 462780 3324
rect 445720 3284 462780 3312
rect 445720 3272 445726 3284
rect 462774 3272 462780 3284
rect 462832 3272 462838 3324
rect 473262 3272 473268 3324
rect 473320 3312 473326 3324
rect 493502 3312 493508 3324
rect 473320 3284 493508 3312
rect 473320 3272 473326 3284
rect 493502 3272 493508 3284
rect 493560 3272 493566 3324
rect 500862 3272 500868 3324
rect 500920 3312 500926 3324
rect 525426 3312 525432 3324
rect 500920 3284 525432 3312
rect 500920 3272 500926 3284
rect 525426 3272 525432 3284
rect 525484 3272 525490 3324
rect 528462 3272 528468 3324
rect 528520 3312 528526 3324
rect 556154 3312 556160 3324
rect 528520 3284 556160 3312
rect 528520 3272 528526 3284
rect 556154 3272 556160 3284
rect 556212 3272 556218 3324
rect 101030 3204 101036 3256
rect 101088 3244 101094 3256
rect 102042 3244 102048 3256
rect 101088 3216 102048 3244
rect 101088 3204 101094 3216
rect 102042 3204 102048 3216
rect 102100 3204 102106 3256
rect 183738 3204 183744 3256
rect 183796 3244 183802 3256
rect 184842 3244 184848 3256
rect 183796 3216 184848 3244
rect 183796 3204 183802 3216
rect 184842 3204 184848 3216
rect 184900 3204 184906 3256
rect 200298 3204 200304 3256
rect 200356 3244 200362 3256
rect 201402 3244 201408 3256
rect 200356 3216 201408 3244
rect 200356 3204 200362 3216
rect 201402 3204 201408 3216
rect 201460 3204 201466 3256
rect 225138 3204 225144 3256
rect 225196 3244 225202 3256
rect 226242 3244 226248 3256
rect 225196 3216 226248 3244
rect 225196 3204 225202 3216
rect 226242 3204 226248 3216
rect 226300 3204 226306 3256
rect 258258 3204 258264 3256
rect 258316 3244 258322 3256
rect 259362 3244 259368 3256
rect 258316 3216 259368 3244
rect 258316 3204 258322 3216
rect 259362 3204 259368 3216
rect 259420 3204 259426 3256
rect 336642 3204 336648 3256
rect 336700 3244 336706 3256
rect 340966 3244 340972 3256
rect 336700 3216 340972 3244
rect 336700 3204 336706 3216
rect 340966 3204 340972 3216
rect 341024 3204 341030 3256
rect 346302 3204 346308 3256
rect 346360 3244 346366 3256
rect 351638 3244 351644 3256
rect 346360 3216 351644 3244
rect 346360 3204 346366 3216
rect 351638 3204 351644 3216
rect 351696 3204 351702 3256
rect 405642 3204 405648 3256
rect 405700 3244 405706 3256
rect 417878 3244 417884 3256
rect 405700 3216 417884 3244
rect 405700 3204 405706 3216
rect 417878 3204 417884 3216
rect 417936 3204 417942 3256
rect 420822 3204 420828 3256
rect 420880 3244 420886 3256
rect 434438 3244 434444 3256
rect 420880 3216 434444 3244
rect 420880 3204 420886 3216
rect 434438 3204 434444 3216
rect 434496 3204 434502 3256
rect 441430 3204 441436 3256
rect 441488 3244 441494 3256
rect 458082 3244 458088 3256
rect 441488 3216 458088 3244
rect 441488 3204 441494 3216
rect 458082 3204 458088 3216
rect 458140 3204 458146 3256
rect 464982 3204 464988 3256
rect 465040 3244 465046 3256
rect 484026 3244 484032 3256
rect 465040 3216 484032 3244
rect 465040 3204 465046 3216
rect 484026 3204 484032 3216
rect 484084 3204 484090 3256
rect 485682 3204 485688 3256
rect 485740 3244 485746 3256
rect 507670 3244 507676 3256
rect 485740 3216 507676 3244
rect 485740 3204 485746 3216
rect 507670 3204 507676 3216
rect 507728 3204 507734 3256
rect 507762 3204 507768 3256
rect 507820 3244 507826 3256
rect 532510 3244 532516 3256
rect 507820 3216 532516 3244
rect 507820 3204 507826 3216
rect 532510 3204 532516 3216
rect 532568 3204 532574 3256
rect 539502 3204 539508 3256
rect 539560 3244 539566 3256
rect 568022 3244 568028 3256
rect 539560 3216 568028 3244
rect 539560 3204 539566 3216
rect 568022 3204 568028 3216
rect 568080 3204 568086 3256
rect 241698 3136 241704 3188
rect 241756 3176 241762 3188
rect 242802 3176 242808 3188
rect 241756 3148 242808 3176
rect 241756 3136 241762 3148
rect 242802 3136 242808 3148
rect 242860 3136 242866 3188
rect 321370 3136 321376 3188
rect 321428 3176 321434 3188
rect 324406 3176 324412 3188
rect 321428 3148 324412 3176
rect 321428 3136 321434 3148
rect 324406 3136 324412 3148
rect 324464 3136 324470 3188
rect 329742 3136 329748 3188
rect 329800 3176 329806 3188
rect 332686 3176 332692 3188
rect 329800 3148 332692 3176
rect 329800 3136 329806 3148
rect 332686 3136 332692 3148
rect 332744 3136 332750 3188
rect 419442 3136 419448 3188
rect 419500 3176 419506 3188
rect 433242 3176 433248 3188
rect 419500 3148 433248 3176
rect 419500 3136 419506 3148
rect 433242 3136 433248 3148
rect 433300 3136 433306 3188
rect 438762 3136 438768 3188
rect 438820 3176 438826 3188
rect 454494 3176 454500 3188
rect 438820 3148 454500 3176
rect 438820 3136 438826 3148
rect 454494 3136 454500 3148
rect 454552 3136 454558 3188
rect 457990 3136 457996 3188
rect 458048 3176 458054 3188
rect 476942 3176 476948 3188
rect 458048 3148 476948 3176
rect 458048 3136 458054 3148
rect 476942 3136 476948 3148
rect 477000 3136 477006 3188
rect 482922 3136 482928 3188
rect 482980 3176 482986 3188
rect 504174 3176 504180 3188
rect 482980 3148 504180 3176
rect 482980 3136 482986 3148
rect 504174 3136 504180 3148
rect 504232 3136 504238 3188
rect 504818 3136 504824 3188
rect 504876 3176 504882 3188
rect 529014 3176 529020 3188
rect 504876 3148 529020 3176
rect 504876 3136 504882 3148
rect 529014 3136 529020 3148
rect 529072 3136 529078 3188
rect 536742 3136 536748 3188
rect 536800 3176 536806 3188
rect 564434 3176 564440 3188
rect 536800 3148 564440 3176
rect 536800 3136 536806 3148
rect 564434 3136 564440 3148
rect 564492 3136 564498 3188
rect 118786 3068 118792 3120
rect 118844 3108 118850 3120
rect 119798 3108 119804 3120
rect 118844 3080 119804 3108
rect 118844 3068 118850 3080
rect 119798 3068 119804 3080
rect 119856 3068 119862 3120
rect 246390 3068 246396 3120
rect 246448 3108 246454 3120
rect 246942 3108 246948 3120
rect 246448 3080 246948 3108
rect 246448 3068 246454 3080
rect 246942 3068 246948 3080
rect 247000 3068 247006 3120
rect 360102 3068 360108 3120
rect 360160 3108 360166 3120
rect 367002 3108 367008 3120
rect 360160 3080 367008 3108
rect 360160 3068 360166 3080
rect 367002 3068 367008 3080
rect 367060 3068 367066 3120
rect 368382 3068 368388 3120
rect 368440 3108 368446 3120
rect 376478 3108 376484 3120
rect 368440 3080 376484 3108
rect 368440 3068 368446 3080
rect 376478 3068 376484 3080
rect 376536 3068 376542 3120
rect 427722 3068 427728 3120
rect 427780 3108 427786 3120
rect 442626 3108 442632 3120
rect 427780 3080 442632 3108
rect 427780 3068 427786 3080
rect 442626 3068 442632 3080
rect 442684 3068 442690 3120
rect 442902 3068 442908 3120
rect 442960 3108 442966 3120
rect 459186 3108 459192 3120
rect 442960 3080 459192 3108
rect 442960 3068 442966 3080
rect 459186 3068 459192 3080
rect 459244 3068 459250 3120
rect 459462 3068 459468 3120
rect 459520 3108 459526 3120
rect 478138 3108 478144 3120
rect 459520 3080 478144 3108
rect 459520 3068 459526 3080
rect 478138 3068 478144 3080
rect 478196 3068 478202 3120
rect 478782 3068 478788 3120
rect 478840 3108 478846 3120
rect 499390 3108 499396 3120
rect 478840 3080 499396 3108
rect 478840 3068 478846 3080
rect 499390 3068 499396 3080
rect 499448 3068 499454 3120
rect 500678 3068 500684 3120
rect 500736 3108 500742 3120
rect 524230 3108 524236 3120
rect 500736 3080 524236 3108
rect 500736 3068 500742 3080
rect 524230 3068 524236 3080
rect 524288 3068 524294 3120
rect 532602 3068 532608 3120
rect 532660 3108 532666 3120
rect 559742 3108 559748 3120
rect 532660 3080 559748 3108
rect 532660 3068 532666 3080
rect 559742 3068 559748 3080
rect 559800 3068 559806 3120
rect 150618 3000 150624 3052
rect 150676 3040 150682 3052
rect 151722 3040 151728 3052
rect 150676 3012 151728 3040
rect 150676 3000 150682 3012
rect 151722 3000 151728 3012
rect 151780 3000 151786 3052
rect 168374 3000 168380 3052
rect 168432 3040 168438 3052
rect 169478 3040 169484 3052
rect 168432 3012 169484 3040
rect 168432 3000 168438 3012
rect 169478 3000 169484 3012
rect 169536 3000 169542 3052
rect 208578 3000 208584 3052
rect 208636 3040 208642 3052
rect 209682 3040 209688 3052
rect 208636 3012 209688 3040
rect 208636 3000 208642 3012
rect 209682 3000 209688 3012
rect 209740 3000 209746 3052
rect 226334 3000 226340 3052
rect 226392 3040 226398 3052
rect 227438 3040 227444 3052
rect 226392 3012 227444 3040
rect 226392 3000 226398 3012
rect 227438 3000 227444 3012
rect 227496 3000 227502 3052
rect 248782 3000 248788 3052
rect 248840 3040 248846 3052
rect 249702 3040 249708 3052
rect 248840 3012 249708 3040
rect 248840 3000 248846 3012
rect 249702 3000 249708 3012
rect 249760 3000 249766 3052
rect 259454 3000 259460 3052
rect 259512 3040 259518 3052
rect 260558 3040 260564 3052
rect 259512 3012 260564 3040
rect 259512 3000 259518 3012
rect 260558 3000 260564 3012
rect 260616 3000 260622 3052
rect 274818 3000 274824 3052
rect 274876 3040 274882 3052
rect 277026 3040 277032 3052
rect 274876 3012 277032 3040
rect 274876 3000 274882 3012
rect 277026 3000 277032 3012
rect 277084 3000 277090 3052
rect 284294 3000 284300 3052
rect 284352 3040 284358 3052
rect 285582 3040 285588 3052
rect 284352 3012 285588 3040
rect 284352 3000 284358 3012
rect 285582 3000 285588 3012
rect 285640 3000 285646 3052
rect 302418 3000 302424 3052
rect 302476 3040 302482 3052
rect 303154 3040 303160 3052
rect 302476 3012 303160 3040
rect 302476 3000 302482 3012
rect 303154 3000 303160 3012
rect 303212 3000 303218 3052
rect 317230 3000 317236 3052
rect 317288 3040 317294 3052
rect 319714 3040 319720 3052
rect 317288 3012 319720 3040
rect 317288 3000 317294 3012
rect 319714 3000 319720 3012
rect 319772 3000 319778 3052
rect 322842 3000 322848 3052
rect 322900 3040 322906 3052
rect 325602 3040 325608 3052
rect 322900 3012 325608 3040
rect 322900 3000 322906 3012
rect 325602 3000 325608 3012
rect 325660 3000 325666 3052
rect 431862 3000 431868 3052
rect 431920 3040 431926 3052
rect 447410 3040 447416 3052
rect 431920 3012 447416 3040
rect 431920 3000 431926 3012
rect 447410 3000 447416 3012
rect 447468 3000 447474 3052
rect 448422 3000 448428 3052
rect 448480 3040 448486 3052
rect 466270 3040 466276 3052
rect 448480 3012 466276 3040
rect 448480 3000 448486 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 471882 3000 471888 3052
rect 471940 3040 471946 3052
rect 492306 3040 492312 3052
rect 471940 3012 492312 3040
rect 471940 3000 471946 3012
rect 492306 3000 492312 3012
rect 492364 3000 492370 3052
rect 525702 3000 525708 3052
rect 525760 3040 525766 3052
rect 552658 3040 552664 3052
rect 525760 3012 552664 3040
rect 525760 3000 525766 3012
rect 552658 3000 552664 3012
rect 552716 3000 552722 3052
rect 73798 2932 73804 2984
rect 73856 2972 73862 2984
rect 74442 2972 74448 2984
rect 73856 2944 74448 2972
rect 73856 2932 73862 2944
rect 74442 2932 74448 2944
rect 74500 2932 74506 2984
rect 313182 2932 313188 2984
rect 313240 2972 313246 2984
rect 315022 2972 315028 2984
rect 313240 2944 315028 2972
rect 313240 2932 313246 2944
rect 315022 2932 315028 2944
rect 315080 2932 315086 2984
rect 463602 2932 463608 2984
rect 463660 2972 463666 2984
rect 482830 2972 482836 2984
rect 463660 2944 482836 2972
rect 463660 2932 463666 2944
rect 482830 2932 482836 2944
rect 482888 2932 482894 2984
rect 526898 2932 526904 2984
rect 526956 2972 526962 2984
rect 553762 2972 553768 2984
rect 526956 2944 553768 2972
rect 526956 2932 526962 2944
rect 553762 2932 553768 2944
rect 553820 2932 553826 2984
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 8110 2904 8116 2916
rect 624 2876 8116 2904
rect 624 2864 630 2876
rect 8110 2864 8116 2876
rect 8168 2864 8174 2916
rect 135254 2864 135260 2916
rect 135312 2904 135318 2916
rect 136542 2904 136548 2916
rect 135312 2876 136548 2904
rect 135312 2864 135318 2876
rect 136542 2864 136548 2876
rect 136600 2864 136606 2916
rect 349062 2864 349068 2916
rect 349120 2904 349126 2916
rect 355226 2904 355232 2916
rect 349120 2876 355232 2904
rect 349120 2864 349126 2876
rect 355226 2864 355232 2876
rect 355284 2864 355290 2916
rect 365622 2864 365628 2916
rect 365680 2904 365686 2916
rect 372890 2904 372896 2916
rect 365680 2876 372896 2904
rect 365680 2864 365686 2876
rect 372890 2864 372896 2876
rect 372948 2864 372954 2916
rect 456702 2864 456708 2916
rect 456760 2904 456766 2916
rect 474550 2904 474556 2916
rect 456760 2876 474556 2904
rect 456760 2864 456766 2876
rect 474550 2864 474556 2876
rect 474608 2864 474614 2916
rect 529842 2864 529848 2916
rect 529900 2904 529906 2916
rect 557350 2904 557356 2916
rect 529900 2876 557356 2904
rect 529900 2864 529906 2876
rect 557350 2864 557356 2876
rect 557408 2864 557414 2916
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 8018 2836 8024 2848
rect 1728 2808 8024 2836
rect 1728 2796 1734 2808
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 449710 2796 449716 2848
rect 449768 2836 449774 2848
rect 467466 2836 467472 2848
rect 449768 2808 467472 2836
rect 449768 2796 449774 2808
rect 467466 2796 467472 2808
rect 467524 2796 467530 2848
rect 522942 2796 522948 2848
rect 523000 2836 523006 2848
rect 549070 2836 549076 2848
rect 523000 2808 549076 2836
rect 523000 2796 523006 2808
rect 549070 2796 549076 2808
rect 549128 2796 549134 2848
<< via1 >>
rect 154120 700952 154172 701004
rect 329840 700952 329892 701004
rect 137836 700884 137888 700936
rect 325700 700884 325752 700936
rect 257988 700816 258040 700868
rect 462320 700816 462372 700868
rect 263508 700748 263560 700800
rect 478512 700748 478564 700800
rect 89168 700680 89220 700732
rect 343640 700680 343692 700732
rect 72976 700612 73028 700664
rect 339500 700612 339552 700664
rect 244188 700544 244240 700596
rect 527180 700544 527232 700596
rect 249708 700476 249760 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 347872 700408 347924 700460
rect 349804 700408 349856 700460
rect 364984 700408 365036 700460
rect 24308 700340 24360 700392
rect 357440 700340 357492 700392
rect 8116 700272 8168 700324
rect 353300 700272 353352 700324
rect 356704 700272 356756 700324
rect 494796 700272 494848 700324
rect 275928 700204 275980 700256
rect 413652 700204 413704 700256
rect 271788 700136 271840 700188
rect 397460 700136 397512 700188
rect 202788 700068 202840 700120
rect 311900 700068 311952 700120
rect 218980 700000 219032 700052
rect 316040 700000 316092 700052
rect 289728 699932 289780 699984
rect 348792 699932 348844 699984
rect 285588 699864 285640 699916
rect 332508 699864 332560 699916
rect 235172 699796 235224 699848
rect 238024 699796 238076 699848
rect 267648 699796 267700 699848
rect 298100 699796 298152 699848
rect 283840 699728 283892 699780
rect 302240 699728 302292 699780
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 555424 699660 555476 699712
rect 559656 699660 559708 699712
rect 230388 696940 230440 696992
rect 580172 696940 580224 696992
rect 235908 683204 235960 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 361580 683136 361632 683188
rect 294236 675996 294288 676048
rect 299480 675996 299532 676048
rect 280528 675928 280580 675980
rect 349804 675928 349856 675980
rect 238024 675860 238076 675912
rect 307852 675860 307904 675912
rect 253112 675792 253164 675844
rect 356704 675792 356756 675844
rect 171048 675724 171100 675776
rect 321560 675724 321612 675776
rect 266820 675656 266872 675708
rect 429200 675656 429252 675708
rect 106188 675588 106240 675640
rect 335268 675588 335320 675640
rect 239496 675520 239548 675572
rect 555424 675520 555476 675572
rect 175556 675452 175608 675504
rect 554136 675452 554188 675504
rect 157340 675384 157392 675436
rect 558276 675384 558328 675436
rect 143632 675316 143684 675368
rect 576216 675316 576268 675368
rect 130016 675248 130068 675300
rect 574836 675248 574888 675300
rect 25596 675180 25648 675232
rect 499488 675180 499540 675232
rect 29736 675112 29788 675164
rect 513104 675112 513156 675164
rect 75276 675044 75328 675096
rect 565084 675044 565136 675096
rect 43352 674976 43404 675028
rect 552664 674976 552716 675028
rect 7564 674908 7616 674960
rect 526812 674908 526864 674960
rect 52460 674840 52512 674892
rect 576124 674840 576176 674892
rect 218060 674772 218112 674824
rect 412824 674772 412876 674824
rect 152832 674704 152884 674756
rect 382280 674704 382332 674756
rect 125416 674636 125468 674688
rect 368664 674636 368716 674688
rect 200120 674568 200172 674620
rect 481180 674568 481232 674620
rect 14556 674500 14608 674552
rect 408224 674500 408276 674552
rect 180156 674432 180208 674484
rect 572076 674432 572128 674484
rect 166448 674364 166500 674416
rect 571984 674364 572036 674416
rect 111708 674296 111760 674348
rect 155776 674296 155828 674348
rect 161940 674296 161992 674348
rect 570604 674296 570656 674348
rect 26884 674228 26936 674280
rect 440148 674228 440200 674280
rect 17316 674160 17368 674212
rect 435548 674160 435600 674212
rect 148232 674092 148284 674144
rect 565176 674092 565228 674144
rect 18696 674024 18748 674076
rect 449256 674024 449308 674076
rect 11796 673956 11848 674008
rect 453856 673956 453908 674008
rect 120908 673888 120960 673940
rect 561036 673888 561088 673940
rect 31024 673820 31076 673872
rect 476672 673820 476724 673872
rect 107200 673752 107252 673804
rect 555516 673752 555568 673804
rect 17224 673684 17276 673736
rect 494888 673684 494940 673736
rect 22744 673616 22796 673668
rect 503996 673616 504048 673668
rect 25504 673548 25556 673600
rect 517704 673548 517756 673600
rect 4896 673480 4948 673532
rect 522212 673480 522264 673532
rect 212080 673344 212132 673396
rect 558368 673344 558420 673396
rect 3516 673276 3568 673328
rect 200120 673276 200172 673328
rect 225788 673276 225840 673328
rect 579528 673276 579580 673328
rect 198372 673208 198424 673260
rect 556988 673208 557040 673260
rect 7748 673140 7800 673192
rect 376300 673140 376352 673192
rect 184756 673072 184808 673124
rect 554228 673072 554280 673124
rect 11888 673004 11940 673056
rect 390008 673004 390060 673056
rect 171048 672936 171100 672988
rect 552756 672936 552808 672988
rect 14648 672868 14700 672920
rect 403624 672868 403676 672920
rect 16028 672800 16080 672852
rect 417332 672800 417384 672852
rect 155776 672732 155828 672784
rect 580264 672732 580316 672784
rect 17408 672664 17460 672716
rect 431040 672664 431092 672716
rect 139124 672596 139176 672648
rect 556896 672596 556948 672648
rect 18788 672528 18840 672580
rect 444748 672528 444800 672580
rect 21456 672460 21508 672512
rect 458364 672460 458416 672512
rect 31116 672392 31168 672444
rect 472072 672392 472124 672444
rect 22836 672324 22888 672376
rect 485780 672324 485832 672376
rect 98092 672256 98144 672308
rect 578884 672256 578936 672308
rect 84384 672188 84436 672240
rect 569224 672188 569276 672240
rect 61568 672120 61620 672172
rect 562324 672120 562376 672172
rect 3424 672052 3476 672104
rect 508596 672052 508648 672104
rect 3608 671984 3660 672036
rect 218060 671984 218112 672036
rect 221464 671984 221516 672036
rect 557080 671984 557132 672036
rect 27068 671916 27120 671968
rect 367284 671916 367336 671968
rect 368664 671916 368716 671968
rect 580356 671916 580408 671968
rect 28356 671848 28408 671900
rect 380992 671848 381044 671900
rect 217048 671780 217100 671832
rect 569500 671780 569552 671832
rect 26976 671712 27028 671764
rect 385132 671712 385184 671764
rect 421564 671755 421616 671764
rect 421564 671721 421573 671755
rect 421573 671721 421607 671755
rect 421607 671721 421616 671755
rect 421564 671712 421616 671721
rect 207848 671644 207900 671696
rect 569408 671644 569460 671696
rect 203248 671576 203300 671628
rect 566648 671576 566700 671628
rect 3332 671508 3384 671560
rect 371332 671508 371384 671560
rect 382280 671508 382332 671560
rect 580448 671508 580500 671560
rect 66260 671483 66312 671492
rect 66260 671449 66269 671483
rect 66269 671449 66303 671483
rect 66303 671449 66312 671483
rect 66260 671440 66312 671449
rect 70952 671483 71004 671492
rect 70952 671449 70961 671483
rect 70961 671449 70995 671483
rect 70995 671449 71004 671483
rect 70952 671440 71004 671449
rect 79968 671483 80020 671492
rect 79968 671449 79977 671483
rect 79977 671449 80011 671483
rect 80011 671449 80020 671483
rect 79968 671440 80020 671449
rect 93676 671483 93728 671492
rect 93676 671449 93685 671483
rect 93685 671449 93719 671483
rect 93719 671449 93728 671483
rect 93676 671440 93728 671449
rect 134800 671483 134852 671492
rect 134800 671449 134809 671483
rect 134809 671449 134843 671483
rect 134843 671449 134852 671483
rect 134800 671440 134852 671449
rect 194232 671440 194284 671492
rect 578976 671440 579028 671492
rect 7656 671372 7708 671424
rect 398840 671372 398892 671424
rect 28264 671304 28316 671356
rect 426256 671372 426308 671424
rect 15936 671236 15988 671288
rect 462596 671372 462648 671424
rect 467196 671415 467248 671424
rect 467196 671381 467205 671415
rect 467205 671381 467239 671415
rect 467239 671381 467248 671415
rect 467196 671372 467248 671381
rect 490104 671415 490156 671424
rect 490104 671381 490113 671415
rect 490113 671381 490147 671415
rect 490147 671381 490156 671415
rect 490104 671372 490156 671381
rect 21364 671100 21416 671152
rect 562416 671168 562468 671220
rect 10324 671032 10376 671084
rect 14464 670964 14516 671016
rect 573364 670896 573416 670948
rect 558184 670828 558236 670880
rect 574744 670760 574796 670812
rect 566464 670692 566516 670744
rect 3332 658180 3384 658232
rect 27068 658180 27120 658232
rect 569500 644376 569552 644428
rect 580172 644376 580224 644428
rect 3332 633360 3384 633412
rect 7748 633360 7800 633412
rect 557080 632000 557132 632052
rect 579712 632000 579764 632052
rect 3332 619556 3384 619608
rect 26976 619556 27028 619608
rect 558368 618196 558420 618248
rect 579804 618196 579856 618248
rect 3056 607112 3108 607164
rect 28356 607112 28408 607164
rect 566648 591948 566700 592000
rect 580172 591948 580224 592000
rect 3332 580932 3384 580984
rect 11888 580932 11940 580984
rect 569408 578144 569460 578196
rect 580172 578144 580224 578196
rect 3148 567060 3200 567112
rect 7656 567060 7708 567112
rect 556988 564340 557040 564392
rect 580172 564340 580224 564392
rect 2964 554684 3016 554736
rect 10416 554684 10468 554736
rect 552848 538160 552900 538212
rect 580172 538160 580224 538212
rect 3148 528504 3200 528556
rect 14648 528504 14700 528556
rect 554228 511912 554280 511964
rect 580172 511912 580224 511964
rect 2964 502256 3016 502308
rect 14556 502256 14608 502308
rect 554136 485732 554188 485784
rect 580172 485732 580224 485784
rect 3240 476008 3292 476060
rect 16028 476008 16080 476060
rect 572076 471928 572128 471980
rect 580172 471928 580224 471980
rect 3056 463632 3108 463684
rect 28264 463632 28316 463684
rect 552756 458124 552808 458176
rect 580172 458124 580224 458176
rect 3332 449828 3384 449880
rect 15936 449828 15988 449880
rect 570604 431876 570656 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 17408 423580 17460 423632
rect 571984 419432 572036 419484
rect 579712 419432 579764 419484
rect 2964 411204 3016 411256
rect 26884 411204 26936 411256
rect 558276 405628 558328 405680
rect 579804 405628 579856 405680
rect 3332 398760 3384 398812
rect 17316 398760 17368 398812
rect 565176 379448 565228 379500
rect 579804 379448 579856 379500
rect 3332 372512 3384 372564
rect 18788 372512 18840 372564
rect 3332 358708 3384 358760
rect 11796 358708 11848 358760
rect 576216 353200 576268 353252
rect 580172 353200 580224 353252
rect 3332 346332 3384 346384
rect 18696 346332 18748 346384
rect 562416 325592 562468 325644
rect 580172 325592 580224 325644
rect 3332 320084 3384 320136
rect 21456 320084 21508 320136
rect 556896 313216 556948 313268
rect 580172 313216 580224 313268
rect 3332 306280 3384 306332
rect 10324 306280 10376 306332
rect 574836 299412 574888 299464
rect 580172 299412 580224 299464
rect 3332 293904 3384 293956
rect 21364 293904 21416 293956
rect 561036 273164 561088 273216
rect 580172 273164 580224 273216
rect 2964 267656 3016 267708
rect 31116 267656 31168 267708
rect 573456 245556 573508 245608
rect 580172 245556 580224 245608
rect 3516 241408 3568 241460
rect 31024 241408 31076 241460
rect 555516 233180 555568 233232
rect 580172 233180 580224 233232
rect 3332 215228 3384 215280
rect 22836 215228 22888 215280
rect 569316 206932 569368 206984
rect 579804 206932 579856 206984
rect 3056 202784 3108 202836
rect 17224 202784 17276 202836
rect 573364 193128 573416 193180
rect 580172 193128 580224 193180
rect 3516 188980 3568 189032
rect 14464 188980 14516 189032
rect 566556 166948 566608 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 25596 164160 25648 164212
rect 574744 153144 574796 153196
rect 580172 153144 580224 153196
rect 3516 150424 3568 150476
rect 4896 150424 4948 150476
rect 569224 139340 569276 139392
rect 580172 139340 580224 139392
rect 3424 137912 3476 137964
rect 22744 137912 22796 137964
rect 565084 126896 565136 126948
rect 580172 126896 580224 126948
rect 558184 113092 558236 113144
rect 579804 113092 579856 113144
rect 3148 111732 3200 111784
rect 29736 111732 29788 111784
rect 566464 100648 566516 100700
rect 580172 100648 580224 100700
rect 562324 86912 562376 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 25504 85484 25556 85536
rect 576124 73108 576176 73160
rect 580172 73108 580224 73160
rect 3424 71612 3476 71664
rect 7564 71612 7616 71664
rect 554044 60664 554096 60716
rect 580172 60664 580224 60716
rect 2780 58624 2832 58676
rect 4804 58624 4856 58676
rect 560944 46860 560996 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 29644 45500 29696 45552
rect 3148 33056 3200 33108
rect 11704 33056 11756 33108
rect 556804 33056 556856 33108
rect 580172 33056 580224 33108
rect 20628 30268 20680 30320
rect 50344 30268 50396 30320
rect 50988 30268 51040 30320
rect 76748 30268 76800 30320
rect 78588 30268 78640 30320
rect 101036 30268 101088 30320
rect 101956 30268 102008 30320
rect 122104 30268 122156 30320
rect 128268 30268 128320 30320
rect 145288 30268 145340 30320
rect 146208 30268 146260 30320
rect 162216 30268 162268 30320
rect 168288 30268 168340 30320
rect 181168 30268 181220 30320
rect 183468 30268 183520 30320
rect 194876 30268 194928 30320
rect 200028 30268 200080 30320
rect 209688 30268 209740 30320
rect 224868 30268 224920 30320
rect 231768 30268 231820 30320
rect 244096 30268 244148 30320
rect 248696 30268 248748 30320
rect 255228 30268 255280 30320
rect 259184 30268 259236 30320
rect 277308 30268 277360 30320
rect 278228 30268 278280 30320
rect 286968 30268 287020 30320
rect 287704 30268 287756 30320
rect 315120 30268 315172 30320
rect 316224 30268 316276 30320
rect 16488 30200 16540 30252
rect 40960 30200 41012 30252
rect 48228 30200 48280 30252
rect 54576 30200 54628 30252
rect 56508 30200 56560 30252
rect 81992 30200 82044 30252
rect 86868 30200 86920 30252
rect 109408 30200 109460 30252
rect 111616 30200 111668 30252
rect 130568 30200 130620 30252
rect 155776 30200 155828 30252
rect 170588 30200 170640 30252
rect 179328 30200 179380 30252
rect 191748 30200 191800 30252
rect 193128 30200 193180 30252
rect 203340 30200 203392 30252
rect 205548 30200 205600 30252
rect 214932 30200 214984 30252
rect 223488 30200 223540 30252
rect 230756 30200 230808 30252
rect 253848 30200 253900 30252
rect 258172 30200 258224 30252
rect 470140 30200 470192 30252
rect 471336 30200 471388 30252
rect 23388 30132 23440 30184
rect 52460 30132 52512 30184
rect 53656 30132 53708 30184
rect 78864 30132 78916 30184
rect 88248 30132 88300 30184
rect 110512 30132 110564 30184
rect 113088 30132 113140 30184
rect 132684 30132 132736 30184
rect 133788 30132 133840 30184
rect 150624 30132 150676 30184
rect 158628 30132 158680 30184
rect 172704 30132 172756 30184
rect 175188 30132 175240 30184
rect 187516 30132 187568 30184
rect 190368 30132 190420 30184
rect 201224 30132 201276 30184
rect 202788 30132 202840 30184
rect 211712 30132 211764 30184
rect 216588 30132 216640 30184
rect 224408 30132 224460 30184
rect 244188 30132 244240 30184
rect 249708 30132 249760 30184
rect 10968 30064 11020 30116
rect 40776 30064 40828 30116
rect 36636 29996 36688 30048
rect 38568 29996 38620 30048
rect 66168 30064 66220 30116
rect 67548 30064 67600 30116
rect 91560 30064 91612 30116
rect 92388 30064 92440 30116
rect 113640 30064 113692 30116
rect 124128 30064 124180 30116
rect 142160 30064 142212 30116
rect 147588 30064 147640 30116
rect 163228 30064 163280 30116
rect 166908 30064 166960 30116
rect 180156 30064 180208 30116
rect 182088 30064 182140 30116
rect 193864 30064 193916 30116
rect 195888 30064 195940 30116
rect 206468 30064 206520 30116
rect 206928 30064 206980 30116
rect 215944 30064 215996 30116
rect 217968 30064 218020 30116
rect 225512 30064 225564 30116
rect 226248 30064 226300 30116
rect 232872 30064 232924 30116
rect 233148 30064 233200 30116
rect 239220 30064 239272 30116
rect 63040 29996 63092 30048
rect 63408 29996 63460 30048
rect 88340 29996 88392 30048
rect 89628 29996 89680 30048
rect 111524 29996 111576 30048
rect 111708 29996 111760 30048
rect 131580 29996 131632 30048
rect 132408 29996 132460 30048
rect 149520 29996 149572 30048
rect 154488 29996 154540 30048
rect 169576 29996 169628 30048
rect 173716 29996 173768 30048
rect 186412 29996 186464 30048
rect 197268 29996 197320 30048
rect 207572 29996 207624 30048
rect 13728 29928 13780 29980
rect 15108 29860 15160 29912
rect 40960 29928 41012 29980
rect 46204 29928 46256 29980
rect 71504 29928 71556 29980
rect 82728 29928 82780 29980
rect 105268 29928 105320 29980
rect 108948 29928 109000 29980
rect 128452 29928 128504 29980
rect 131028 29928 131080 29980
rect 148508 29928 148560 29980
rect 148968 29928 149020 29980
rect 164332 29928 164384 29980
rect 171048 29928 171100 29980
rect 184296 29928 184348 29980
rect 188988 29928 189040 29980
rect 200120 29928 200172 29980
rect 204168 29928 204220 29980
rect 213828 29928 213880 29980
rect 215208 29928 215260 29980
rect 223396 29928 223448 29980
rect 227444 29928 227496 29980
rect 233884 29928 233936 29980
rect 523960 29928 524012 29980
rect 529296 29928 529348 29980
rect 44088 29860 44140 29912
rect 45468 29860 45520 29912
rect 72516 29860 72568 29912
rect 75828 29860 75880 29912
rect 98920 29860 98972 29912
rect 100668 29860 100720 29912
rect 121092 29860 121144 29912
rect 122748 29860 122800 29912
rect 141056 29860 141108 29912
rect 143448 29860 143500 29912
rect 158996 29860 159048 29912
rect 164148 29860 164200 29912
rect 178040 29860 178092 29912
rect 180708 29860 180760 29912
rect 192760 29860 192812 29912
rect 194508 29860 194560 29912
rect 205456 29860 205508 29912
rect 209688 29860 209740 29912
rect 218060 29860 218112 29912
rect 219348 29860 219400 29912
rect 227536 29860 227588 29912
rect 227628 29860 227680 29912
rect 234988 29860 235040 29912
rect 248328 29860 248380 29912
rect 252928 29860 252980 29912
rect 257988 29860 258040 29912
rect 261300 29860 261352 29912
rect 546132 29860 546184 29912
rect 556804 29860 556856 29912
rect 12256 29792 12308 29844
rect 41972 29792 42024 29844
rect 45376 29792 45428 29844
rect 6828 29724 6880 29776
rect 37740 29724 37792 29776
rect 45100 29724 45152 29776
rect 3976 29656 4028 29708
rect 35624 29656 35676 29708
rect 35808 29656 35860 29708
rect 42708 29656 42760 29708
rect 69388 29792 69440 29844
rect 70308 29792 70360 29844
rect 94688 29792 94740 29844
rect 96528 29792 96580 29844
rect 117872 29792 117924 29844
rect 118608 29792 118660 29844
rect 136824 29792 136876 29844
rect 137928 29792 137980 29844
rect 154764 29792 154816 29844
rect 157248 29792 157300 29844
rect 171692 29792 171744 29844
rect 172428 29792 172480 29844
rect 185400 29792 185452 29844
rect 187608 29792 187660 29844
rect 199108 29792 199160 29844
rect 201408 29792 201460 29844
rect 210700 29792 210752 29844
rect 212448 29792 212500 29844
rect 221280 29792 221332 29844
rect 222108 29792 222160 29844
rect 229652 29792 229704 29844
rect 530308 29792 530360 29844
rect 557540 29792 557592 29844
rect 67272 29724 67324 29776
rect 68928 29724 68980 29776
rect 92572 29724 92624 29776
rect 93768 29724 93820 29776
rect 114744 29724 114796 29776
rect 119896 29724 119948 29776
rect 138940 29724 138992 29776
rect 144736 29724 144788 29776
rect 161112 29724 161164 29776
rect 162768 29724 162820 29776
rect 176936 29724 176988 29776
rect 177856 29724 177908 29776
rect 189632 29724 189684 29776
rect 198648 29724 198700 29776
rect 208584 29724 208636 29776
rect 211068 29724 211120 29776
rect 220176 29724 220228 29776
rect 238668 29724 238720 29776
rect 244464 29724 244516 29776
rect 256608 29724 256660 29776
rect 260288 29724 260340 29776
rect 536656 29724 536708 29776
rect 564532 29724 564584 29776
rect 73620 29656 73672 29708
rect 78496 29656 78548 29708
rect 102048 29656 102100 29708
rect 107568 29656 107620 29708
rect 127348 29656 127400 29708
rect 136456 29656 136508 29708
rect 153752 29656 153804 29708
rect 161296 29656 161348 29708
rect 175924 29656 175976 29708
rect 177948 29656 178000 29708
rect 190644 29656 190696 29708
rect 194416 29656 194468 29708
rect 204352 29656 204404 29708
rect 208308 29656 208360 29708
rect 217048 29656 217100 29708
rect 219256 29656 219308 29708
rect 226524 29656 226576 29708
rect 229008 29656 229060 29708
rect 236000 29656 236052 29708
rect 237288 29656 237340 29708
rect 243360 29656 243412 29708
rect 246948 29656 247000 29708
rect 251824 29656 251876 29708
rect 508136 29656 508188 29708
rect 511356 29656 511408 29708
rect 514484 29656 514536 29708
rect 525064 29656 525116 29708
rect 539784 29656 539836 29708
rect 568580 29656 568632 29708
rect 5448 29588 5500 29640
rect 33048 29588 33100 29640
rect 44088 29588 44140 29640
rect 70400 29588 70452 29640
rect 71688 29588 71740 29640
rect 95700 29588 95752 29640
rect 100760 29588 100812 29640
rect 103152 29588 103204 29640
rect 103336 29588 103388 29640
rect 124220 29588 124272 29640
rect 128176 29588 128228 29640
rect 146392 29588 146444 29640
rect 153016 29588 153068 29640
rect 168472 29588 168524 29640
rect 169576 29588 169628 29640
rect 182180 29588 182232 29640
rect 186136 29588 186188 29640
rect 198004 29588 198056 29640
rect 202696 29588 202748 29640
rect 212816 29588 212868 29640
rect 213828 29588 213880 29640
rect 222292 29588 222344 29640
rect 235816 29588 235868 29640
rect 242348 29588 242400 29640
rect 498660 29588 498712 29640
rect 520924 29588 520976 29640
rect 20536 29520 20588 29572
rect 49332 29520 49384 29572
rect 49608 29520 49660 29572
rect 75736 29520 75788 29572
rect 81348 29520 81400 29572
rect 104164 29520 104216 29572
rect 104808 29520 104860 29572
rect 125232 29520 125284 29572
rect 125508 29520 125560 29572
rect 143172 29520 143224 29572
rect 144828 29520 144880 29572
rect 160100 29520 160152 29572
rect 165528 29520 165580 29572
rect 179052 29520 179104 29572
rect 186228 29520 186280 29572
rect 196992 29520 197044 29572
rect 235908 29520 235960 29572
rect 241244 29520 241296 29572
rect 542912 29520 542964 29572
rect 572812 29588 572864 29640
rect 28816 29452 28868 29504
rect 57796 29452 57848 29504
rect 57888 29452 57940 29504
rect 83096 29452 83148 29504
rect 86776 29452 86828 29504
rect 108396 29452 108448 29504
rect 31668 29384 31720 29436
rect 60924 29384 60976 29436
rect 64788 29384 64840 29436
rect 89444 29384 89496 29436
rect 91008 29384 91060 29436
rect 24768 29316 24820 29368
rect 53564 29316 53616 29368
rect 53748 29316 53800 29368
rect 79876 29316 79928 29368
rect 85488 29316 85540 29368
rect 107292 29384 107344 29436
rect 112628 29452 112680 29504
rect 114468 29452 114520 29504
rect 133696 29452 133748 29504
rect 140688 29452 140740 29504
rect 156880 29452 156932 29504
rect 160008 29452 160060 29504
rect 173808 29452 173860 29504
rect 176568 29452 176620 29504
rect 188528 29452 188580 29504
rect 191748 29452 191800 29504
rect 202236 29452 202288 29504
rect 266268 29452 266320 29504
rect 268752 29452 268804 29504
rect 110328 29384 110380 29436
rect 129464 29384 129516 29436
rect 129648 29384 129700 29436
rect 147404 29384 147456 29436
rect 153108 29384 153160 29436
rect 167460 29384 167512 29436
rect 169668 29384 169720 29436
rect 183284 29384 183336 29436
rect 184848 29384 184900 29436
rect 195796 29384 195848 29436
rect 106188 29316 106240 29368
rect 126336 29316 126388 29368
rect 126888 29316 126940 29368
rect 144276 29316 144328 29368
rect 150348 29316 150400 29368
rect 165344 29316 165396 29368
rect 19248 29248 19300 29300
rect 39948 29248 40000 29300
rect 61936 29248 61988 29300
rect 86224 29248 86276 29300
rect 95148 29248 95200 29300
rect 116860 29248 116912 29300
rect 28908 29180 28960 29232
rect 56692 29180 56744 29232
rect 60648 29180 60700 29232
rect 85212 29180 85264 29232
rect 97908 29180 97960 29232
rect 118976 29248 119028 29300
rect 121368 29248 121420 29300
rect 140044 29248 140096 29300
rect 142068 29248 142120 29300
rect 157984 29248 158036 29300
rect 161388 29248 161440 29300
rect 174820 29248 174872 29300
rect 234528 29248 234580 29300
rect 240232 29248 240284 29300
rect 267556 29248 267608 29300
rect 269764 29248 269816 29300
rect 117228 29180 117280 29232
rect 135812 29180 135864 29232
rect 136548 29180 136600 29232
rect 152648 29180 152700 29232
rect 241428 29180 241480 29232
rect 246580 29180 246632 29232
rect 249708 29180 249760 29232
rect 253940 29180 253992 29232
rect 262128 29180 262180 29232
rect 265532 29180 265584 29232
rect 270408 29180 270460 29232
rect 272892 29180 272944 29232
rect 26148 29112 26200 29164
rect 46848 29112 46900 29164
rect 74448 29112 74500 29164
rect 97816 29112 97868 29164
rect 103428 29112 103480 29164
rect 123116 29112 123168 29164
rect 135168 29112 135220 29164
rect 151636 29112 151688 29164
rect 151728 29112 151780 29164
rect 166356 29112 166408 29164
rect 210976 29112 211028 29164
rect 219164 29112 219216 29164
rect 230388 29112 230440 29164
rect 237104 29112 237156 29164
rect 240048 29112 240100 29164
rect 245476 29112 245528 29164
rect 245568 29112 245620 29164
rect 250812 29112 250864 29164
rect 252468 29112 252520 29164
rect 256056 29112 256108 29164
rect 260656 29112 260708 29164
rect 263416 29112 263468 29164
rect 264888 29112 264940 29164
rect 267648 29112 267700 29164
rect 271788 29112 271840 29164
rect 273996 29112 274048 29164
rect 274548 29112 274600 29164
rect 276112 29112 276164 29164
rect 277216 29112 277268 29164
rect 279240 29112 279292 29164
rect 281448 29112 281500 29164
rect 282460 29112 282512 29164
rect 289912 29112 289964 29164
rect 290832 29112 290884 29164
rect 296720 29112 296772 29164
rect 297180 29112 297232 29164
rect 299572 29112 299624 29164
rect 300308 29112 300360 29164
rect 305644 29112 305696 29164
rect 306288 29112 306340 29164
rect 306656 29112 306708 29164
rect 307668 29112 307720 29164
rect 309876 29112 309928 29164
rect 310428 29112 310480 29164
rect 310888 29112 310940 29164
rect 311808 29112 311860 29164
rect 316132 29112 316184 29164
rect 317328 29112 317380 29164
rect 318248 29112 318300 29164
rect 318708 29112 318760 29164
rect 320364 29112 320416 29164
rect 321284 29112 321336 29164
rect 323584 29112 323636 29164
rect 324228 29112 324280 29164
rect 327816 29112 327868 29164
rect 328368 29112 328420 29164
rect 328828 29112 328880 29164
rect 329748 29112 329800 29164
rect 329840 29112 329892 29164
rect 331128 29112 331180 29164
rect 331956 29112 332008 29164
rect 332508 29112 332560 29164
rect 333060 29112 333112 29164
rect 333888 29112 333940 29164
rect 334072 29112 334124 29164
rect 335084 29112 335136 29164
rect 336188 29112 336240 29164
rect 336648 29112 336700 29164
rect 337292 29112 337344 29164
rect 338028 29112 338080 29164
rect 338304 29112 338356 29164
rect 339316 29112 339368 29164
rect 341524 29112 341576 29164
rect 342168 29112 342220 29164
rect 342536 29112 342588 29164
rect 343548 29112 343600 29164
rect 345664 29112 345716 29164
rect 346308 29112 346360 29164
rect 346768 29112 346820 29164
rect 347688 29112 347740 29164
rect 351000 29112 351052 29164
rect 351828 29112 351880 29164
rect 352012 29112 352064 29164
rect 353208 29112 353260 29164
rect 354128 29112 354180 29164
rect 354588 29112 354640 29164
rect 356244 29112 356296 29164
rect 357256 29112 357308 29164
rect 359372 29112 359424 29164
rect 360108 29112 360160 29164
rect 360476 29112 360528 29164
rect 361396 29112 361448 29164
rect 363604 29112 363656 29164
rect 364248 29112 364300 29164
rect 364708 29112 364760 29164
rect 365628 29112 365680 29164
rect 365720 29112 365772 29164
rect 367008 29112 367060 29164
rect 367836 29112 367888 29164
rect 368388 29112 368440 29164
rect 368940 29112 368992 29164
rect 369768 29112 369820 29164
rect 369952 29112 370004 29164
rect 370964 29112 371016 29164
rect 372068 29112 372120 29164
rect 372528 29112 372580 29164
rect 373172 29112 373224 29164
rect 373908 29112 373960 29164
rect 374184 29112 374236 29164
rect 375288 29112 375340 29164
rect 377312 29112 377364 29164
rect 378048 29112 378100 29164
rect 378416 29112 378468 29164
rect 379244 29112 379296 29164
rect 381544 29112 381596 29164
rect 382188 29112 382240 29164
rect 382648 29112 382700 29164
rect 383568 29112 383620 29164
rect 386880 29112 386932 29164
rect 387708 29112 387760 29164
rect 387892 29112 387944 29164
rect 388904 29112 388956 29164
rect 390008 29112 390060 29164
rect 390468 29112 390520 29164
rect 391020 29112 391072 29164
rect 391848 29112 391900 29164
rect 392124 29112 392176 29164
rect 393044 29112 393096 29164
rect 395252 29112 395304 29164
rect 395988 29112 396040 29164
rect 396356 29112 396408 29164
rect 397276 29112 397328 29164
rect 399484 29112 399536 29164
rect 400128 29112 400180 29164
rect 400588 29112 400640 29164
rect 401508 29112 401560 29164
rect 403716 29112 403768 29164
rect 404268 29112 404320 29164
rect 404728 29112 404780 29164
rect 405648 29112 405700 29164
rect 407948 29112 408000 29164
rect 408408 29112 408460 29164
rect 408960 29112 409012 29164
rect 409788 29112 409840 29164
rect 410064 29112 410116 29164
rect 411168 29112 411220 29164
rect 414296 29112 414348 29164
rect 415124 29112 415176 29164
rect 417424 29112 417476 29164
rect 418068 29112 418120 29164
rect 418528 29112 418580 29164
rect 419448 29112 419500 29164
rect 419540 29112 419592 29164
rect 420828 29112 420880 29164
rect 421656 29112 421708 29164
rect 422208 29112 422260 29164
rect 422668 29112 422720 29164
rect 423588 29112 423640 29164
rect 423772 29112 423824 29164
rect 424968 29112 425020 29164
rect 425888 29112 425940 29164
rect 426348 29112 426400 29164
rect 426900 29112 426952 29164
rect 427728 29112 427780 29164
rect 428004 29112 428056 29164
rect 428924 29112 428976 29164
rect 435364 29112 435416 29164
rect 436008 29112 436060 29164
rect 436376 29112 436428 29164
rect 437388 29112 437440 29164
rect 437480 29112 437532 29164
rect 438768 29112 438820 29164
rect 439596 29112 439648 29164
rect 440148 29112 440200 29164
rect 440608 29112 440660 29164
rect 441528 29112 441580 29164
rect 441712 29112 441764 29164
rect 442908 29112 442960 29164
rect 443828 29112 443880 29164
rect 444288 29112 444340 29164
rect 444840 29112 444892 29164
rect 445668 29112 445720 29164
rect 445944 29112 445996 29164
rect 446864 29112 446916 29164
rect 449072 29112 449124 29164
rect 449808 29112 449860 29164
rect 450084 29112 450136 29164
rect 451096 29112 451148 29164
rect 453304 29112 453356 29164
rect 453948 29112 454000 29164
rect 454316 29112 454368 29164
rect 455328 29112 455380 29164
rect 455420 29112 455472 29164
rect 456708 29112 456760 29164
rect 457536 29112 457588 29164
rect 458088 29112 458140 29164
rect 458548 29112 458600 29164
rect 459468 29112 459520 29164
rect 461768 29112 461820 29164
rect 462228 29112 462280 29164
rect 462780 29112 462832 29164
rect 463608 29112 463660 29164
rect 463792 29112 463844 29164
rect 464988 29112 465040 29164
rect 465908 29112 465960 29164
rect 466368 29112 466420 29164
rect 467012 29112 467064 29164
rect 467748 29112 467800 29164
rect 468024 29112 468076 29164
rect 469036 29112 469088 29164
rect 471244 29112 471296 29164
rect 471888 29112 471940 29164
rect 472256 29112 472308 29164
rect 473268 29112 473320 29164
rect 473360 29112 473412 29164
rect 475384 29112 475436 29164
rect 475476 29112 475528 29164
rect 476028 29112 476080 29164
rect 476488 29112 476540 29164
rect 477408 29112 477460 29164
rect 477592 29112 477644 29164
rect 478788 29112 478840 29164
rect 479616 29112 479668 29164
rect 480168 29112 480220 29164
rect 480720 29112 480772 29164
rect 481548 29112 481600 29164
rect 481732 29112 481784 29164
rect 482928 29112 482980 29164
rect 483848 29112 483900 29164
rect 484308 29112 484360 29164
rect 484952 29112 485004 29164
rect 485688 29112 485740 29164
rect 485964 29112 486016 29164
rect 486976 29112 487028 29164
rect 489184 29112 489236 29164
rect 489828 29112 489880 29164
rect 490196 29112 490248 29164
rect 491208 29112 491260 29164
rect 491300 29112 491352 29164
rect 492588 29112 492640 29164
rect 493324 29112 493376 29164
rect 493968 29112 494020 29164
rect 494428 29112 494480 29164
rect 495348 29112 495400 29164
rect 495440 29112 495492 29164
rect 497464 29112 497516 29164
rect 497556 29112 497608 29164
rect 498108 29112 498160 29164
rect 499672 29112 499724 29164
rect 500684 29112 500736 29164
rect 501788 29112 501840 29164
rect 502248 29112 502300 29164
rect 502892 29112 502944 29164
rect 503628 29112 503680 29164
rect 503904 29112 503956 29164
rect 504824 29112 504876 29164
rect 507124 29112 507176 29164
rect 507768 29112 507820 29164
rect 511264 29112 511316 29164
rect 511908 29112 511960 29164
rect 512368 29112 512420 29164
rect 513288 29112 513340 29164
rect 513380 29112 513432 29164
rect 514668 29112 514720 29164
rect 515496 29112 515548 29164
rect 516048 29112 516100 29164
rect 516600 29112 516652 29164
rect 517428 29112 517480 29164
rect 517612 29112 517664 29164
rect 518624 29112 518676 29164
rect 519728 29112 519780 29164
rect 520188 29112 520240 29164
rect 520832 29112 520884 29164
rect 521568 29112 521620 29164
rect 521844 29112 521896 29164
rect 522948 29112 523000 29164
rect 524972 29112 525024 29164
rect 525708 29112 525760 29164
rect 531320 29112 531372 29164
rect 532608 29112 532660 29164
rect 533436 29112 533488 29164
rect 533988 29112 534040 29164
rect 534540 29112 534592 29164
rect 535368 29112 535420 29164
rect 535552 29112 535604 29164
rect 536748 29112 536800 29164
rect 537668 29112 537720 29164
rect 538128 29112 538180 29164
rect 538680 29112 538732 29164
rect 539508 29112 539560 29164
rect 544016 29112 544068 29164
rect 544936 29112 544988 29164
rect 548248 29112 548300 29164
rect 549168 29112 549220 29164
rect 9588 28976 9640 29028
rect 39856 29044 39908 29096
rect 59912 29044 59964 29096
rect 95056 29044 95108 29096
rect 115756 29044 115808 29096
rect 115848 29044 115900 29096
rect 134800 29044 134852 29096
rect 139308 29044 139360 29096
rect 155868 29044 155920 29096
rect 220728 29044 220780 29096
rect 228640 29044 228692 29096
rect 242808 29044 242860 29096
rect 247592 29044 247644 29096
rect 251088 29044 251140 29096
rect 255044 29044 255096 29096
rect 259368 29044 259420 29096
rect 262404 29044 262456 29096
rect 263508 29044 263560 29096
rect 266636 29044 266688 29096
rect 269028 29044 269080 29096
rect 270776 29044 270828 29096
rect 273904 29044 273956 29096
rect 275008 29044 275060 29096
rect 278688 29044 278740 29096
rect 280344 29044 280396 29096
rect 311992 29044 312044 29096
rect 313280 29044 313332 29096
rect 319352 29044 319404 29096
rect 321560 29044 321612 29096
rect 324596 29044 324648 29096
rect 325608 29044 325660 29096
rect 347780 29044 347832 29096
rect 348976 29044 349028 29096
rect 355232 29044 355284 29096
rect 355968 29044 356020 29096
rect 383660 29044 383712 29096
rect 384856 29044 384908 29096
rect 405832 29044 405884 29096
rect 406936 29044 406988 29096
rect 413192 29044 413244 29096
rect 413928 29044 413980 29096
rect 431132 29044 431184 29096
rect 431868 29044 431920 29096
rect 432236 29044 432288 29096
rect 433064 29044 433116 29096
rect 492312 29044 492364 29096
rect 493416 29044 493468 29096
rect 526076 29044 526128 29096
rect 526904 29044 526956 29096
rect 547144 29044 547196 29096
rect 547788 29044 547840 29096
rect 549260 29044 549312 29096
rect 550456 29044 550508 29096
rect 37188 28976 37240 29028
rect 64052 28976 64104 29028
rect 99288 28976 99340 29028
rect 119712 28976 119764 29028
rect 119804 28976 119856 29028
rect 137836 28976 137888 29028
rect 231768 28976 231820 29028
rect 238116 28976 238168 29028
rect 252376 28976 252428 29028
rect 257068 28976 257120 29028
rect 260748 28976 260800 29028
rect 264520 28976 264572 29028
rect 268936 28976 268988 29028
rect 271880 28976 271932 29028
rect 282828 28976 282880 29028
rect 283472 28976 283524 29028
rect 314108 28976 314160 29028
rect 314568 28976 314620 29028
rect 325700 28976 325752 29028
rect 327724 28976 327776 29028
rect 343640 28976 343692 29028
rect 344836 28976 344888 29028
rect 349896 28976 349948 29028
rect 350448 28976 350500 29028
rect 385776 28976 385828 29028
rect 386328 28976 386380 29028
rect 401600 28976 401652 29028
rect 402796 28976 402848 29028
rect 459652 28976 459704 29028
rect 460756 28976 460808 29028
rect 529204 28976 529256 29028
rect 529848 28976 529900 29028
rect 66168 28568 66220 28620
rect 90456 28568 90508 28620
rect 52368 28500 52420 28552
rect 77760 28500 77812 28552
rect 79968 28500 80020 28552
rect 100760 28500 100812 28552
rect 30288 28432 30340 28484
rect 58808 28432 58860 28484
rect 59268 28432 59320 28484
rect 84108 28432 84160 28484
rect 17868 28364 17920 28416
rect 47216 28364 47268 28416
rect 48228 28364 48280 28416
rect 74632 28364 74684 28416
rect 77208 28364 77260 28416
rect 99932 28364 99984 28416
rect 22008 28296 22060 28348
rect 51448 28296 51500 28348
rect 55128 28296 55180 28348
rect 80980 28296 81032 28348
rect 84108 28296 84160 28348
rect 106280 28296 106332 28348
rect 8208 28228 8260 28280
rect 38752 28228 38804 28280
rect 41328 28228 41380 28280
rect 68284 28228 68336 28280
rect 73068 28228 73120 28280
rect 96804 28228 96856 28280
rect 51724 27616 51776 27668
rect 55680 27616 55732 27668
rect 60832 26732 60884 26784
rect 62028 26732 62080 26784
rect 3424 20612 3476 20664
rect 18604 20612 18656 20664
rect 552664 20612 552716 20664
rect 579988 20612 580040 20664
rect 299572 11704 299624 11756
rect 300768 11704 300820 11756
rect 3424 6808 3476 6860
rect 15844 6808 15896 6860
rect 555424 6808 555476 6860
rect 580172 6808 580224 6860
rect 69112 6128 69164 6180
rect 93584 6128 93636 6180
rect 526996 6128 527048 6180
rect 554964 6128 555016 6180
rect 62212 5244 62264 5296
rect 65156 5244 65208 5296
rect 475384 5244 475436 5296
rect 494704 5244 494756 5296
rect 511356 5244 511408 5296
rect 533712 5244 533764 5296
rect 493416 5176 493468 5228
rect 515956 5176 516008 5228
rect 471336 5108 471388 5160
rect 491116 5108 491168 5160
rect 497464 5108 497516 5160
rect 519544 5108 519596 5160
rect 525064 5108 525116 5160
rect 540796 5108 540848 5160
rect 477408 5040 477460 5092
rect 498200 5040 498252 5092
rect 502248 5040 502300 5092
rect 526628 5040 526680 5092
rect 529296 5040 529348 5092
rect 551468 5040 551520 5092
rect 8116 4972 8168 5024
rect 31760 4972 31812 5024
rect 486976 4972 487028 5024
rect 508872 4972 508924 5024
rect 511908 4972 511960 5024
rect 537208 4972 537260 5024
rect 8024 4904 8076 4956
rect 33508 4904 33560 4956
rect 33600 4904 33652 4956
rect 60832 4904 60884 4956
rect 467748 4904 467800 4956
rect 487620 4904 487672 4956
rect 489828 4904 489880 4956
rect 512460 4904 512512 4956
rect 518624 4904 518676 4956
rect 544384 4904 544436 4956
rect 12348 4836 12400 4888
rect 42984 4836 43036 4888
rect 482836 4836 482888 4888
rect 505376 4836 505428 4888
rect 521568 4836 521620 4888
rect 547880 4836 547932 4888
rect 556804 4836 556856 4888
rect 576308 4836 576360 4888
rect 2872 4768 2924 4820
rect 34520 4768 34572 4820
rect 62120 4768 62172 4820
rect 87328 4768 87380 4820
rect 480168 4768 480220 4820
rect 501788 4768 501840 4820
rect 504916 4768 504968 4820
rect 530124 4768 530176 4820
rect 533988 4768 534040 4820
rect 562048 4768 562100 4820
rect 520924 4156 520976 4208
rect 523040 4156 523092 4208
rect 314568 4088 314620 4140
rect 316224 4088 316276 4140
rect 325608 4088 325660 4140
rect 328000 4088 328052 4140
rect 342168 4088 342220 4140
rect 346952 4088 347004 4140
rect 350448 4088 350500 4140
rect 356336 4088 356388 4140
rect 358728 4088 358780 4140
rect 365812 4088 365864 4140
rect 382188 4088 382240 4140
rect 391848 4088 391900 4140
rect 397276 4088 397328 4140
rect 408408 4088 408460 4140
rect 413928 4088 413980 4140
rect 427268 4088 427320 4140
rect 430488 4088 430540 4140
rect 446220 4088 446272 4140
rect 455328 4088 455380 4140
rect 473452 4088 473504 4140
rect 481548 4088 481600 4140
rect 502984 4088 503036 4140
rect 503628 4088 503680 4140
rect 527824 4088 527876 4140
rect 538128 4088 538180 4140
rect 566832 4088 566884 4140
rect 340788 4020 340840 4072
rect 345756 4020 345808 4072
rect 375288 4020 375340 4072
rect 383476 4020 383528 4072
rect 384856 4020 384908 4072
rect 394240 4020 394292 4072
rect 394608 4020 394660 4072
rect 406016 4020 406068 4072
rect 411168 4020 411220 4072
rect 423772 4020 423824 4072
rect 424968 4020 425020 4072
rect 439136 4020 439188 4072
rect 440148 4020 440200 4072
rect 456892 4020 456944 4072
rect 460756 4020 460808 4072
rect 479340 4020 479392 4072
rect 487068 4020 487120 4072
rect 510068 4020 510120 4072
rect 513288 4020 513340 4072
rect 538404 4020 538456 4072
rect 544936 4020 544988 4072
rect 573916 4020 573968 4072
rect 333888 3952 333940 4004
rect 337476 3952 337528 4004
rect 353208 3952 353260 4004
rect 358728 3952 358780 4004
rect 369768 3952 369820 4004
rect 377680 3952 377732 4004
rect 383568 3952 383620 4004
rect 392952 3952 393004 4004
rect 393044 3952 393096 4004
rect 403624 3952 403676 4004
rect 404268 3952 404320 4004
rect 416688 3952 416740 4004
rect 418068 3952 418120 4004
rect 432052 3952 432104 4004
rect 433064 3952 433116 4004
rect 448612 3952 448664 4004
rect 451188 3952 451240 4004
rect 469864 3952 469916 4004
rect 476028 3952 476080 4004
rect 497096 3952 497148 4004
rect 506388 3952 506440 4004
rect 531320 3952 531372 4004
rect 532516 3952 532568 4004
rect 560852 3952 560904 4004
rect 373908 3884 373960 3936
rect 382372 3884 382424 3936
rect 387708 3884 387760 3936
rect 397736 3884 397788 3936
rect 398748 3884 398800 3936
rect 410800 3884 410852 3936
rect 416596 3884 416648 3936
rect 430856 3884 430908 3936
rect 436008 3884 436060 3936
rect 452108 3884 452160 3936
rect 452568 3884 452620 3936
rect 471060 3884 471112 3936
rect 478696 3884 478748 3936
rect 500592 3884 500644 3936
rect 509148 3884 509200 3936
rect 534908 3884 534960 3936
rect 542268 3884 542320 3936
rect 571524 3884 571576 3936
rect 367008 3816 367060 3868
rect 374092 3816 374144 3868
rect 376668 3816 376720 3868
rect 385960 3816 386012 3868
rect 386328 3816 386380 3868
rect 396540 3816 396592 3868
rect 397368 3816 397420 3868
rect 344928 3748 344980 3800
rect 350448 3748 350500 3800
rect 351828 3748 351880 3800
rect 357532 3748 357584 3800
rect 361396 3748 361448 3800
rect 368204 3748 368256 3800
rect 378048 3748 378100 3800
rect 387156 3748 387208 3800
rect 389088 3748 389140 3800
rect 354588 3680 354640 3732
rect 361120 3680 361172 3732
rect 361488 3680 361540 3732
rect 369400 3680 369452 3732
rect 372528 3680 372580 3732
rect 381176 3680 381228 3732
rect 384948 3680 385000 3732
rect 395344 3680 395396 3732
rect 400128 3680 400180 3732
rect 402888 3816 402940 3868
rect 415492 3816 415544 3868
rect 422208 3816 422260 3868
rect 436744 3816 436796 3868
rect 437388 3816 437440 3868
rect 453304 3816 453356 3868
rect 456616 3816 456668 3868
rect 475752 3816 475804 3868
rect 491208 3816 491260 3868
rect 513564 3816 513616 3868
rect 517428 3816 517480 3868
rect 543188 3816 543240 3868
rect 545028 3816 545080 3868
rect 575112 3816 575164 3868
rect 400312 3748 400364 3800
rect 411904 3748 411956 3800
rect 412548 3748 412600 3800
rect 426164 3748 426216 3800
rect 428924 3748 428976 3800
rect 443828 3748 443880 3800
rect 444288 3748 444340 3800
rect 461584 3748 461636 3800
rect 462228 3748 462280 3800
rect 481732 3748 481784 3800
rect 492588 3748 492640 3800
rect 514760 3748 514812 3800
rect 516048 3748 516100 3800
rect 541992 3748 542044 3800
rect 549168 3748 549220 3800
rect 578608 3748 578660 3800
rect 409604 3680 409656 3732
rect 409788 3680 409840 3732
rect 422576 3680 422628 3732
rect 423588 3680 423640 3732
rect 437940 3680 437992 3732
rect 442816 3680 442868 3732
rect 460388 3680 460440 3732
rect 466368 3680 466420 3732
rect 486424 3680 486476 3732
rect 488448 3680 488500 3732
rect 511264 3680 511316 3732
rect 514668 3680 514720 3732
rect 539600 3680 539652 3732
rect 547788 3680 547840 3732
rect 577412 3680 577464 3732
rect 324228 3612 324280 3664
rect 326804 3612 326856 3664
rect 332508 3612 332560 3664
rect 336280 3612 336332 3664
rect 357348 3612 357400 3664
rect 364616 3612 364668 3664
rect 370964 3612 371016 3664
rect 378876 3612 378928 3664
rect 379244 3612 379296 3664
rect 388260 3612 388312 3664
rect 393228 3612 393280 3664
rect 404820 3612 404872 3664
rect 407028 3612 407080 3664
rect 420184 3612 420236 3664
rect 420736 3612 420788 3664
rect 435548 3612 435600 3664
rect 438676 3612 438728 3664
rect 455696 3612 455748 3664
rect 460848 3612 460900 3664
rect 480536 3612 480588 3664
rect 484308 3612 484360 3664
rect 506480 3612 506532 3664
rect 510528 3612 510580 3664
rect 536104 3612 536156 3664
rect 540888 3612 540940 3664
rect 570328 3612 570380 3664
rect 27712 3544 27764 3596
rect 28816 3544 28868 3596
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12256 3476 12308 3528
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 25320 3476 25372 3528
rect 26148 3476 26200 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 51724 3544 51776 3596
rect 26516 3408 26568 3460
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 51356 3476 51408 3528
rect 52368 3476 52420 3528
rect 52552 3476 52604 3528
rect 53656 3476 53708 3528
rect 34796 3408 34848 3460
rect 35808 3408 35860 3460
rect 35992 3408 36044 3460
rect 37188 3408 37240 3460
rect 40684 3408 40736 3460
rect 41328 3408 41380 3460
rect 41880 3408 41932 3460
rect 42708 3408 42760 3460
rect 43076 3408 43128 3460
rect 44088 3408 44140 3460
rect 44272 3408 44324 3460
rect 45376 3408 45428 3460
rect 48964 3408 49016 3460
rect 49608 3408 49660 3460
rect 19432 3272 19484 3324
rect 20536 3272 20588 3324
rect 37188 3272 37240 3324
rect 62212 3544 62264 3596
rect 77392 3544 77444 3596
rect 78496 3544 78548 3596
rect 307760 3544 307812 3596
rect 309048 3544 309100 3596
rect 326988 3544 327040 3596
rect 330392 3544 330444 3596
rect 335268 3544 335320 3596
rect 339868 3544 339920 3596
rect 353116 3544 353168 3596
rect 359924 3544 359976 3596
rect 362868 3544 362920 3596
rect 370596 3544 370648 3596
rect 371148 3544 371200 3596
rect 379980 3544 380032 3596
rect 380808 3544 380860 3596
rect 390652 3544 390704 3596
rect 401508 3544 401560 3596
rect 413100 3544 413152 3596
rect 415216 3544 415268 3596
rect 429660 3544 429712 3596
rect 433156 3544 433208 3596
rect 449808 3544 449860 3596
rect 451096 3544 451148 3596
rect 468668 3544 468720 3596
rect 469036 3544 469088 3596
rect 488816 3544 488868 3596
rect 495348 3544 495400 3596
rect 518348 3544 518400 3596
rect 518808 3544 518860 3596
rect 545488 3544 545540 3596
rect 550548 3544 550600 3596
rect 582196 3544 582248 3596
rect 56048 3476 56100 3528
rect 56508 3476 56560 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 60832 3476 60884 3528
rect 62028 3476 62080 3528
rect 64328 3476 64380 3528
rect 64788 3476 64840 3528
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 66720 3476 66772 3528
rect 67548 3476 67600 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 82084 3476 82136 3528
rect 82728 3476 82780 3528
rect 83280 3476 83332 3528
rect 84108 3476 84160 3528
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 92388 3476 92440 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 105728 3476 105780 3528
rect 106188 3476 106240 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 109316 3476 109368 3528
rect 110328 3476 110380 3528
rect 110512 3476 110564 3528
rect 111524 3476 111576 3528
rect 114008 3476 114060 3528
rect 114468 3476 114520 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 116400 3476 116452 3528
rect 117228 3476 117280 3528
rect 117596 3476 117648 3528
rect 118608 3476 118660 3528
rect 122288 3476 122340 3528
rect 122748 3476 122800 3528
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 125876 3476 125928 3528
rect 126888 3476 126940 3528
rect 126980 3476 127032 3528
rect 128268 3476 128320 3528
rect 130568 3476 130620 3528
rect 131028 3476 131080 3528
rect 132960 3476 133012 3528
rect 133788 3476 133840 3528
rect 134156 3476 134208 3528
rect 135168 3476 135220 3528
rect 138848 3476 138900 3528
rect 139308 3476 139360 3528
rect 140044 3476 140096 3528
rect 140688 3476 140740 3528
rect 141240 3476 141292 3528
rect 142068 3476 142120 3528
rect 142436 3476 142488 3528
rect 143448 3476 143500 3528
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 149520 3476 149572 3528
rect 150348 3476 150400 3528
rect 151820 3476 151872 3528
rect 153108 3476 153160 3528
rect 156604 3476 156656 3528
rect 157248 3476 157300 3528
rect 157800 3476 157852 3528
rect 158628 3476 158680 3528
rect 158904 3476 158956 3528
rect 160008 3476 160060 3528
rect 160100 3476 160152 3528
rect 161388 3476 161440 3528
rect 163688 3476 163740 3528
rect 164148 3476 164200 3528
rect 164884 3476 164936 3528
rect 165528 3476 165580 3528
rect 166080 3476 166132 3528
rect 166908 3476 166960 3528
rect 167184 3476 167236 3528
rect 168288 3476 168340 3528
rect 171968 3476 172020 3528
rect 172428 3476 172480 3528
rect 173164 3476 173216 3528
rect 173808 3476 173860 3528
rect 174268 3476 174320 3528
rect 175188 3476 175240 3528
rect 175464 3476 175516 3528
rect 176568 3476 176620 3528
rect 176660 3476 176712 3528
rect 177764 3476 177816 3528
rect 180248 3476 180300 3528
rect 180708 3476 180760 3528
rect 181444 3476 181496 3528
rect 182088 3476 182140 3528
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 184940 3476 184992 3528
rect 186228 3476 186280 3528
rect 188528 3476 188580 3528
rect 188988 3476 189040 3528
rect 190828 3476 190880 3528
rect 191748 3476 191800 3528
rect 192024 3476 192076 3528
rect 193128 3476 193180 3528
rect 193220 3476 193272 3528
rect 194324 3476 194376 3528
rect 197912 3476 197964 3528
rect 198648 3476 198700 3528
rect 199108 3476 199160 3528
rect 200028 3476 200080 3528
rect 201500 3476 201552 3528
rect 202788 3476 202840 3528
rect 205088 3476 205140 3528
rect 205548 3476 205600 3528
rect 206192 3476 206244 3528
rect 206928 3476 206980 3528
rect 207388 3476 207440 3528
rect 208308 3476 208360 3528
rect 209780 3476 209832 3528
rect 210884 3476 210936 3528
rect 213368 3476 213420 3528
rect 213828 3476 213880 3528
rect 214472 3476 214524 3528
rect 215208 3476 215260 3528
rect 215668 3476 215720 3528
rect 216588 3476 216640 3528
rect 216864 3476 216916 3528
rect 217968 3476 218020 3528
rect 218060 3476 218112 3528
rect 219164 3476 219216 3528
rect 222752 3476 222804 3528
rect 223488 3476 223540 3528
rect 223948 3476 224000 3528
rect 224868 3476 224920 3528
rect 229836 3476 229888 3528
rect 230388 3476 230440 3528
rect 231032 3476 231084 3528
rect 231768 3476 231820 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 234620 3476 234672 3528
rect 235908 3476 235960 3528
rect 238116 3476 238168 3528
rect 238668 3476 238720 3528
rect 239312 3476 239364 3528
rect 240048 3476 240100 3528
rect 240508 3476 240560 3528
rect 241428 3476 241480 3528
rect 242900 3476 242952 3528
rect 244004 3476 244056 3528
rect 247592 3476 247644 3528
rect 248328 3476 248380 3528
rect 249984 3476 250036 3528
rect 251088 3476 251140 3528
rect 251180 3476 251232 3528
rect 252468 3476 252520 3528
rect 254676 3476 254728 3528
rect 255228 3476 255280 3528
rect 255872 3476 255924 3528
rect 256608 3476 256660 3528
rect 257068 3476 257120 3528
rect 257988 3476 258040 3528
rect 264152 3476 264204 3528
rect 264888 3476 264940 3528
rect 265348 3476 265400 3528
rect 266268 3476 266320 3528
rect 266544 3476 266596 3528
rect 267556 3476 267608 3528
rect 267740 3476 267792 3528
rect 269028 3476 269080 3528
rect 273628 3476 273680 3528
rect 274548 3476 274600 3528
rect 276020 3476 276072 3528
rect 277308 3476 277360 3528
rect 280712 3476 280764 3528
rect 281448 3476 281500 3528
rect 281908 3476 281960 3528
rect 282828 3476 282880 3528
rect 283104 3476 283156 3528
rect 284576 3476 284628 3528
rect 285404 3476 285456 3528
rect 286600 3476 286652 3528
rect 288992 3476 289044 3528
rect 289728 3476 289780 3528
rect 291384 3476 291436 3528
rect 291936 3476 291988 3528
rect 301412 3476 301464 3528
rect 301964 3476 302016 3528
rect 303528 3476 303580 3528
rect 304356 3476 304408 3528
rect 304908 3476 304960 3528
rect 305552 3476 305604 3528
rect 310428 3476 310480 3528
rect 311440 3476 311492 3528
rect 311808 3476 311860 3528
rect 312636 3476 312688 3528
rect 318708 3476 318760 3528
rect 320916 3476 320968 3528
rect 321284 3476 321336 3528
rect 323308 3476 323360 3528
rect 327724 3476 327776 3528
rect 329196 3476 329248 3528
rect 331128 3476 331180 3528
rect 333888 3476 333940 3528
rect 335084 3476 335136 3528
rect 338672 3476 338724 3528
rect 339408 3476 339460 3528
rect 344560 3476 344612 3528
rect 344836 3476 344888 3528
rect 349252 3476 349304 3528
rect 357256 3476 357308 3528
rect 363512 3476 363564 3528
rect 364248 3476 364300 3528
rect 371700 3476 371752 3528
rect 375196 3476 375248 3528
rect 384764 3476 384816 3528
rect 388904 3476 388956 3528
rect 398932 3476 398984 3528
rect 402796 3476 402848 3528
rect 414296 3476 414348 3528
rect 415124 3476 415176 3528
rect 428464 3476 428516 3528
rect 429108 3476 429160 3528
rect 445024 3476 445076 3528
rect 446864 3476 446916 3528
rect 463976 3476 464028 3528
rect 464896 3476 464948 3528
rect 485228 3476 485280 3528
rect 493968 3476 494020 3528
rect 517152 3476 517204 3528
rect 520188 3476 520240 3528
rect 546684 3476 546736 3528
rect 551928 3476 551980 3528
rect 583392 3476 583444 3528
rect 57244 3408 57296 3460
rect 57888 3408 57940 3460
rect 102232 3408 102284 3460
rect 103428 3408 103480 3460
rect 106924 3408 106976 3460
rect 107568 3408 107620 3460
rect 131764 3408 131816 3460
rect 132408 3408 132460 3460
rect 189724 3408 189776 3460
rect 190368 3408 190420 3460
rect 272432 3408 272484 3460
rect 273904 3408 273956 3460
rect 279516 3408 279568 3460
rect 281356 3408 281408 3460
rect 328368 3408 328420 3460
rect 331588 3408 331640 3460
rect 338028 3408 338080 3460
rect 342168 3408 342220 3460
rect 343548 3408 343600 3460
rect 348056 3408 348108 3460
rect 348976 3408 349028 3460
rect 354036 3408 354088 3460
rect 366916 3408 366968 3460
rect 375288 3408 375340 3460
rect 379336 3408 379388 3460
rect 389456 3408 389508 3460
rect 395988 3408 396040 3460
rect 407212 3408 407264 3460
rect 411076 3408 411128 3460
rect 424968 3408 425020 3460
rect 434628 3408 434680 3460
rect 331036 3340 331088 3392
rect 335084 3340 335136 3392
rect 390468 3340 390520 3392
rect 401324 3340 401376 3392
rect 408316 3340 408368 3392
rect 421380 3340 421432 3392
rect 424876 3340 424928 3392
rect 440332 3340 440384 3392
rect 447048 3408 447100 3460
rect 465172 3408 465224 3460
rect 469128 3408 469180 3460
rect 489920 3408 489972 3460
rect 498108 3408 498160 3460
rect 521844 3408 521896 3460
rect 522856 3408 522908 3460
rect 550272 3408 550324 3460
rect 550456 3408 550508 3460
rect 581000 3408 581052 3460
rect 450912 3340 450964 3392
rect 453948 3340 454000 3392
rect 472256 3340 472308 3392
rect 474648 3340 474700 3392
rect 495900 3340 495952 3392
rect 496728 3340 496780 3392
rect 520740 3340 520792 3392
rect 535368 3340 535420 3392
rect 563244 3340 563296 3392
rect 80888 3272 80940 3324
rect 81348 3272 81400 3324
rect 85672 3272 85724 3324
rect 86776 3272 86828 3324
rect 89168 3272 89220 3324
rect 89628 3272 89680 3324
rect 93952 3272 94004 3324
rect 95056 3272 95108 3324
rect 97448 3272 97500 3324
rect 97908 3272 97960 3324
rect 196808 3272 196860 3324
rect 197268 3272 197320 3324
rect 221556 3272 221608 3324
rect 222108 3272 222160 3324
rect 262956 3272 263008 3324
rect 263508 3272 263560 3324
rect 271236 3272 271288 3324
rect 271788 3272 271840 3324
rect 287796 3272 287848 3324
rect 288348 3272 288400 3324
rect 317328 3272 317380 3324
rect 318524 3272 318576 3324
rect 339316 3272 339368 3324
rect 343364 3272 343416 3324
rect 347688 3272 347740 3324
rect 352840 3272 352892 3324
rect 355968 3272 356020 3324
rect 362316 3272 362368 3324
rect 391756 3272 391808 3324
rect 402520 3272 402572 3324
rect 406936 3272 406988 3324
rect 418988 3272 419040 3324
rect 426348 3272 426400 3324
rect 441528 3272 441580 3324
rect 445668 3272 445720 3324
rect 462780 3272 462832 3324
rect 473268 3272 473320 3324
rect 493508 3272 493560 3324
rect 500868 3272 500920 3324
rect 525432 3272 525484 3324
rect 528468 3272 528520 3324
rect 556160 3272 556212 3324
rect 101036 3204 101088 3256
rect 102048 3204 102100 3256
rect 183744 3204 183796 3256
rect 184848 3204 184900 3256
rect 200304 3204 200356 3256
rect 201408 3204 201460 3256
rect 225144 3204 225196 3256
rect 226248 3204 226300 3256
rect 258264 3204 258316 3256
rect 259368 3204 259420 3256
rect 336648 3204 336700 3256
rect 340972 3204 341024 3256
rect 346308 3204 346360 3256
rect 351644 3204 351696 3256
rect 405648 3204 405700 3256
rect 417884 3204 417936 3256
rect 420828 3204 420880 3256
rect 434444 3204 434496 3256
rect 441436 3204 441488 3256
rect 458088 3204 458140 3256
rect 464988 3204 465040 3256
rect 484032 3204 484084 3256
rect 485688 3204 485740 3256
rect 507676 3204 507728 3256
rect 507768 3204 507820 3256
rect 532516 3204 532568 3256
rect 539508 3204 539560 3256
rect 568028 3204 568080 3256
rect 241704 3136 241756 3188
rect 242808 3136 242860 3188
rect 321376 3136 321428 3188
rect 324412 3136 324464 3188
rect 329748 3136 329800 3188
rect 332692 3136 332744 3188
rect 419448 3136 419500 3188
rect 433248 3136 433300 3188
rect 438768 3136 438820 3188
rect 454500 3136 454552 3188
rect 457996 3136 458048 3188
rect 476948 3136 477000 3188
rect 482928 3136 482980 3188
rect 504180 3136 504232 3188
rect 504824 3136 504876 3188
rect 529020 3136 529072 3188
rect 536748 3136 536800 3188
rect 564440 3136 564492 3188
rect 118792 3068 118844 3120
rect 119804 3068 119856 3120
rect 246396 3068 246448 3120
rect 246948 3068 247000 3120
rect 360108 3068 360160 3120
rect 367008 3068 367060 3120
rect 368388 3068 368440 3120
rect 376484 3068 376536 3120
rect 427728 3068 427780 3120
rect 442632 3068 442684 3120
rect 442908 3068 442960 3120
rect 459192 3068 459244 3120
rect 459468 3068 459520 3120
rect 478144 3068 478196 3120
rect 478788 3068 478840 3120
rect 499396 3068 499448 3120
rect 500684 3068 500736 3120
rect 524236 3068 524288 3120
rect 532608 3068 532660 3120
rect 559748 3068 559800 3120
rect 150624 3000 150676 3052
rect 151728 3000 151780 3052
rect 168380 3000 168432 3052
rect 169484 3000 169536 3052
rect 208584 3000 208636 3052
rect 209688 3000 209740 3052
rect 226340 3000 226392 3052
rect 227444 3000 227496 3052
rect 248788 3000 248840 3052
rect 249708 3000 249760 3052
rect 259460 3000 259512 3052
rect 260564 3000 260616 3052
rect 274824 3000 274876 3052
rect 277032 3000 277084 3052
rect 284300 3000 284352 3052
rect 285588 3000 285640 3052
rect 302424 3000 302476 3052
rect 303160 3000 303212 3052
rect 317236 3000 317288 3052
rect 319720 3000 319772 3052
rect 322848 3000 322900 3052
rect 325608 3000 325660 3052
rect 431868 3000 431920 3052
rect 447416 3000 447468 3052
rect 448428 3000 448480 3052
rect 466276 3000 466328 3052
rect 471888 3000 471940 3052
rect 492312 3000 492364 3052
rect 525708 3000 525760 3052
rect 552664 3000 552716 3052
rect 73804 2932 73856 2984
rect 74448 2932 74500 2984
rect 313188 2932 313240 2984
rect 315028 2932 315080 2984
rect 463608 2932 463660 2984
rect 482836 2932 482888 2984
rect 526904 2932 526956 2984
rect 553768 2932 553820 2984
rect 572 2864 624 2916
rect 8116 2864 8168 2916
rect 135260 2864 135312 2916
rect 136548 2864 136600 2916
rect 349068 2864 349120 2916
rect 355232 2864 355284 2916
rect 365628 2864 365680 2916
rect 372896 2864 372948 2916
rect 456708 2864 456760 2916
rect 474556 2864 474608 2916
rect 529848 2864 529900 2916
rect 557356 2864 557408 2916
rect 1676 2796 1728 2848
rect 8024 2796 8076 2848
rect 449716 2796 449768 2848
rect 467472 2796 467524 2848
rect 522948 2796 523000 2848
rect 549076 2796 549128 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700670 73016 703520
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 105464 699718 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 170324 699718 170352 703520
rect 202800 700126 202828 703520
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 218992 700058 219020 703520
rect 218980 700052 219032 700058
rect 218980 699994 219032 700000
rect 235184 699854 235212 703520
rect 257988 700868 258040 700874
rect 257988 700810 258040 700816
rect 244188 700596 244240 700602
rect 244188 700538 244240 700544
rect 235172 699848 235224 699854
rect 235172 699790 235224 699796
rect 238024 699848 238076 699854
rect 238024 699790 238076 699796
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 106200 675646 106228 699654
rect 171060 675782 171088 699654
rect 230388 696992 230440 696998
rect 230388 696934 230440 696940
rect 171048 675776 171100 675782
rect 171048 675718 171100 675724
rect 106188 675640 106240 675646
rect 106188 675582 106240 675588
rect 175556 675504 175608 675510
rect 175556 675446 175608 675452
rect 157340 675436 157392 675442
rect 157340 675378 157392 675384
rect 143632 675368 143684 675374
rect 143632 675310 143684 675316
rect 130016 675300 130068 675306
rect 130016 675242 130068 675248
rect 25596 675232 25648 675238
rect 25596 675174 25648 675180
rect 7564 674960 7616 674966
rect 7564 674902 7616 674908
rect 4802 673840 4858 673849
rect 4802 673775 4858 673784
rect 3516 673328 3568 673334
rect 3516 673270 3568 673276
rect 3424 672104 3476 672110
rect 3424 672046 3476 672052
rect 3332 671560 3384 671566
rect 3332 671502 3384 671508
rect 3344 671265 3372 671502
rect 3330 671256 3386 671265
rect 3330 671191 3386 671200
rect 3332 658232 3384 658238
rect 3330 658200 3332 658209
rect 3384 658200 3386 658209
rect 3330 658135 3386 658144
rect 3332 633412 3384 633418
rect 3332 633354 3384 633360
rect 3344 632097 3372 633354
rect 3330 632088 3386 632097
rect 3330 632023 3386 632032
rect 3332 619608 3384 619614
rect 3332 619550 3384 619556
rect 3344 619177 3372 619550
rect 3330 619168 3386 619177
rect 3330 619103 3386 619112
rect 3056 607164 3108 607170
rect 3056 607106 3108 607112
rect 3068 606121 3096 607106
rect 3054 606112 3110 606121
rect 3054 606047 3110 606056
rect 3332 580984 3384 580990
rect 3332 580926 3384 580932
rect 3344 580009 3372 580926
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3148 567112 3200 567118
rect 3148 567054 3200 567060
rect 3160 566953 3188 567054
rect 3146 566944 3202 566953
rect 3146 566879 3202 566888
rect 2964 554736 3016 554742
rect 2964 554678 3016 554684
rect 2976 553897 3004 554678
rect 2962 553888 3018 553897
rect 2962 553823 3018 553832
rect 3148 528556 3200 528562
rect 3148 528498 3200 528504
rect 3160 527921 3188 528498
rect 3146 527912 3202 527921
rect 3146 527847 3202 527856
rect 2964 502308 3016 502314
rect 2964 502250 3016 502256
rect 2976 501809 3004 502250
rect 2962 501800 3018 501809
rect 2962 501735 3018 501744
rect 3240 476060 3292 476066
rect 3240 476002 3292 476008
rect 3252 475697 3280 476002
rect 3238 475688 3294 475697
rect 3238 475623 3294 475632
rect 3056 463684 3108 463690
rect 3056 463626 3108 463632
rect 3068 462641 3096 463626
rect 3054 462632 3110 462641
rect 3054 462567 3110 462576
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3332 293956 3384 293962
rect 3332 293898 3384 293904
rect 3344 293185 3372 293898
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3436 149841 3464 672046
rect 3528 254153 3556 673270
rect 3608 672036 3660 672042
rect 3608 671978 3660 671984
rect 3620 514865 3648 671978
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150476 3568 150482
rect 3516 150418 3568 150424
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3424 137964 3476 137970
rect 3424 137906 3476 137912
rect 3436 136785 3464 137906
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3528 97617 3556 150418
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71664 3476 71670
rect 3422 71632 3424 71641
rect 3476 71632 3478 71641
rect 3422 71567 3478 71576
rect 4816 58682 4844 673775
rect 4896 673532 4948 673538
rect 4896 673474 4948 673480
rect 4908 150482 4936 673474
rect 4896 150476 4948 150482
rect 4896 150418 4948 150424
rect 7576 71670 7604 674902
rect 14556 674552 14608 674558
rect 14556 674494 14608 674500
rect 11796 674008 11848 674014
rect 11796 673950 11848 673956
rect 7748 673192 7800 673198
rect 7748 673134 7800 673140
rect 7656 671424 7708 671430
rect 7656 671366 7708 671372
rect 7668 567118 7696 671366
rect 7760 633418 7788 673134
rect 10324 671084 10376 671090
rect 10324 671026 10376 671032
rect 7748 633412 7800 633418
rect 7748 633354 7800 633360
rect 7656 567112 7708 567118
rect 7656 567054 7708 567060
rect 10336 306338 10364 671026
rect 11702 670032 11758 670041
rect 11702 669967 11758 669976
rect 10414 669760 10470 669769
rect 10414 669695 10470 669704
rect 10428 554742 10456 669695
rect 10416 554736 10468 554742
rect 10416 554678 10468 554684
rect 10324 306332 10376 306338
rect 10324 306274 10376 306280
rect 7564 71664 7616 71670
rect 7564 71606 7616 71612
rect 2780 58676 2832 58682
rect 2780 58618 2832 58624
rect 4804 58676 4856 58682
rect 4804 58618 4856 58624
rect 2792 58585 2820 58618
rect 2778 58576 2834 58585
rect 2778 58511 2834 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 11716 33114 11744 669967
rect 11808 358766 11836 673950
rect 11888 673056 11940 673062
rect 11888 672998 11940 673004
rect 11900 580990 11928 672998
rect 14464 671016 14516 671022
rect 14464 670958 14516 670964
rect 11888 580984 11940 580990
rect 11888 580926 11940 580932
rect 11796 358760 11848 358766
rect 11796 358702 11848 358708
rect 14476 189038 14504 670958
rect 14568 502314 14596 674494
rect 17316 674212 17368 674218
rect 17316 674154 17368 674160
rect 17224 673736 17276 673742
rect 15842 673704 15898 673713
rect 17224 673678 17276 673684
rect 15842 673639 15898 673648
rect 14648 672920 14700 672926
rect 14648 672862 14700 672868
rect 14660 528562 14688 672862
rect 14648 528556 14700 528562
rect 14648 528498 14700 528504
rect 14556 502308 14608 502314
rect 14556 502250 14608 502256
rect 14464 189032 14516 189038
rect 14464 188974 14516 188980
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 11704 33108 11756 33114
rect 11704 33050 11756 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 10968 30116 11020 30122
rect 10968 30058 11020 30064
rect 6828 29776 6880 29782
rect 6828 29718 6880 29724
rect 3976 29708 4028 29714
rect 3976 29650 4028 29656
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3988 16574 4016 29650
rect 5448 29640 5500 29646
rect 5448 29582 5500 29588
rect 3988 16546 4108 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 584 480 612 2858
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1688 480 1716 2790
rect 2884 480 2912 4762
rect 4080 480 4108 16546
rect 5460 6914 5488 29582
rect 6840 6914 6868 29718
rect 9588 29028 9640 29034
rect 9588 28970 9640 28976
rect 8208 28280 8260 28286
rect 8208 28222 8260 28228
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8024 4956 8076 4962
rect 8024 4898 8076 4904
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 480 7696 3470
rect 8036 2854 8064 4898
rect 8128 2922 8156 4966
rect 8220 3534 8248 28222
rect 9600 3534 9628 28970
rect 10980 3534 11008 30058
rect 13728 29980 13780 29986
rect 13728 29922 13780 29928
rect 12256 29844 12308 29850
rect 12256 29786 12308 29792
rect 12268 3534 12296 29786
rect 13740 6914 13768 29922
rect 15108 29912 15160 29918
rect 15108 29854 15160 29860
rect 15120 6914 15148 29854
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12348 4888 12400 4894
rect 12348 4830 12400 4836
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 12360 480 12388 4830
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 15856 6866 15884 673639
rect 16028 672852 16080 672858
rect 16028 672794 16080 672800
rect 15936 671288 15988 671294
rect 15936 671230 15988 671236
rect 15948 449886 15976 671230
rect 16040 476066 16068 672794
rect 16028 476060 16080 476066
rect 16028 476002 16080 476008
rect 15936 449880 15988 449886
rect 15936 449822 15988 449828
rect 17236 202842 17264 673678
rect 17328 398818 17356 674154
rect 18696 674076 18748 674082
rect 18696 674018 18748 674024
rect 17408 672716 17460 672722
rect 17408 672658 17460 672664
rect 17420 423638 17448 672658
rect 18602 669896 18658 669905
rect 18602 669831 18658 669840
rect 17408 423632 17460 423638
rect 17408 423574 17460 423580
rect 17316 398812 17368 398818
rect 17316 398754 17368 398760
rect 17224 202836 17276 202842
rect 17224 202778 17276 202784
rect 16488 30252 16540 30258
rect 16488 30194 16540 30200
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 16500 3534 16528 30194
rect 17868 28416 17920 28422
rect 17868 28358 17920 28364
rect 17880 3534 17908 28358
rect 18616 20670 18644 669831
rect 18708 346390 18736 674018
rect 22744 673668 22796 673674
rect 22744 673610 22796 673616
rect 18788 672580 18840 672586
rect 18788 672522 18840 672528
rect 18800 372570 18828 672522
rect 21456 672512 21508 672518
rect 21456 672454 21508 672460
rect 21364 671152 21416 671158
rect 21364 671094 21416 671100
rect 18788 372564 18840 372570
rect 18788 372506 18840 372512
rect 18696 346384 18748 346390
rect 18696 346326 18748 346332
rect 21376 293962 21404 671094
rect 21468 320142 21496 672454
rect 21456 320136 21508 320142
rect 21456 320078 21508 320084
rect 21364 293956 21416 293962
rect 21364 293898 21416 293904
rect 22756 137970 22784 673610
rect 25504 673600 25556 673606
rect 25504 673542 25556 673548
rect 22836 672376 22888 672382
rect 22836 672318 22888 672324
rect 22848 215286 22876 672318
rect 22836 215280 22888 215286
rect 22836 215222 22888 215228
rect 22744 137964 22796 137970
rect 22744 137906 22796 137912
rect 25516 85542 25544 673542
rect 25608 164218 25636 675174
rect 29736 675164 29788 675170
rect 29736 675106 29788 675112
rect 26884 674280 26936 674286
rect 26884 674222 26936 674228
rect 26896 411262 26924 674222
rect 27068 671968 27120 671974
rect 27068 671910 27120 671916
rect 26976 671764 27028 671770
rect 26976 671706 27028 671712
rect 26988 619614 27016 671706
rect 27080 658238 27108 671910
rect 28356 671900 28408 671906
rect 28356 671842 28408 671848
rect 28264 671356 28316 671362
rect 28264 671298 28316 671304
rect 27068 658232 27120 658238
rect 27068 658174 27120 658180
rect 26976 619608 27028 619614
rect 26976 619550 27028 619556
rect 28276 463690 28304 671298
rect 28368 607170 28396 671842
rect 29642 670712 29698 670721
rect 29642 670647 29698 670656
rect 28356 607164 28408 607170
rect 28356 607106 28408 607112
rect 28264 463684 28316 463690
rect 28264 463626 28316 463632
rect 26884 411256 26936 411262
rect 26884 411198 26936 411204
rect 25596 164212 25648 164218
rect 25596 164154 25648 164160
rect 25504 85536 25556 85542
rect 25504 85478 25556 85484
rect 29656 45558 29684 670647
rect 29748 111790 29776 675106
rect 75276 675096 75328 675102
rect 75276 675038 75328 675044
rect 43352 675028 43404 675034
rect 43352 674970 43404 674976
rect 31024 673872 31076 673878
rect 31024 673814 31076 673820
rect 31036 241466 31064 673814
rect 31116 672444 31168 672450
rect 31116 672386 31168 672392
rect 31128 267714 31156 672386
rect 34242 672208 34298 672217
rect 34242 672143 34298 672152
rect 34256 671908 34284 672143
rect 43364 671908 43392 674970
rect 52460 674892 52512 674898
rect 52460 674834 52512 674840
rect 47858 672344 47914 672353
rect 47858 672279 47914 672288
rect 47872 671908 47900 672279
rect 52472 671908 52500 674834
rect 61568 672172 61620 672178
rect 61568 672114 61620 672120
rect 61580 671908 61608 672114
rect 75288 671908 75316 675038
rect 125416 674688 125468 674694
rect 125416 674630 125468 674636
rect 111708 674348 111760 674354
rect 111708 674290 111760 674296
rect 107200 673804 107252 673810
rect 107200 673746 107252 673752
rect 98092 672308 98144 672314
rect 98092 672250 98144 672256
rect 84384 672240 84436 672246
rect 84384 672182 84436 672188
rect 84396 671908 84424 672182
rect 98104 671908 98132 672250
rect 107212 671908 107240 673746
rect 111720 671908 111748 674290
rect 120908 673940 120960 673946
rect 120908 673882 120960 673888
rect 120920 671908 120948 673882
rect 125428 671908 125456 674630
rect 130028 671908 130056 675242
rect 139124 672648 139176 672654
rect 139124 672590 139176 672596
rect 139136 671908 139164 672590
rect 143644 671908 143672 675310
rect 152832 674756 152884 674762
rect 152832 674698 152884 674704
rect 148232 674144 148284 674150
rect 148232 674086 148284 674092
rect 148244 671908 148272 674086
rect 152844 671908 152872 674698
rect 155776 674348 155828 674354
rect 155776 674290 155828 674296
rect 155788 672790 155816 674290
rect 155776 672784 155828 672790
rect 155776 672726 155828 672732
rect 157352 671908 157380 675378
rect 166448 674416 166500 674422
rect 166448 674358 166500 674364
rect 161940 674348 161992 674354
rect 161940 674290 161992 674296
rect 161952 671908 161980 674290
rect 166460 671908 166488 674358
rect 171048 672988 171100 672994
rect 171048 672930 171100 672936
rect 171060 671908 171088 672930
rect 175568 671908 175596 675446
rect 218060 674824 218112 674830
rect 218060 674766 218112 674772
rect 200120 674620 200172 674626
rect 200120 674562 200172 674568
rect 180156 674484 180208 674490
rect 180156 674426 180208 674432
rect 180168 671908 180196 674426
rect 200132 673334 200160 674562
rect 212080 673396 212132 673402
rect 212080 673338 212132 673344
rect 200120 673328 200172 673334
rect 200120 673270 200172 673276
rect 198372 673260 198424 673266
rect 198372 673202 198424 673208
rect 184756 673124 184808 673130
rect 184756 673066 184808 673072
rect 184768 671908 184796 673066
rect 198384 671908 198412 673202
rect 212092 671908 212120 673338
rect 218072 672042 218100 674766
rect 225788 673328 225840 673334
rect 225788 673270 225840 673276
rect 218060 672036 218112 672042
rect 218060 671978 218112 671984
rect 221464 672036 221516 672042
rect 221464 671978 221516 671984
rect 221476 671922 221504 671978
rect 221214 671894 221504 671922
rect 225800 671908 225828 673270
rect 230400 671922 230428 696934
rect 235908 683256 235960 683262
rect 235908 683198 235960 683204
rect 235920 673454 235948 683198
rect 238036 675918 238064 699790
rect 238024 675912 238076 675918
rect 238024 675854 238076 675860
rect 239496 675572 239548 675578
rect 239496 675514 239548 675520
rect 235368 673426 235948 673454
rect 235368 671922 235396 673426
rect 230322 671894 230428 671922
rect 234922 671894 235396 671922
rect 239508 671908 239536 675514
rect 244200 671922 244228 700538
rect 249708 700528 249760 700534
rect 249708 700470 249760 700476
rect 249720 673454 249748 700470
rect 253112 675844 253164 675850
rect 253112 675786 253164 675792
rect 248984 673426 249748 673454
rect 248984 671922 249012 673426
rect 244030 671894 244228 671922
rect 248630 671894 249012 671922
rect 253124 671908 253152 675786
rect 258000 671922 258028 700810
rect 263508 700800 263560 700806
rect 263508 700742 263560 700748
rect 263520 673454 263548 700742
rect 267660 699854 267688 703520
rect 275928 700256 275980 700262
rect 275928 700198 275980 700204
rect 271788 700188 271840 700194
rect 271788 700130 271840 700136
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 266820 675708 266872 675714
rect 266820 675650 266872 675656
rect 262600 673426 263548 673454
rect 262600 671922 262628 673426
rect 257738 671894 258028 671922
rect 262246 671894 262628 671922
rect 266832 671908 266860 675650
rect 271800 671922 271828 700130
rect 271446 671894 271828 671922
rect 275940 671908 275968 700198
rect 283852 699786 283880 703520
rect 289728 699984 289780 699990
rect 289728 699926 289780 699932
rect 285588 699916 285640 699922
rect 285588 699858 285640 699864
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 280528 675980 280580 675986
rect 280528 675922 280580 675928
rect 280540 671908 280568 675922
rect 285600 673454 285628 699858
rect 285416 673426 285628 673454
rect 285416 671922 285444 673426
rect 289740 671922 289768 699926
rect 298100 699848 298152 699854
rect 298100 699790 298152 699796
rect 298112 692774 298140 699790
rect 298112 692746 298416 692774
rect 294236 676048 294288 676054
rect 294236 675990 294288 675996
rect 285062 671894 285444 671922
rect 289662 671894 289768 671922
rect 294248 671908 294276 675990
rect 298388 671922 298416 692746
rect 299492 676054 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 329840 701004 329892 701010
rect 329840 700946 329892 700952
rect 325700 700936 325752 700942
rect 325700 700878 325752 700884
rect 311900 700120 311952 700126
rect 311900 700062 311952 700068
rect 302240 699780 302292 699786
rect 302240 699722 302292 699728
rect 302252 692774 302280 699722
rect 311912 692774 311940 700062
rect 316040 700052 316092 700058
rect 316040 699994 316092 700000
rect 316052 692774 316080 699994
rect 325712 692774 325740 700878
rect 329852 692774 329880 700946
rect 332520 699922 332548 703520
rect 343640 700732 343692 700738
rect 343640 700674 343692 700680
rect 339500 700664 339552 700670
rect 339500 700606 339552 700612
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 302252 692746 303016 692774
rect 311912 692746 312032 692774
rect 316052 692746 316632 692774
rect 325712 692746 325832 692774
rect 329852 692746 330248 692774
rect 299480 676048 299532 676054
rect 299480 675990 299532 675996
rect 302988 671922 303016 692746
rect 307852 675912 307904 675918
rect 307852 675854 307904 675860
rect 298388 671894 298770 671922
rect 302988 671894 303370 671922
rect 307864 671908 307892 675854
rect 312004 671922 312032 692746
rect 316604 671922 316632 692746
rect 321560 675776 321612 675782
rect 321560 675718 321612 675724
rect 312004 671894 312478 671922
rect 316604 671894 316986 671922
rect 321572 671908 321600 675718
rect 325804 671922 325832 692746
rect 330220 671922 330248 692746
rect 335268 675640 335320 675646
rect 335268 675582 335320 675588
rect 325804 671894 326186 671922
rect 330220 671894 330694 671922
rect 335280 671908 335308 675582
rect 339512 671922 339540 700606
rect 343652 692774 343680 700674
rect 347872 700460 347924 700466
rect 347872 700402 347924 700408
rect 347884 692774 347912 700402
rect 348804 699990 348832 703520
rect 364996 700466 365024 703520
rect 349804 700460 349856 700466
rect 349804 700402 349856 700408
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 343652 692746 344048 692774
rect 347884 692746 348464 692774
rect 344020 671922 344048 692746
rect 348436 671922 348464 692746
rect 349816 675986 349844 700402
rect 357440 700392 357492 700398
rect 357440 700334 357492 700340
rect 353300 700324 353352 700330
rect 353300 700266 353352 700272
rect 356704 700324 356756 700330
rect 356704 700266 356756 700272
rect 349804 675980 349856 675986
rect 349804 675922 349856 675928
rect 353312 671922 353340 700266
rect 356716 675850 356744 700266
rect 357452 692774 357480 700334
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 357452 692746 357664 692774
rect 356704 675844 356756 675850
rect 356704 675786 356756 675792
rect 357636 671922 357664 692746
rect 361580 683188 361632 683194
rect 361580 683130 361632 683136
rect 361592 673454 361620 683130
rect 429212 675714 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 494808 700330 494836 703520
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 559668 699718 559696 703520
rect 555424 699712 555476 699718
rect 555424 699654 555476 699660
rect 559656 699712 559708 699718
rect 559656 699654 559708 699660
rect 429200 675708 429252 675714
rect 429200 675650 429252 675656
rect 555436 675578 555464 699654
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 555424 675572 555476 675578
rect 555424 675514 555476 675520
rect 554136 675504 554188 675510
rect 554136 675446 554188 675452
rect 499488 675232 499540 675238
rect 499488 675174 499540 675180
rect 412824 674824 412876 674830
rect 412824 674766 412876 674772
rect 382280 674756 382332 674762
rect 382280 674698 382332 674704
rect 368664 674688 368716 674694
rect 368664 674630 368716 674636
rect 361592 673426 362264 673454
rect 362236 671922 362264 673426
rect 368676 671974 368704 674630
rect 376300 673192 376352 673198
rect 376300 673134 376352 673140
rect 367284 671968 367336 671974
rect 339512 671894 339802 671922
rect 344020 671894 344402 671922
rect 348436 671894 348910 671922
rect 353312 671894 353510 671922
rect 357636 671894 358110 671922
rect 362236 671894 362618 671922
rect 367218 671916 367284 671922
rect 367218 671910 367336 671916
rect 368664 671968 368716 671974
rect 368664 671910 368716 671916
rect 367218 671894 367324 671910
rect 376312 671908 376340 673134
rect 380926 671906 381032 671922
rect 380926 671900 381044 671906
rect 380926 671894 380992 671900
rect 380992 671842 381044 671848
rect 217048 671832 217100 671838
rect 216706 671780 217048 671786
rect 216706 671774 217100 671780
rect 216706 671758 217088 671774
rect 207848 671696 207900 671702
rect 202998 671634 203288 671650
rect 207598 671644 207848 671650
rect 207598 671638 207900 671644
rect 202998 671628 203300 671634
rect 202998 671622 203248 671628
rect 207598 671622 207888 671638
rect 203248 671570 203300 671576
rect 382292 671566 382320 674698
rect 408224 674552 408276 674558
rect 408224 674494 408276 674500
rect 390008 673056 390060 673062
rect 390008 672998 390060 673004
rect 390020 671908 390048 672998
rect 403624 672920 403676 672926
rect 403624 672862 403676 672868
rect 403636 671908 403664 672862
rect 408236 671908 408264 674494
rect 412836 671908 412864 674766
rect 481180 674620 481232 674626
rect 481180 674562 481232 674568
rect 440148 674280 440200 674286
rect 440148 674222 440200 674228
rect 435548 674212 435600 674218
rect 435548 674154 435600 674160
rect 417332 672852 417384 672858
rect 417332 672794 417384 672800
rect 417344 671908 417372 672794
rect 431040 672716 431092 672722
rect 431040 672658 431092 672664
rect 431052 671908 431080 672658
rect 435560 671908 435588 674154
rect 440160 671908 440188 674222
rect 449256 674076 449308 674082
rect 449256 674018 449308 674024
rect 444748 672580 444800 672586
rect 444748 672522 444800 672528
rect 444760 671908 444788 672522
rect 449268 671908 449296 674018
rect 453856 674008 453908 674014
rect 453856 673950 453908 673956
rect 453868 671908 453896 673950
rect 476672 673872 476724 673878
rect 476672 673814 476724 673820
rect 458364 672512 458416 672518
rect 458364 672454 458416 672460
rect 458376 671908 458404 672454
rect 472072 672444 472124 672450
rect 472072 672386 472124 672392
rect 472084 671908 472112 672386
rect 476684 671908 476712 673814
rect 481192 671908 481220 674562
rect 494888 673736 494940 673742
rect 494888 673678 494940 673684
rect 485780 672376 485832 672382
rect 485780 672318 485832 672324
rect 485792 671908 485820 672318
rect 494900 671908 494928 673678
rect 499500 671908 499528 675174
rect 513104 675164 513156 675170
rect 513104 675106 513156 675112
rect 503996 673668 504048 673674
rect 503996 673610 504048 673616
rect 504008 671908 504036 673610
rect 508596 672104 508648 672110
rect 508596 672046 508648 672052
rect 508608 671908 508636 672046
rect 513116 671908 513144 675106
rect 552664 675028 552716 675034
rect 552664 674970 552716 674976
rect 526812 674960 526864 674966
rect 526812 674902 526864 674908
rect 517704 673600 517756 673606
rect 517704 673542 517756 673548
rect 517716 671908 517744 673542
rect 522212 673532 522264 673538
rect 522212 673474 522264 673480
rect 522224 671908 522252 673474
rect 526824 671908 526852 674902
rect 535918 673840 535974 673849
rect 535918 673775 535974 673784
rect 535932 671908 535960 673775
rect 545026 673704 545082 673713
rect 545026 673639 545082 673648
rect 545040 671908 545068 673639
rect 385144 671770 385434 671786
rect 421576 671770 421958 671786
rect 385132 671764 385434 671770
rect 385184 671758 385434 671764
rect 421564 671764 421958 671770
rect 385132 671706 385184 671712
rect 421616 671758 421958 671764
rect 421564 671706 421616 671712
rect 371332 671560 371384 671566
rect 66194 671498 66300 671514
rect 70702 671498 70992 671514
rect 79810 671498 80008 671514
rect 93518 671498 93716 671514
rect 134550 671498 134840 671514
rect 193890 671498 194272 671514
rect 382280 671560 382332 671566
rect 371384 671508 371726 671514
rect 371332 671502 371726 671508
rect 382280 671502 382332 671508
rect 66194 671492 66312 671498
rect 66194 671486 66260 671492
rect 70702 671492 71004 671498
rect 70702 671486 70952 671492
rect 66260 671434 66312 671440
rect 79810 671492 80020 671498
rect 79810 671486 79968 671492
rect 70952 671434 71004 671440
rect 93518 671492 93728 671498
rect 93518 671486 93676 671492
rect 79968 671434 80020 671440
rect 134550 671492 134852 671498
rect 134550 671486 134800 671492
rect 93676 671434 93728 671440
rect 193890 671492 194284 671498
rect 193890 671486 194232 671492
rect 134800 671434 134852 671440
rect 371344 671486 371726 671502
rect 194232 671434 194284 671440
rect 398840 671424 398892 671430
rect 39026 671392 39082 671401
rect 38778 671350 39026 671378
rect 57334 671392 57390 671401
rect 56994 671350 57334 671378
rect 39026 671327 39082 671336
rect 89074 671392 89130 671401
rect 88918 671350 89074 671378
rect 57334 671327 57390 671336
rect 102874 671392 102930 671401
rect 102626 671350 102874 671378
rect 89074 671327 89130 671336
rect 116490 671392 116546 671401
rect 116334 671350 116490 671378
rect 102874 671327 102930 671336
rect 189630 671392 189686 671401
rect 189290 671350 189630 671378
rect 116490 671327 116546 671336
rect 189630 671327 189686 671336
rect 394146 671392 394202 671401
rect 394202 671350 394542 671378
rect 426256 671424 426308 671430
rect 398892 671372 399142 671378
rect 398840 671366 399142 671372
rect 462596 671424 462648 671430
rect 426308 671372 426466 671378
rect 426256 671366 426466 671372
rect 467196 671424 467248 671430
rect 462648 671372 462990 671378
rect 462596 671366 462990 671372
rect 490104 671424 490156 671430
rect 467248 671372 467590 671378
rect 467196 671366 467590 671372
rect 531226 671392 531282 671401
rect 490156 671372 490314 671378
rect 490104 671366 490314 671372
rect 398852 671350 399142 671366
rect 426268 671350 426466 671366
rect 462608 671350 462990 671366
rect 467208 671350 467590 671366
rect 490116 671350 490314 671366
rect 394146 671327 394202 671336
rect 540334 671392 540390 671401
rect 531282 671350 531438 671378
rect 531226 671327 531282 671336
rect 549350 671392 549406 671401
rect 540390 671350 540546 671378
rect 540334 671327 540390 671336
rect 549406 671350 549654 671378
rect 549350 671327 549406 671336
rect 31116 267708 31168 267714
rect 31116 267650 31168 267656
rect 31024 241460 31076 241466
rect 31024 241402 31076 241408
rect 29736 111784 29788 111790
rect 29736 111726 29788 111732
rect 29644 45552 29696 45558
rect 29644 45494 29696 45500
rect 31772 32014 32522 32042
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20536 29572 20588 29578
rect 20536 29514 20588 29520
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 18604 20664 18656 20670
rect 18604 20606 18656 20612
rect 19260 3534 19288 29242
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 15948 480 15976 3470
rect 17052 480 17080 3470
rect 18248 480 18276 3470
rect 20548 3330 20576 29514
rect 19432 3324 19484 3330
rect 19432 3266 19484 3272
rect 20536 3324 20588 3330
rect 20536 3266 20588 3272
rect 19444 480 19472 3266
rect 20640 480 20668 30262
rect 23388 30184 23440 30190
rect 23388 30126 23440 30132
rect 22008 28348 22060 28354
rect 22008 28290 22060 28296
rect 22020 6914 22048 28290
rect 23400 6914 23428 30126
rect 28816 29504 28868 29510
rect 28816 29446 28868 29452
rect 24768 29368 24820 29374
rect 24768 29310 24820 29316
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3534 24808 29310
rect 26148 29164 26200 29170
rect 26148 29106 26200 29112
rect 26160 3534 26188 29106
rect 28828 16574 28856 29446
rect 31668 29436 31720 29442
rect 31668 29378 31720 29384
rect 28908 29232 28960 29238
rect 28908 29174 28960 29180
rect 28736 16546 28856 16574
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 24228 480 24256 3470
rect 25332 480 25360 3470
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 26528 480 26556 3402
rect 27724 480 27752 3538
rect 28736 3482 28764 16546
rect 28920 6914 28948 29174
rect 30288 28484 30340 28490
rect 30288 28426 30340 28432
rect 30300 6914 30328 28426
rect 31680 6914 31708 29378
rect 28828 6886 28948 6914
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 28828 3602 28856 6886
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 28736 3454 28948 3482
rect 28920 480 28948 3454
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 31772 5030 31800 32014
rect 33048 29640 33100 29646
rect 33048 29582 33100 29588
rect 31760 5024 31812 5030
rect 31760 4966 31812 4972
rect 33060 3534 33088 29582
rect 33520 4962 33548 32028
rect 33508 4956 33560 4962
rect 33508 4898 33560 4904
rect 33600 4956 33652 4962
rect 33600 4898 33652 4904
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 32416 480 32444 3470
rect 33612 480 33640 4898
rect 34532 4826 34560 32028
rect 35636 29714 35664 32028
rect 36648 30054 36676 32028
rect 36636 30048 36688 30054
rect 36636 29990 36688 29996
rect 37752 29782 37780 32028
rect 38568 30048 38620 30054
rect 38568 29990 38620 29996
rect 37740 29776 37792 29782
rect 37740 29718 37792 29724
rect 35624 29708 35676 29714
rect 35624 29650 35676 29656
rect 35808 29708 35860 29714
rect 35808 29650 35860 29656
rect 34520 4820 34572 4826
rect 34520 4762 34572 4768
rect 35820 3466 35848 29650
rect 37188 29028 37240 29034
rect 37188 28970 37240 28976
rect 37200 3466 37228 28970
rect 38580 6914 38608 29990
rect 38764 28286 38792 32028
rect 39868 29102 39896 32028
rect 40880 30138 40908 32028
rect 40960 30252 41012 30258
rect 40960 30194 41012 30200
rect 40788 30122 40908 30138
rect 40776 30116 40908 30122
rect 40828 30110 40908 30116
rect 40776 30058 40828 30064
rect 40972 29986 41000 30194
rect 40960 29980 41012 29986
rect 40960 29922 41012 29928
rect 41984 29850 42012 32028
rect 41972 29844 42024 29850
rect 41972 29786 42024 29792
rect 42708 29708 42760 29714
rect 42708 29650 42760 29656
rect 39948 29300 40000 29306
rect 39948 29242 40000 29248
rect 39856 29096 39908 29102
rect 39856 29038 39908 29044
rect 38752 28280 38804 28286
rect 38752 28222 38804 28228
rect 39960 6914 39988 29242
rect 41328 28280 41380 28286
rect 41328 28222 41380 28228
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 34796 3460 34848 3466
rect 34796 3402 34848 3408
rect 35808 3460 35860 3466
rect 35808 3402 35860 3408
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 37188 3460 37240 3466
rect 37188 3402 37240 3408
rect 34808 480 34836 3402
rect 36004 480 36032 3402
rect 37188 3324 37240 3330
rect 37188 3266 37240 3272
rect 37200 480 37228 3266
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3466 41368 28222
rect 42720 3466 42748 29650
rect 42996 4894 43024 32028
rect 44100 29918 44128 32028
rect 44088 29912 44140 29918
rect 44088 29854 44140 29860
rect 45112 29782 45140 32028
rect 46216 29986 46244 32028
rect 46204 29980 46256 29986
rect 46204 29922 46256 29928
rect 45468 29912 45520 29918
rect 45468 29854 45520 29860
rect 45376 29844 45428 29850
rect 45376 29786 45428 29792
rect 45100 29776 45152 29782
rect 45100 29718 45152 29724
rect 44088 29640 44140 29646
rect 44088 29582 44140 29588
rect 42984 4888 43036 4894
rect 42984 4830 43036 4836
rect 44100 3466 44128 29582
rect 45388 3466 45416 29786
rect 40684 3460 40736 3466
rect 40684 3402 40736 3408
rect 41328 3460 41380 3466
rect 41328 3402 41380 3408
rect 41880 3460 41932 3466
rect 41880 3402 41932 3408
rect 42708 3460 42760 3466
rect 42708 3402 42760 3408
rect 43076 3460 43128 3466
rect 43076 3402 43128 3408
rect 44088 3460 44140 3466
rect 44088 3402 44140 3408
rect 44272 3460 44324 3466
rect 44272 3402 44324 3408
rect 45376 3460 45428 3466
rect 45376 3402 45428 3408
rect 40696 480 40724 3402
rect 41892 480 41920 3402
rect 43088 480 43116 3402
rect 44284 480 44312 3402
rect 45480 480 45508 29854
rect 46848 29164 46900 29170
rect 46848 29106 46900 29112
rect 46860 6914 46888 29106
rect 47228 28422 47256 32028
rect 48240 30258 48268 32028
rect 48228 30252 48280 30258
rect 48228 30194 48280 30200
rect 49344 29578 49372 32028
rect 50356 30326 50384 32028
rect 50344 30320 50396 30326
rect 50344 30262 50396 30268
rect 50988 30320 51040 30326
rect 50988 30262 51040 30268
rect 49332 29572 49384 29578
rect 49332 29514 49384 29520
rect 49608 29572 49660 29578
rect 49608 29514 49660 29520
rect 47216 28416 47268 28422
rect 47216 28358 47268 28364
rect 48228 28416 48280 28422
rect 48228 28358 48280 28364
rect 48240 6914 48268 28358
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3466 49648 29514
rect 51000 3534 51028 30262
rect 51460 28354 51488 32028
rect 52472 30190 52500 32028
rect 52460 30184 52512 30190
rect 52460 30126 52512 30132
rect 53576 29374 53604 32028
rect 54588 30258 54616 32028
rect 54576 30252 54628 30258
rect 54576 30194 54628 30200
rect 53656 30184 53708 30190
rect 53656 30126 53708 30132
rect 53564 29368 53616 29374
rect 53564 29310 53616 29316
rect 52368 28552 52420 28558
rect 52368 28494 52420 28500
rect 51448 28348 51500 28354
rect 51448 28290 51500 28296
rect 51724 27668 51776 27674
rect 51724 27610 51776 27616
rect 51736 3602 51764 27610
rect 51724 3596 51776 3602
rect 51724 3538 51776 3544
rect 52380 3534 52408 28494
rect 53668 3534 53696 30126
rect 53748 29368 53800 29374
rect 53748 29310 53800 29316
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 53656 3528 53708 3534
rect 53656 3470 53708 3476
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 49608 3460 49660 3466
rect 49608 3402 49660 3408
rect 48976 480 49004 3402
rect 50172 480 50200 3470
rect 51368 480 51396 3470
rect 52564 480 52592 3470
rect 53760 480 53788 29310
rect 55128 28348 55180 28354
rect 55128 28290 55180 28296
rect 55140 6914 55168 28290
rect 55692 27674 55720 32028
rect 56508 30252 56560 30258
rect 56508 30194 56560 30200
rect 55680 27668 55732 27674
rect 55680 27610 55732 27616
rect 54956 6886 55168 6914
rect 54956 480 54984 6886
rect 56520 3534 56548 30194
rect 56704 29238 56732 32028
rect 57808 29510 57836 32028
rect 57796 29504 57848 29510
rect 57796 29446 57848 29452
rect 57888 29504 57940 29510
rect 57888 29446 57940 29452
rect 56692 29232 56744 29238
rect 56692 29174 56744 29180
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56508 3528 56560 3534
rect 56508 3470 56560 3476
rect 56060 480 56088 3470
rect 57900 3466 57928 29446
rect 58820 28490 58848 32028
rect 59924 29102 59952 32028
rect 60936 29442 60964 32028
rect 60924 29436 60976 29442
rect 60924 29378 60976 29384
rect 61936 29300 61988 29306
rect 61936 29242 61988 29248
rect 60648 29232 60700 29238
rect 60648 29174 60700 29180
rect 59912 29096 59964 29102
rect 59912 29038 59964 29044
rect 58808 28484 58860 28490
rect 58808 28426 58860 28432
rect 59268 28484 59320 28490
rect 59268 28426 59320 28432
rect 59280 3534 59308 28426
rect 60660 3534 60688 29174
rect 60832 26784 60884 26790
rect 60832 26726 60884 26732
rect 60844 4962 60872 26726
rect 61948 26234 61976 29242
rect 62040 26790 62068 32028
rect 63052 30054 63080 32028
rect 63040 30048 63092 30054
rect 63040 29990 63092 29996
rect 63408 30048 63460 30054
rect 63408 29990 63460 29996
rect 62028 26784 62080 26790
rect 62028 26726 62080 26732
rect 61948 26206 62068 26234
rect 60832 4956 60884 4962
rect 60832 4898 60884 4904
rect 62040 3534 62068 26206
rect 63420 6914 63448 29990
rect 64064 29034 64092 32028
rect 64788 29436 64840 29442
rect 64788 29378 64840 29384
rect 64052 29028 64104 29034
rect 64052 28970 64104 28976
rect 63236 6886 63448 6914
rect 62212 5296 62264 5302
rect 62212 5238 62264 5244
rect 62120 4820 62172 4826
rect 62120 4762 62172 4768
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 60832 3528 60884 3534
rect 60832 3470 60884 3476
rect 62028 3528 62080 3534
rect 62028 3470 62080 3476
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 57888 3460 57940 3466
rect 57888 3402 57940 3408
rect 57256 480 57284 3402
rect 58452 480 58480 3470
rect 59648 480 59676 3470
rect 60844 480 60872 3470
rect 62132 2802 62160 4762
rect 62224 3602 62252 5238
rect 62212 3596 62264 3602
rect 62212 3538 62264 3544
rect 62040 2774 62160 2802
rect 62040 480 62068 2774
rect 63236 480 63264 6886
rect 64800 3534 64828 29378
rect 65168 5302 65196 32028
rect 66180 30122 66208 32028
rect 66168 30116 66220 30122
rect 66168 30058 66220 30064
rect 67284 29782 67312 32028
rect 67548 30116 67600 30122
rect 67548 30058 67600 30064
rect 67272 29776 67324 29782
rect 67272 29718 67324 29724
rect 66168 28620 66220 28626
rect 66168 28562 66220 28568
rect 65156 5296 65208 5302
rect 65156 5238 65208 5244
rect 66180 3534 66208 28562
rect 67560 3534 67588 30058
rect 68296 28286 68324 32028
rect 69400 29850 69428 32028
rect 69388 29844 69440 29850
rect 69388 29786 69440 29792
rect 70308 29844 70360 29850
rect 70308 29786 70360 29792
rect 68928 29776 68980 29782
rect 68928 29718 68980 29724
rect 68284 28280 68336 28286
rect 68284 28222 68336 28228
rect 68940 3534 68968 29718
rect 69112 6180 69164 6186
rect 69112 6122 69164 6128
rect 64328 3528 64380 3534
rect 64328 3470 64380 3476
rect 64788 3528 64840 3534
rect 64788 3470 64840 3476
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 66720 3528 66772 3534
rect 66720 3470 66772 3476
rect 67548 3528 67600 3534
rect 67548 3470 67600 3476
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 64340 480 64368 3470
rect 65536 480 65564 3470
rect 66732 480 66760 3470
rect 67928 480 67956 3470
rect 69124 480 69152 6122
rect 70320 480 70348 29786
rect 70412 29646 70440 32028
rect 71516 29986 71544 32028
rect 71504 29980 71556 29986
rect 71504 29922 71556 29928
rect 72528 29918 72556 32028
rect 72516 29912 72568 29918
rect 72516 29854 72568 29860
rect 73632 29714 73660 32028
rect 73620 29708 73672 29714
rect 73620 29650 73672 29656
rect 70400 29640 70452 29646
rect 70400 29582 70452 29588
rect 71688 29640 71740 29646
rect 71688 29582 71740 29588
rect 71700 6914 71728 29582
rect 74448 29164 74500 29170
rect 74448 29106 74500 29112
rect 73068 28280 73120 28286
rect 73068 28222 73120 28228
rect 71516 6886 71728 6914
rect 71516 480 71544 6886
rect 73080 3534 73108 28222
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 72620 480 72648 3470
rect 74460 2990 74488 29106
rect 74644 28422 74672 32028
rect 75748 29578 75776 32028
rect 76760 30326 76788 32028
rect 76748 30320 76800 30326
rect 76748 30262 76800 30268
rect 75828 29912 75880 29918
rect 75828 29854 75880 29860
rect 75736 29572 75788 29578
rect 75736 29514 75788 29520
rect 74632 28416 74684 28422
rect 74632 28358 74684 28364
rect 75840 3534 75868 29854
rect 77772 28558 77800 32028
rect 78588 30320 78640 30326
rect 78588 30262 78640 30268
rect 78496 29708 78548 29714
rect 78496 29650 78548 29656
rect 77760 28552 77812 28558
rect 77760 28494 77812 28500
rect 77208 28416 77260 28422
rect 77208 28358 77260 28364
rect 77220 3534 77248 28358
rect 78508 16574 78536 29650
rect 78416 16546 78536 16574
rect 77392 3596 77444 3602
rect 77392 3538 77444 3544
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 73804 2984 73856 2990
rect 73804 2926 73856 2932
rect 74448 2984 74500 2990
rect 74448 2926 74500 2932
rect 73816 480 73844 2926
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77404 480 77432 3538
rect 78416 3482 78444 16546
rect 78600 6914 78628 30262
rect 78876 30190 78904 32028
rect 78864 30184 78916 30190
rect 78864 30126 78916 30132
rect 79888 29374 79916 32028
rect 79876 29368 79928 29374
rect 79876 29310 79928 29316
rect 79968 28552 80020 28558
rect 79968 28494 80020 28500
rect 79980 6914 80008 28494
rect 80992 28354 81020 32028
rect 82004 30258 82032 32028
rect 81992 30252 82044 30258
rect 81992 30194 82044 30200
rect 82728 29980 82780 29986
rect 82728 29922 82780 29928
rect 81348 29572 81400 29578
rect 81348 29514 81400 29520
rect 80980 28348 81032 28354
rect 80980 28290 81032 28296
rect 78508 6886 78628 6914
rect 79704 6886 80008 6914
rect 78508 3602 78536 6886
rect 78496 3596 78548 3602
rect 78496 3538 78548 3544
rect 78416 3454 78628 3482
rect 78600 480 78628 3454
rect 79704 480 79732 6886
rect 81360 3330 81388 29514
rect 82740 3534 82768 29922
rect 83108 29510 83136 32028
rect 83096 29504 83148 29510
rect 83096 29446 83148 29452
rect 84120 28490 84148 32028
rect 85224 29238 85252 32028
rect 85488 29368 85540 29374
rect 85488 29310 85540 29316
rect 85212 29232 85264 29238
rect 85212 29174 85264 29180
rect 84108 28484 84160 28490
rect 84108 28426 84160 28432
rect 84108 28348 84160 28354
rect 84108 28290 84160 28296
rect 84120 3534 84148 28290
rect 85500 3534 85528 29310
rect 86236 29306 86264 32028
rect 86868 30252 86920 30258
rect 86868 30194 86920 30200
rect 86776 29504 86828 29510
rect 86776 29446 86828 29452
rect 86224 29300 86276 29306
rect 86224 29242 86276 29248
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 82728 3528 82780 3534
rect 82728 3470 82780 3476
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 84108 3528 84160 3534
rect 84108 3470 84160 3476
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 80888 3324 80940 3330
rect 80888 3266 80940 3272
rect 81348 3324 81400 3330
rect 81348 3266 81400 3272
rect 80900 480 80928 3266
rect 82096 480 82124 3470
rect 83292 480 83320 3470
rect 84488 480 84516 3470
rect 86788 3330 86816 29446
rect 85672 3324 85724 3330
rect 85672 3266 85724 3272
rect 86776 3324 86828 3330
rect 86776 3266 86828 3272
rect 85684 480 85712 3266
rect 86880 480 86908 30194
rect 87340 4826 87368 32028
rect 88248 30184 88300 30190
rect 88248 30126 88300 30132
rect 88260 6914 88288 30126
rect 88352 30054 88380 32028
rect 88340 30048 88392 30054
rect 88340 29990 88392 29996
rect 89456 29442 89484 32028
rect 89628 30048 89680 30054
rect 89628 29990 89680 29996
rect 89444 29436 89496 29442
rect 89444 29378 89496 29384
rect 87984 6886 88288 6914
rect 87328 4820 87380 4826
rect 87328 4762 87380 4768
rect 87984 480 88012 6886
rect 89640 3330 89668 29990
rect 90468 28626 90496 32028
rect 91572 30122 91600 32028
rect 91560 30116 91612 30122
rect 91560 30058 91612 30064
rect 92388 30116 92440 30122
rect 92388 30058 92440 30064
rect 91008 29436 91060 29442
rect 91008 29378 91060 29384
rect 90456 28620 90508 28626
rect 90456 28562 90508 28568
rect 91020 3534 91048 29378
rect 92400 3534 92428 30058
rect 92584 29782 92612 32028
rect 92572 29776 92624 29782
rect 92572 29718 92624 29724
rect 93596 6186 93624 32028
rect 94700 29850 94728 32028
rect 94688 29844 94740 29850
rect 94688 29786 94740 29792
rect 93768 29776 93820 29782
rect 93768 29718 93820 29724
rect 93584 6180 93636 6186
rect 93584 6122 93636 6128
rect 93780 3534 93808 29718
rect 95712 29646 95740 32028
rect 96528 29844 96580 29850
rect 96528 29786 96580 29792
rect 95700 29640 95752 29646
rect 95700 29582 95752 29588
rect 95148 29300 95200 29306
rect 95148 29242 95200 29248
rect 95056 29096 95108 29102
rect 95056 29038 95108 29044
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 92388 3528 92440 3534
rect 92388 3470 92440 3476
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 89168 3324 89220 3330
rect 89168 3266 89220 3272
rect 89628 3324 89680 3330
rect 89628 3266 89680 3272
rect 89180 480 89208 3266
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 92768 480 92796 3470
rect 95068 3330 95096 29038
rect 93952 3324 94004 3330
rect 93952 3266 94004 3272
rect 95056 3324 95108 3330
rect 95056 3266 95108 3272
rect 93964 480 93992 3266
rect 95160 480 95188 29242
rect 96540 6914 96568 29786
rect 96816 28286 96844 32028
rect 97828 29170 97856 32028
rect 98932 29918 98960 32028
rect 98920 29912 98972 29918
rect 98920 29854 98972 29860
rect 97908 29232 97960 29238
rect 97908 29174 97960 29180
rect 97816 29164 97868 29170
rect 97816 29106 97868 29112
rect 96804 28280 96856 28286
rect 96804 28222 96856 28228
rect 96264 6886 96568 6914
rect 96264 480 96292 6886
rect 97920 3330 97948 29174
rect 99288 29028 99340 29034
rect 99288 28970 99340 28976
rect 99300 3534 99328 28970
rect 99944 28422 99972 32028
rect 101048 30326 101076 32028
rect 101036 30320 101088 30326
rect 101036 30262 101088 30268
rect 101956 30320 102008 30326
rect 101956 30262 102008 30268
rect 100668 29912 100720 29918
rect 100668 29854 100720 29860
rect 99932 28416 99984 28422
rect 99932 28358 99984 28364
rect 100680 3534 100708 29854
rect 100760 29640 100812 29646
rect 100760 29582 100812 29588
rect 100772 28558 100800 29582
rect 100760 28552 100812 28558
rect 100760 28494 100812 28500
rect 101968 26234 101996 30262
rect 102060 29714 102088 32028
rect 102048 29708 102100 29714
rect 102048 29650 102100 29656
rect 103164 29646 103192 32028
rect 103152 29640 103204 29646
rect 103152 29582 103204 29588
rect 103336 29640 103388 29646
rect 103336 29582 103388 29588
rect 101968 26206 102088 26234
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 97448 3324 97500 3330
rect 97448 3266 97500 3272
rect 97908 3324 97960 3330
rect 97908 3266 97960 3272
rect 97460 480 97488 3266
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 102060 3262 102088 26206
rect 102232 3460 102284 3466
rect 102232 3402 102284 3408
rect 101036 3256 101088 3262
rect 101036 3198 101088 3204
rect 102048 3256 102100 3262
rect 102048 3198 102100 3204
rect 101048 480 101076 3198
rect 102244 480 102272 3402
rect 103348 480 103376 29582
rect 104176 29578 104204 32028
rect 105280 29986 105308 32028
rect 105268 29980 105320 29986
rect 105268 29922 105320 29928
rect 104164 29572 104216 29578
rect 104164 29514 104216 29520
rect 104808 29572 104860 29578
rect 104808 29514 104860 29520
rect 103428 29164 103480 29170
rect 103428 29106 103480 29112
rect 103440 3466 103468 29106
rect 104820 6914 104848 29514
rect 106188 29368 106240 29374
rect 106188 29310 106240 29316
rect 104544 6886 104848 6914
rect 103428 3460 103480 3466
rect 103428 3402 103480 3408
rect 104544 480 104572 6886
rect 106200 3534 106228 29310
rect 106292 28354 106320 32028
rect 107304 29442 107332 32028
rect 107568 29708 107620 29714
rect 107568 29650 107620 29656
rect 107292 29436 107344 29442
rect 107292 29378 107344 29384
rect 106280 28348 106332 28354
rect 106280 28290 106332 28296
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 105740 480 105768 3470
rect 107580 3466 107608 29650
rect 108408 29510 108436 32028
rect 109420 30258 109448 32028
rect 109408 30252 109460 30258
rect 109408 30194 109460 30200
rect 110524 30190 110552 32028
rect 110512 30184 110564 30190
rect 110512 30126 110564 30132
rect 111536 30054 111564 32028
rect 111616 30252 111668 30258
rect 111616 30194 111668 30200
rect 111524 30048 111576 30054
rect 111524 29990 111576 29996
rect 108948 29980 109000 29986
rect 108948 29922 109000 29928
rect 108396 29504 108448 29510
rect 108396 29446 108448 29452
rect 108960 3534 108988 29922
rect 110328 29436 110380 29442
rect 110328 29378 110380 29384
rect 110340 3534 110368 29378
rect 111628 16574 111656 30194
rect 111708 30048 111760 30054
rect 111708 29990 111760 29996
rect 111536 16546 111656 16574
rect 111536 3534 111564 16546
rect 111720 6914 111748 29990
rect 112640 29510 112668 32028
rect 113088 30184 113140 30190
rect 113088 30126 113140 30132
rect 112628 29504 112680 29510
rect 112628 29446 112680 29452
rect 113100 6914 113128 30126
rect 113652 30122 113680 32028
rect 113640 30116 113692 30122
rect 113640 30058 113692 30064
rect 114756 29782 114784 32028
rect 114744 29776 114796 29782
rect 114744 29718 114796 29724
rect 114468 29504 114520 29510
rect 114468 29446 114520 29452
rect 111628 6886 111748 6914
rect 112824 6886 113128 6914
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 110328 3528 110380 3534
rect 110328 3470 110380 3476
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 111524 3528 111576 3534
rect 111524 3470 111576 3476
rect 106924 3460 106976 3466
rect 106924 3402 106976 3408
rect 107568 3460 107620 3466
rect 107568 3402 107620 3408
rect 106936 480 106964 3402
rect 108132 480 108160 3470
rect 109328 480 109356 3470
rect 110524 480 110552 3470
rect 111628 480 111656 6886
rect 112824 480 112852 6886
rect 114480 3534 114508 29446
rect 115768 29102 115796 32028
rect 116872 29306 116900 32028
rect 117884 29850 117912 32028
rect 117872 29844 117924 29850
rect 117872 29786 117924 29792
rect 118608 29844 118660 29850
rect 118608 29786 118660 29792
rect 116860 29300 116912 29306
rect 116860 29242 116912 29248
rect 117228 29232 117280 29238
rect 117228 29174 117280 29180
rect 115756 29096 115808 29102
rect 115756 29038 115808 29044
rect 115848 29096 115900 29102
rect 115848 29038 115900 29044
rect 115860 3534 115888 29038
rect 117240 3534 117268 29174
rect 118620 3534 118648 29786
rect 118988 29306 119016 32028
rect 120000 29866 120028 32028
rect 121104 29918 121132 32028
rect 122116 30326 122144 32028
rect 122104 30320 122156 30326
rect 122104 30262 122156 30268
rect 119724 29838 120028 29866
rect 121092 29912 121144 29918
rect 121092 29854 121144 29860
rect 122748 29912 122800 29918
rect 122748 29854 122800 29860
rect 118976 29300 119028 29306
rect 118976 29242 119028 29248
rect 119724 29034 119752 29838
rect 119896 29776 119948 29782
rect 119896 29718 119948 29724
rect 119712 29028 119764 29034
rect 119712 28970 119764 28976
rect 119804 29028 119856 29034
rect 119804 28970 119856 28976
rect 114008 3528 114060 3534
rect 114008 3470 114060 3476
rect 114468 3528 114520 3534
rect 114468 3470 114520 3476
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 117228 3528 117280 3534
rect 117228 3470 117280 3476
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 118608 3528 118660 3534
rect 118608 3470 118660 3476
rect 114020 480 114048 3470
rect 115216 480 115244 3470
rect 116412 480 116440 3470
rect 117608 480 117636 3470
rect 119816 3126 119844 28970
rect 118792 3120 118844 3126
rect 118792 3062 118844 3068
rect 119804 3120 119856 3126
rect 119804 3062 119856 3068
rect 118804 480 118832 3062
rect 119908 480 119936 29718
rect 121368 29300 121420 29306
rect 121368 29242 121420 29248
rect 121380 6914 121408 29242
rect 121104 6886 121408 6914
rect 121104 480 121132 6886
rect 122760 3534 122788 29854
rect 123128 29170 123156 32028
rect 124128 30116 124180 30122
rect 124128 30058 124180 30064
rect 123116 29164 123168 29170
rect 123116 29106 123168 29112
rect 124140 3534 124168 30058
rect 124232 29646 124260 32028
rect 124220 29640 124272 29646
rect 124220 29582 124272 29588
rect 125244 29578 125272 32028
rect 125232 29572 125284 29578
rect 125232 29514 125284 29520
rect 125508 29572 125560 29578
rect 125508 29514 125560 29520
rect 125520 3534 125548 29514
rect 126348 29374 126376 32028
rect 127360 29714 127388 32028
rect 128268 30320 128320 30326
rect 128268 30262 128320 30268
rect 127348 29708 127400 29714
rect 127348 29650 127400 29656
rect 128176 29640 128228 29646
rect 128176 29582 128228 29588
rect 126336 29368 126388 29374
rect 126336 29310 126388 29316
rect 126888 29368 126940 29374
rect 126888 29310 126940 29316
rect 126900 3534 126928 29310
rect 122288 3528 122340 3534
rect 122288 3470 122340 3476
rect 122748 3528 122800 3534
rect 122748 3470 122800 3476
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 122300 480 122328 3470
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 126992 480 127020 3470
rect 128188 480 128216 29582
rect 128280 3534 128308 30262
rect 128464 29986 128492 32028
rect 128452 29980 128504 29986
rect 128452 29922 128504 29928
rect 129476 29442 129504 32028
rect 130580 30258 130608 32028
rect 130568 30252 130620 30258
rect 130568 30194 130620 30200
rect 131592 30054 131620 32028
rect 132696 30190 132724 32028
rect 132684 30184 132736 30190
rect 132684 30126 132736 30132
rect 131580 30048 131632 30054
rect 131580 29990 131632 29996
rect 132408 30048 132460 30054
rect 132408 29990 132460 29996
rect 131028 29980 131080 29986
rect 131028 29922 131080 29928
rect 129464 29436 129516 29442
rect 129464 29378 129516 29384
rect 129648 29436 129700 29442
rect 129648 29378 129700 29384
rect 129660 6914 129688 29378
rect 129384 6886 129688 6914
rect 128268 3528 128320 3534
rect 128268 3470 128320 3476
rect 129384 480 129412 6886
rect 131040 3534 131068 29922
rect 130568 3528 130620 3534
rect 130568 3470 130620 3476
rect 131028 3528 131080 3534
rect 131028 3470 131080 3476
rect 130580 480 130608 3470
rect 132420 3466 132448 29990
rect 133708 29510 133736 32028
rect 133788 30184 133840 30190
rect 133788 30126 133840 30132
rect 133696 29504 133748 29510
rect 133696 29446 133748 29452
rect 133800 3534 133828 30126
rect 134812 29102 134840 32028
rect 135824 29238 135852 32028
rect 136836 29850 136864 32028
rect 137940 30002 137968 32028
rect 137848 29974 137968 30002
rect 136824 29844 136876 29850
rect 136824 29786 136876 29792
rect 136456 29708 136508 29714
rect 136456 29650 136508 29656
rect 135812 29232 135864 29238
rect 135812 29174 135864 29180
rect 135168 29164 135220 29170
rect 135168 29106 135220 29112
rect 134800 29096 134852 29102
rect 134800 29038 134852 29044
rect 135180 3534 135208 29106
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 134156 3528 134208 3534
rect 134156 3470 134208 3476
rect 135168 3528 135220 3534
rect 135168 3470 135220 3476
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 132408 3460 132460 3466
rect 132408 3402 132460 3408
rect 131776 480 131804 3402
rect 132972 480 133000 3470
rect 134168 480 134196 3470
rect 135260 2916 135312 2922
rect 135260 2858 135312 2864
rect 135272 480 135300 2858
rect 136468 480 136496 29650
rect 136548 29232 136600 29238
rect 136548 29174 136600 29180
rect 136560 2922 136588 29174
rect 137848 29034 137876 29974
rect 137928 29844 137980 29850
rect 137928 29786 137980 29792
rect 137836 29028 137888 29034
rect 137836 28970 137888 28976
rect 137940 6914 137968 29786
rect 138952 29782 138980 32028
rect 138940 29776 138992 29782
rect 138940 29718 138992 29724
rect 140056 29306 140084 32028
rect 141068 29918 141096 32028
rect 142172 30122 142200 32028
rect 142160 30116 142212 30122
rect 142160 30058 142212 30064
rect 141056 29912 141108 29918
rect 141056 29854 141108 29860
rect 143184 29578 143212 32028
rect 143448 29912 143500 29918
rect 143448 29854 143500 29860
rect 143172 29572 143224 29578
rect 143172 29514 143224 29520
rect 140688 29504 140740 29510
rect 140688 29446 140740 29452
rect 140044 29300 140096 29306
rect 140044 29242 140096 29248
rect 139308 29096 139360 29102
rect 139308 29038 139360 29044
rect 137664 6886 137968 6914
rect 136548 2916 136600 2922
rect 136548 2858 136600 2864
rect 137664 480 137692 6886
rect 139320 3534 139348 29038
rect 140700 3534 140728 29446
rect 142068 29300 142120 29306
rect 142068 29242 142120 29248
rect 142080 3534 142108 29242
rect 143460 3534 143488 29854
rect 144288 29374 144316 32028
rect 145300 30326 145328 32028
rect 145288 30320 145340 30326
rect 145288 30262 145340 30268
rect 146208 30320 146260 30326
rect 146208 30262 146260 30268
rect 144736 29776 144788 29782
rect 144736 29718 144788 29724
rect 144276 29368 144328 29374
rect 144276 29310 144328 29316
rect 138848 3528 138900 3534
rect 138848 3470 138900 3476
rect 139308 3528 139360 3534
rect 139308 3470 139360 3476
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 140688 3528 140740 3534
rect 140688 3470 140740 3476
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 142068 3528 142120 3534
rect 142068 3470 142120 3476
rect 142436 3528 142488 3534
rect 142436 3470 142488 3476
rect 143448 3528 143500 3534
rect 143448 3470 143500 3476
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 138860 480 138888 3470
rect 140056 480 140084 3470
rect 141252 480 141280 3470
rect 142448 480 142476 3470
rect 143552 480 143580 3470
rect 144748 480 144776 29718
rect 144828 29572 144880 29578
rect 144828 29514 144880 29520
rect 144840 3534 144868 29514
rect 146220 6914 146248 30262
rect 146404 29646 146432 32028
rect 146392 29640 146444 29646
rect 146392 29582 146444 29588
rect 147416 29442 147444 32028
rect 147588 30116 147640 30122
rect 147588 30058 147640 30064
rect 147404 29436 147456 29442
rect 147404 29378 147456 29384
rect 145944 6886 146248 6914
rect 144828 3528 144880 3534
rect 144828 3470 144880 3476
rect 145944 480 145972 6886
rect 147600 3534 147628 30058
rect 148520 29986 148548 32028
rect 149532 30054 149560 32028
rect 150636 30190 150664 32028
rect 150624 30184 150676 30190
rect 150624 30126 150676 30132
rect 149520 30048 149572 30054
rect 149520 29990 149572 29996
rect 148508 29980 148560 29986
rect 148508 29922 148560 29928
rect 148968 29980 149020 29986
rect 148968 29922 149020 29928
rect 148980 3534 149008 29922
rect 150348 29368 150400 29374
rect 150348 29310 150400 29316
rect 150360 3534 150388 29310
rect 151648 29170 151676 32028
rect 152660 29238 152688 32028
rect 153764 29714 153792 32028
rect 154488 30048 154540 30054
rect 154488 29990 154540 29996
rect 153752 29708 153804 29714
rect 153752 29650 153804 29656
rect 153016 29640 153068 29646
rect 153016 29582 153068 29588
rect 152648 29232 152700 29238
rect 152648 29174 152700 29180
rect 151636 29164 151688 29170
rect 151636 29106 151688 29112
rect 151728 29164 151780 29170
rect 151728 29106 151780 29112
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 150348 3528 150400 3534
rect 150348 3470 150400 3476
rect 147140 480 147168 3470
rect 148336 480 148364 3470
rect 149532 480 149560 3470
rect 151740 3058 151768 29106
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 150624 3052 150676 3058
rect 150624 2994 150676 3000
rect 151728 3052 151780 3058
rect 151728 2994 151780 3000
rect 150636 480 150664 2994
rect 151832 480 151860 3470
rect 153028 480 153056 29582
rect 153108 29436 153160 29442
rect 153108 29378 153160 29384
rect 153120 3534 153148 29378
rect 154500 6914 154528 29990
rect 154776 29850 154804 32028
rect 155776 30252 155828 30258
rect 155776 30194 155828 30200
rect 154764 29844 154816 29850
rect 154764 29786 154816 29792
rect 154224 6886 154528 6914
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 154224 480 154252 6886
rect 155420 598 155632 626
rect 155420 480 155448 598
rect 155604 490 155632 598
rect 155788 490 155816 30194
rect 155880 29102 155908 32028
rect 156892 29510 156920 32028
rect 157248 29844 157300 29850
rect 157248 29786 157300 29792
rect 156880 29504 156932 29510
rect 156880 29446 156932 29452
rect 155868 29096 155920 29102
rect 155868 29038 155920 29044
rect 157260 3534 157288 29786
rect 157996 29306 158024 32028
rect 158628 30184 158680 30190
rect 158628 30126 158680 30132
rect 157984 29300 158036 29306
rect 157984 29242 158036 29248
rect 158640 3534 158668 30126
rect 159008 29918 159036 32028
rect 158996 29912 159048 29918
rect 158996 29854 159048 29860
rect 160112 29578 160140 32028
rect 161124 29782 161152 32028
rect 162228 30326 162256 32028
rect 162216 30320 162268 30326
rect 162216 30262 162268 30268
rect 163240 30122 163268 32028
rect 163228 30116 163280 30122
rect 163228 30058 163280 30064
rect 164344 29986 164372 32028
rect 164332 29980 164384 29986
rect 164332 29922 164384 29928
rect 164148 29912 164200 29918
rect 164148 29854 164200 29860
rect 161112 29776 161164 29782
rect 161112 29718 161164 29724
rect 162768 29776 162820 29782
rect 162768 29718 162820 29724
rect 161296 29708 161348 29714
rect 161296 29650 161348 29656
rect 160100 29572 160152 29578
rect 160100 29514 160152 29520
rect 160008 29504 160060 29510
rect 160008 29446 160060 29452
rect 160020 3534 160048 29446
rect 156604 3528 156656 3534
rect 156604 3470 156656 3476
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 157800 3528 157852 3534
rect 157800 3470 157852 3476
rect 158628 3528 158680 3534
rect 158628 3470 158680 3476
rect 158904 3528 158956 3534
rect 158904 3470 158956 3476
rect 160008 3528 160060 3534
rect 160008 3470 160060 3476
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 155604 462 155816 490
rect 156616 480 156644 3470
rect 157812 480 157840 3470
rect 158916 480 158944 3470
rect 160112 480 160140 3470
rect 161308 480 161336 29650
rect 161388 29300 161440 29306
rect 161388 29242 161440 29248
rect 161400 3534 161428 29242
rect 162780 6914 162808 29718
rect 162504 6886 162808 6914
rect 161388 3528 161440 3534
rect 161388 3470 161440 3476
rect 162504 480 162532 6886
rect 164160 3534 164188 29854
rect 165356 29374 165384 32028
rect 165528 29572 165580 29578
rect 165528 29514 165580 29520
rect 165344 29368 165396 29374
rect 165344 29310 165396 29316
rect 165540 3534 165568 29514
rect 166368 29170 166396 32028
rect 166908 30116 166960 30122
rect 166908 30058 166960 30064
rect 166356 29164 166408 29170
rect 166356 29106 166408 29112
rect 166920 3534 166948 30058
rect 167472 29442 167500 32028
rect 168288 30320 168340 30326
rect 168288 30262 168340 30268
rect 167460 29436 167512 29442
rect 167460 29378 167512 29384
rect 168300 3534 168328 30262
rect 168484 29646 168512 32028
rect 169588 30054 169616 32028
rect 170600 30258 170628 32028
rect 170588 30252 170640 30258
rect 170588 30194 170640 30200
rect 169576 30048 169628 30054
rect 169576 29990 169628 29996
rect 171048 29980 171100 29986
rect 171048 29922 171100 29928
rect 168472 29640 168524 29646
rect 168472 29582 168524 29588
rect 169576 29640 169628 29646
rect 169576 29582 169628 29588
rect 169588 16574 169616 29582
rect 169668 29436 169720 29442
rect 169668 29378 169720 29384
rect 169496 16546 169616 16574
rect 163688 3528 163740 3534
rect 163688 3470 163740 3476
rect 164148 3528 164200 3534
rect 164148 3470 164200 3476
rect 164884 3528 164936 3534
rect 164884 3470 164936 3476
rect 165528 3528 165580 3534
rect 165528 3470 165580 3476
rect 166080 3528 166132 3534
rect 166080 3470 166132 3476
rect 166908 3528 166960 3534
rect 166908 3470 166960 3476
rect 167184 3528 167236 3534
rect 167184 3470 167236 3476
rect 168288 3528 168340 3534
rect 168288 3470 168340 3476
rect 163700 480 163728 3470
rect 164896 480 164924 3470
rect 166092 480 166120 3470
rect 167196 480 167224 3470
rect 169496 3058 169524 16546
rect 169680 6914 169708 29378
rect 171060 6914 171088 29922
rect 171704 29850 171732 32028
rect 172716 30190 172744 32028
rect 172704 30184 172756 30190
rect 172704 30126 172756 30132
rect 173716 30048 173768 30054
rect 173716 29990 173768 29996
rect 171692 29844 171744 29850
rect 171692 29786 171744 29792
rect 172428 29844 172480 29850
rect 172428 29786 172480 29792
rect 169588 6886 169708 6914
rect 170784 6886 171088 6914
rect 168380 3052 168432 3058
rect 168380 2994 168432 3000
rect 169484 3052 169536 3058
rect 169484 2994 169536 3000
rect 168392 480 168420 2994
rect 169588 480 169616 6886
rect 170784 480 170812 6886
rect 172440 3534 172468 29786
rect 173728 26234 173756 29990
rect 173820 29510 173848 32028
rect 173808 29504 173860 29510
rect 173808 29446 173860 29452
rect 174832 29306 174860 32028
rect 175188 30184 175240 30190
rect 175188 30126 175240 30132
rect 174820 29300 174872 29306
rect 174820 29242 174872 29248
rect 173728 26206 173848 26234
rect 173820 3534 173848 26206
rect 175200 3534 175228 30126
rect 175936 29714 175964 32028
rect 176948 29782 176976 32028
rect 178052 29918 178080 32028
rect 178040 29912 178092 29918
rect 178040 29854 178092 29860
rect 176936 29776 176988 29782
rect 176936 29718 176988 29724
rect 177856 29776 177908 29782
rect 177856 29718 177908 29724
rect 175924 29708 175976 29714
rect 175924 29650 175976 29656
rect 176568 29504 176620 29510
rect 176568 29446 176620 29452
rect 176580 3534 176608 29446
rect 177868 16574 177896 29718
rect 177948 29708 178000 29714
rect 177948 29650 178000 29656
rect 177776 16546 177896 16574
rect 177776 3534 177804 16546
rect 177960 6914 177988 29650
rect 179064 29578 179092 32028
rect 179328 30252 179380 30258
rect 179328 30194 179380 30200
rect 179052 29572 179104 29578
rect 179052 29514 179104 29520
rect 179340 6914 179368 30194
rect 180168 30122 180196 32028
rect 181180 30326 181208 32028
rect 181168 30320 181220 30326
rect 181168 30262 181220 30268
rect 180156 30116 180208 30122
rect 180156 30058 180208 30064
rect 182088 30116 182140 30122
rect 182088 30058 182140 30064
rect 180708 29912 180760 29918
rect 180708 29854 180760 29860
rect 177868 6886 177988 6914
rect 179064 6886 179368 6914
rect 171968 3528 172020 3534
rect 171968 3470 172020 3476
rect 172428 3528 172480 3534
rect 172428 3470 172480 3476
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 175188 3528 175240 3534
rect 175188 3470 175240 3476
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 176568 3528 176620 3534
rect 176568 3470 176620 3476
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 177764 3528 177816 3534
rect 177764 3470 177816 3476
rect 171980 480 172008 3470
rect 173176 480 173204 3470
rect 174280 480 174308 3470
rect 175476 480 175504 3470
rect 176672 480 176700 3470
rect 177868 480 177896 6886
rect 179064 480 179092 6886
rect 180720 3534 180748 29854
rect 182100 3534 182128 30058
rect 182192 29646 182220 32028
rect 182180 29640 182232 29646
rect 182180 29582 182232 29588
rect 183296 29442 183324 32028
rect 183468 30320 183520 30326
rect 183468 30262 183520 30268
rect 183284 29436 183336 29442
rect 183284 29378 183336 29384
rect 183480 3534 183508 30262
rect 184308 29986 184336 32028
rect 184296 29980 184348 29986
rect 184296 29922 184348 29928
rect 185412 29850 185440 32028
rect 186424 30054 186452 32028
rect 187528 30190 187556 32028
rect 187516 30184 187568 30190
rect 187516 30126 187568 30132
rect 186412 30048 186464 30054
rect 186412 29990 186464 29996
rect 185400 29844 185452 29850
rect 185400 29786 185452 29792
rect 187608 29844 187660 29850
rect 187608 29786 187660 29792
rect 186136 29640 186188 29646
rect 186136 29582 186188 29588
rect 184848 29436 184900 29442
rect 184848 29378 184900 29384
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 181444 3528 181496 3534
rect 181444 3470 181496 3476
rect 182088 3528 182140 3534
rect 182088 3470 182140 3476
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 180260 480 180288 3470
rect 181456 480 181484 3470
rect 182560 480 182588 3470
rect 184860 3262 184888 29378
rect 184940 3528 184992 3534
rect 184940 3470 184992 3476
rect 183744 3256 183796 3262
rect 183744 3198 183796 3204
rect 184848 3256 184900 3262
rect 184848 3198 184900 3204
rect 183756 480 183784 3198
rect 184952 480 184980 3470
rect 186148 480 186176 29582
rect 186228 29572 186280 29578
rect 186228 29514 186280 29520
rect 186240 3534 186268 29514
rect 187620 6914 187648 29786
rect 188540 29510 188568 32028
rect 188988 29980 189040 29986
rect 188988 29922 189040 29928
rect 188528 29504 188580 29510
rect 188528 29446 188580 29452
rect 187344 6886 187648 6914
rect 186228 3528 186280 3534
rect 186228 3470 186280 3476
rect 187344 480 187372 6886
rect 189000 3534 189028 29922
rect 189644 29782 189672 32028
rect 190368 30184 190420 30190
rect 190368 30126 190420 30132
rect 189632 29776 189684 29782
rect 189632 29718 189684 29724
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 188988 3528 189040 3534
rect 188988 3470 189040 3476
rect 188540 480 188568 3470
rect 190380 3466 190408 30126
rect 190656 29714 190684 32028
rect 191760 30258 191788 32028
rect 191748 30252 191800 30258
rect 191748 30194 191800 30200
rect 192772 29918 192800 32028
rect 193128 30252 193180 30258
rect 193128 30194 193180 30200
rect 192760 29912 192812 29918
rect 192760 29854 192812 29860
rect 190644 29708 190696 29714
rect 190644 29650 190696 29656
rect 191748 29504 191800 29510
rect 191748 29446 191800 29452
rect 191760 3534 191788 29446
rect 193140 3534 193168 30194
rect 193876 30122 193904 32028
rect 194888 30326 194916 32028
rect 194876 30320 194928 30326
rect 195900 30274 195928 32028
rect 194876 30262 194928 30268
rect 195808 30246 195928 30274
rect 193864 30116 193916 30122
rect 193864 30058 193916 30064
rect 194508 29912 194560 29918
rect 194508 29854 194560 29860
rect 194416 29708 194468 29714
rect 194416 29650 194468 29656
rect 194428 16574 194456 29650
rect 194336 16546 194456 16574
rect 194336 3534 194364 16546
rect 194520 6914 194548 29854
rect 195808 29442 195836 30246
rect 195888 30116 195940 30122
rect 195888 30058 195940 30064
rect 195796 29436 195848 29442
rect 195796 29378 195848 29384
rect 195900 6914 195928 30058
rect 197004 29578 197032 32028
rect 197268 30048 197320 30054
rect 197268 29990 197320 29996
rect 196992 29572 197044 29578
rect 196992 29514 197044 29520
rect 194428 6886 194548 6914
rect 195624 6886 195928 6914
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 191748 3528 191800 3534
rect 191748 3470 191800 3476
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 193128 3528 193180 3534
rect 193128 3470 193180 3476
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 194324 3528 194376 3534
rect 194324 3470 194376 3476
rect 189724 3460 189776 3466
rect 189724 3402 189776 3408
rect 190368 3460 190420 3466
rect 190368 3402 190420 3408
rect 189736 480 189764 3402
rect 190840 480 190868 3470
rect 192036 480 192064 3470
rect 193232 480 193260 3470
rect 194428 480 194456 6886
rect 195624 480 195652 6886
rect 197280 3330 197308 29990
rect 198016 29646 198044 32028
rect 199120 29850 199148 32028
rect 200028 30320 200080 30326
rect 200028 30262 200080 30268
rect 199108 29844 199160 29850
rect 199108 29786 199160 29792
rect 198648 29776 198700 29782
rect 198648 29718 198700 29724
rect 198004 29640 198056 29646
rect 198004 29582 198056 29588
rect 198660 3534 198688 29718
rect 200040 3534 200068 30262
rect 200132 29986 200160 32028
rect 201236 30190 201264 32028
rect 201224 30184 201276 30190
rect 201224 30126 201276 30132
rect 200120 29980 200172 29986
rect 200120 29922 200172 29928
rect 201408 29844 201460 29850
rect 201408 29786 201460 29792
rect 197912 3528 197964 3534
rect 197912 3470 197964 3476
rect 198648 3528 198700 3534
rect 198648 3470 198700 3476
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 200028 3528 200080 3534
rect 200028 3470 200080 3476
rect 196808 3324 196860 3330
rect 196808 3266 196860 3272
rect 197268 3324 197320 3330
rect 197268 3266 197320 3272
rect 196820 480 196848 3266
rect 197924 480 197952 3470
rect 199120 480 199148 3470
rect 201420 3262 201448 29786
rect 202248 29510 202276 32028
rect 203352 30258 203380 32028
rect 203340 30252 203392 30258
rect 203340 30194 203392 30200
rect 202788 30184 202840 30190
rect 202788 30126 202840 30132
rect 202696 29640 202748 29646
rect 202696 29582 202748 29588
rect 202236 29504 202288 29510
rect 202236 29446 202288 29452
rect 201500 3528 201552 3534
rect 201500 3470 201552 3476
rect 200304 3256 200356 3262
rect 200304 3198 200356 3204
rect 201408 3256 201460 3262
rect 201408 3198 201460 3204
rect 200316 480 200344 3198
rect 201512 480 201540 3470
rect 202708 480 202736 29582
rect 202800 3534 202828 30126
rect 204168 29980 204220 29986
rect 204168 29922 204220 29928
rect 204180 6914 204208 29922
rect 204364 29714 204392 32028
rect 205468 29918 205496 32028
rect 205548 30252 205600 30258
rect 205548 30194 205600 30200
rect 205456 29912 205508 29918
rect 205456 29854 205508 29860
rect 204352 29708 204404 29714
rect 204352 29650 204404 29656
rect 203904 6886 204208 6914
rect 202788 3528 202840 3534
rect 202788 3470 202840 3476
rect 203904 480 203932 6886
rect 205560 3534 205588 30194
rect 206480 30122 206508 32028
rect 206468 30116 206520 30122
rect 206468 30058 206520 30064
rect 206928 30116 206980 30122
rect 206928 30058 206980 30064
rect 206940 3534 206968 30058
rect 207584 30054 207612 32028
rect 207572 30048 207624 30054
rect 207572 29990 207624 29996
rect 208596 29782 208624 32028
rect 209700 30326 209728 32028
rect 209688 30320 209740 30326
rect 209688 30262 209740 30268
rect 209688 29912 209740 29918
rect 209688 29854 209740 29860
rect 208584 29776 208636 29782
rect 208584 29718 208636 29724
rect 208308 29708 208360 29714
rect 208308 29650 208360 29656
rect 208320 3534 208348 29650
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 206192 3528 206244 3534
rect 206192 3470 206244 3476
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 207388 3528 207440 3534
rect 207388 3470 207440 3476
rect 208308 3528 208360 3534
rect 208308 3470 208360 3476
rect 205100 480 205128 3470
rect 206204 480 206232 3470
rect 207400 480 207428 3470
rect 209700 3058 209728 29854
rect 210712 29850 210740 32028
rect 211724 30190 211752 32028
rect 211712 30184 211764 30190
rect 211712 30126 211764 30132
rect 210700 29844 210752 29850
rect 210700 29786 210752 29792
rect 212448 29844 212500 29850
rect 212448 29786 212500 29792
rect 211068 29776 211120 29782
rect 211068 29718 211120 29724
rect 210976 29164 211028 29170
rect 210976 29106 211028 29112
rect 210988 16574 211016 29106
rect 210896 16546 211016 16574
rect 210896 3534 210924 16546
rect 211080 6914 211108 29718
rect 212460 6914 212488 29786
rect 212828 29646 212856 32028
rect 213840 29986 213868 32028
rect 214944 30258 214972 32028
rect 214932 30252 214984 30258
rect 214932 30194 214984 30200
rect 215956 30122 215984 32028
rect 216588 30184 216640 30190
rect 216588 30126 216640 30132
rect 215944 30116 215996 30122
rect 215944 30058 215996 30064
rect 213828 29980 213880 29986
rect 213828 29922 213880 29928
rect 215208 29980 215260 29986
rect 215208 29922 215260 29928
rect 212816 29640 212868 29646
rect 212816 29582 212868 29588
rect 213828 29640 213880 29646
rect 213828 29582 213880 29588
rect 210988 6886 211108 6914
rect 212184 6886 212488 6914
rect 209780 3528 209832 3534
rect 209780 3470 209832 3476
rect 210884 3528 210936 3534
rect 210884 3470 210936 3476
rect 208584 3052 208636 3058
rect 208584 2994 208636 3000
rect 209688 3052 209740 3058
rect 209688 2994 209740 3000
rect 208596 480 208624 2994
rect 209792 480 209820 3470
rect 210988 480 211016 6886
rect 212184 480 212212 6886
rect 213840 3534 213868 29582
rect 215220 3534 215248 29922
rect 216600 3534 216628 30126
rect 217060 29714 217088 32028
rect 217968 30116 218020 30122
rect 217968 30058 218020 30064
rect 217048 29708 217100 29714
rect 217048 29650 217100 29656
rect 217980 3534 218008 30058
rect 218072 29918 218100 32028
rect 218060 29912 218112 29918
rect 218060 29854 218112 29860
rect 219176 29170 219204 32028
rect 219348 29912 219400 29918
rect 219348 29854 219400 29860
rect 219256 29708 219308 29714
rect 219256 29650 219308 29656
rect 219164 29164 219216 29170
rect 219164 29106 219216 29112
rect 219268 16574 219296 29650
rect 219176 16546 219296 16574
rect 219176 3534 219204 16546
rect 219360 6914 219388 29854
rect 220188 29782 220216 32028
rect 221292 29850 221320 32028
rect 221280 29844 221332 29850
rect 221280 29786 221332 29792
rect 222108 29844 222160 29850
rect 222108 29786 222160 29792
rect 220176 29776 220228 29782
rect 220176 29718 220228 29724
rect 220728 29096 220780 29102
rect 220728 29038 220780 29044
rect 220740 6914 220768 29038
rect 219268 6886 219388 6914
rect 220464 6886 220768 6914
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213828 3528 213880 3534
rect 213828 3470 213880 3476
rect 214472 3528 214524 3534
rect 214472 3470 214524 3476
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 216864 3528 216916 3534
rect 216864 3470 216916 3476
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 219164 3528 219216 3534
rect 219164 3470 219216 3476
rect 213380 480 213408 3470
rect 214484 480 214512 3470
rect 215680 480 215708 3470
rect 216876 480 216904 3470
rect 218072 480 218100 3470
rect 219268 480 219296 6886
rect 220464 480 220492 6886
rect 222120 3330 222148 29786
rect 222304 29646 222332 32028
rect 223408 29986 223436 32028
rect 223488 30252 223540 30258
rect 223488 30194 223540 30200
rect 223396 29980 223448 29986
rect 223396 29922 223448 29928
rect 222292 29640 222344 29646
rect 222292 29582 222344 29588
rect 223500 3534 223528 30194
rect 224420 30190 224448 32028
rect 224868 30320 224920 30326
rect 224868 30262 224920 30268
rect 224408 30184 224460 30190
rect 224408 30126 224460 30132
rect 224880 3534 224908 30262
rect 225524 30122 225552 32028
rect 225512 30116 225564 30122
rect 225512 30058 225564 30064
rect 226248 30116 226300 30122
rect 226248 30058 226300 30064
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 221556 3324 221608 3330
rect 221556 3266 221608 3272
rect 222108 3324 222160 3330
rect 222108 3266 222160 3272
rect 221568 480 221596 3266
rect 222764 480 222792 3470
rect 223960 480 223988 3470
rect 226260 3262 226288 30058
rect 226536 29714 226564 32028
rect 227444 29980 227496 29986
rect 227444 29922 227496 29928
rect 226524 29708 226576 29714
rect 226524 29650 226576 29656
rect 225144 3256 225196 3262
rect 225144 3198 225196 3204
rect 226248 3256 226300 3262
rect 226248 3198 226300 3204
rect 225156 480 225184 3198
rect 227456 3058 227484 29922
rect 227548 29918 227576 32028
rect 227536 29912 227588 29918
rect 227536 29854 227588 29860
rect 227628 29912 227680 29918
rect 227628 29854 227680 29860
rect 227640 6914 227668 29854
rect 228652 29102 228680 32028
rect 229664 29850 229692 32028
rect 230768 30258 230796 32028
rect 231780 30326 231808 32028
rect 231768 30320 231820 30326
rect 231768 30262 231820 30268
rect 230756 30252 230808 30258
rect 230756 30194 230808 30200
rect 232884 30122 232912 32028
rect 232872 30116 232924 30122
rect 232872 30058 232924 30064
rect 233148 30116 233200 30122
rect 233148 30058 233200 30064
rect 229652 29844 229704 29850
rect 229652 29786 229704 29792
rect 229008 29708 229060 29714
rect 229008 29650 229060 29656
rect 228640 29096 228692 29102
rect 228640 29038 228692 29044
rect 229020 6914 229048 29650
rect 230388 29164 230440 29170
rect 230388 29106 230440 29112
rect 227548 6886 227668 6914
rect 228744 6886 229048 6914
rect 226340 3052 226392 3058
rect 226340 2994 226392 3000
rect 227444 3052 227496 3058
rect 227444 2994 227496 3000
rect 226352 480 226380 2994
rect 227548 480 227576 6886
rect 228744 480 228772 6886
rect 230400 3534 230428 29106
rect 231768 29028 231820 29034
rect 231768 28970 231820 28976
rect 231780 3534 231808 28970
rect 233160 3534 233188 30058
rect 233896 29986 233924 32028
rect 233884 29980 233936 29986
rect 233884 29922 233936 29928
rect 235000 29918 235028 32028
rect 234988 29912 235040 29918
rect 234988 29854 235040 29860
rect 236012 29714 236040 32028
rect 236000 29708 236052 29714
rect 236000 29650 236052 29656
rect 235816 29640 235868 29646
rect 235816 29582 235868 29588
rect 234528 29300 234580 29306
rect 234528 29242 234580 29248
rect 234540 3534 234568 29242
rect 229836 3528 229888 3534
rect 229836 3470 229888 3476
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 229848 480 229876 3470
rect 231044 480 231072 3470
rect 232240 480 232268 3470
rect 233436 480 233464 3470
rect 234632 480 234660 3470
rect 235828 480 235856 29582
rect 235908 29572 235960 29578
rect 235908 29514 235960 29520
rect 235920 3534 235948 29514
rect 237116 29170 237144 32028
rect 237288 29708 237340 29714
rect 237288 29650 237340 29656
rect 237104 29164 237156 29170
rect 237104 29106 237156 29112
rect 237300 6914 237328 29650
rect 238128 29034 238156 32028
rect 239232 30122 239260 32028
rect 239220 30116 239272 30122
rect 239220 30058 239272 30064
rect 238668 29776 238720 29782
rect 238668 29718 238720 29724
rect 238116 29028 238168 29034
rect 238116 28970 238168 28976
rect 237024 6886 237328 6914
rect 235908 3528 235960 3534
rect 235908 3470 235960 3476
rect 237024 480 237052 6886
rect 238680 3534 238708 29718
rect 240244 29306 240272 32028
rect 241256 29578 241284 32028
rect 242360 29646 242388 32028
rect 243372 29714 243400 32028
rect 244096 30320 244148 30326
rect 244096 30262 244148 30268
rect 243360 29708 243412 29714
rect 243360 29650 243412 29656
rect 242348 29640 242400 29646
rect 242348 29582 242400 29588
rect 241244 29572 241296 29578
rect 241244 29514 241296 29520
rect 240232 29300 240284 29306
rect 240232 29242 240284 29248
rect 241428 29232 241480 29238
rect 241428 29174 241480 29180
rect 240048 29164 240100 29170
rect 240048 29106 240100 29112
rect 240060 3534 240088 29106
rect 241440 3534 241468 29174
rect 242808 29096 242860 29102
rect 242808 29038 242860 29044
rect 238116 3528 238168 3534
rect 238116 3470 238168 3476
rect 238668 3528 238720 3534
rect 238668 3470 238720 3476
rect 239312 3528 239364 3534
rect 239312 3470 239364 3476
rect 240048 3528 240100 3534
rect 240048 3470 240100 3476
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 238128 480 238156 3470
rect 239324 480 239352 3470
rect 240520 480 240548 3470
rect 242820 3194 242848 29038
rect 244108 16574 244136 30262
rect 244188 30184 244240 30190
rect 244188 30126 244240 30132
rect 244016 16546 244136 16574
rect 244016 3534 244044 16546
rect 244200 6914 244228 30126
rect 244476 29782 244504 32028
rect 244464 29776 244516 29782
rect 244464 29718 244516 29724
rect 245488 29170 245516 32028
rect 246592 29238 246620 32028
rect 246948 29708 247000 29714
rect 246948 29650 247000 29656
rect 246580 29232 246632 29238
rect 246580 29174 246632 29180
rect 245476 29164 245528 29170
rect 245476 29106 245528 29112
rect 245568 29164 245620 29170
rect 245568 29106 245620 29112
rect 244108 6886 244228 6914
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 244004 3528 244056 3534
rect 244004 3470 244056 3476
rect 241704 3188 241756 3194
rect 241704 3130 241756 3136
rect 242808 3188 242860 3194
rect 242808 3130 242860 3136
rect 241716 480 241744 3130
rect 242912 480 242940 3470
rect 244108 480 244136 6886
rect 245212 598 245424 626
rect 245212 480 245240 598
rect 245396 490 245424 598
rect 245580 490 245608 29106
rect 246960 3126 246988 29650
rect 247604 29102 247632 32028
rect 248708 30326 248736 32028
rect 248696 30320 248748 30326
rect 248696 30262 248748 30268
rect 249720 30190 249748 32028
rect 249708 30184 249760 30190
rect 249708 30126 249760 30132
rect 248328 29912 248380 29918
rect 248328 29854 248380 29860
rect 247592 29096 247644 29102
rect 247592 29038 247644 29044
rect 248340 3534 248368 29854
rect 249708 29232 249760 29238
rect 249708 29174 249760 29180
rect 247592 3528 247644 3534
rect 247592 3470 247644 3476
rect 248328 3528 248380 3534
rect 248328 3470 248380 3476
rect 246396 3120 246448 3126
rect 246396 3062 246448 3068
rect 246948 3120 247000 3126
rect 246948 3062 247000 3068
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245396 462 245608 490
rect 246408 480 246436 3062
rect 247604 480 247632 3470
rect 249720 3058 249748 29174
rect 250824 29170 250852 32028
rect 251836 29714 251864 32028
rect 252940 29918 252968 32028
rect 253848 30252 253900 30258
rect 253848 30194 253900 30200
rect 252928 29912 252980 29918
rect 252928 29854 252980 29860
rect 251824 29708 251876 29714
rect 251824 29650 251876 29656
rect 250812 29164 250864 29170
rect 250812 29106 250864 29112
rect 252468 29164 252520 29170
rect 252468 29106 252520 29112
rect 251088 29096 251140 29102
rect 251088 29038 251140 29044
rect 251100 3534 251128 29038
rect 252376 29028 252428 29034
rect 252376 28970 252428 28976
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 248788 3052 248840 3058
rect 248788 2994 248840 3000
rect 249708 3052 249760 3058
rect 249708 2994 249760 3000
rect 248800 480 248828 2994
rect 249996 480 250024 3470
rect 251192 480 251220 3470
rect 252388 480 252416 28970
rect 252480 3534 252508 29106
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 253492 598 253704 626
rect 253492 480 253520 598
rect 253676 490 253704 598
rect 253860 490 253888 30194
rect 253952 29238 253980 32028
rect 253940 29232 253992 29238
rect 253940 29174 253992 29180
rect 255056 29102 255084 32028
rect 255228 30320 255280 30326
rect 255228 30262 255280 30268
rect 255044 29096 255096 29102
rect 255044 29038 255096 29044
rect 255240 3534 255268 30262
rect 256068 29170 256096 32028
rect 256608 29776 256660 29782
rect 256608 29718 256660 29724
rect 256056 29164 256108 29170
rect 256056 29106 256108 29112
rect 256620 3534 256648 29718
rect 257080 29034 257108 32028
rect 258184 30258 258212 32028
rect 259196 30326 259224 32028
rect 259184 30320 259236 30326
rect 259184 30262 259236 30268
rect 258172 30252 258224 30258
rect 258172 30194 258224 30200
rect 257988 29912 258040 29918
rect 257988 29854 258040 29860
rect 257068 29028 257120 29034
rect 257068 28970 257120 28976
rect 258000 3534 258028 29854
rect 260300 29782 260328 32028
rect 261312 29918 261340 32028
rect 261300 29912 261352 29918
rect 261300 29854 261352 29860
rect 260288 29776 260340 29782
rect 260288 29718 260340 29724
rect 262128 29232 262180 29238
rect 262128 29174 262180 29180
rect 260656 29164 260708 29170
rect 260656 29106 260708 29112
rect 259368 29096 259420 29102
rect 259368 29038 259420 29044
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 255228 3528 255280 3534
rect 255228 3470 255280 3476
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 256608 3528 256660 3534
rect 256608 3470 256660 3476
rect 257068 3528 257120 3534
rect 257068 3470 257120 3476
rect 257988 3528 258040 3534
rect 257988 3470 258040 3476
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 253676 462 253888 490
rect 254688 480 254716 3470
rect 255884 480 255912 3470
rect 257080 480 257108 3470
rect 259380 3262 259408 29038
rect 260668 16574 260696 29106
rect 260748 29028 260800 29034
rect 260748 28970 260800 28976
rect 260576 16546 260696 16574
rect 258264 3256 258316 3262
rect 258264 3198 258316 3204
rect 259368 3256 259420 3262
rect 259368 3198 259420 3204
rect 258276 480 258304 3198
rect 260576 3058 260604 16546
rect 260760 6914 260788 28970
rect 260668 6886 260788 6914
rect 259460 3052 259512 3058
rect 259460 2994 259512 3000
rect 260564 3052 260616 3058
rect 260564 2994 260616 3000
rect 259472 480 259500 2994
rect 260668 480 260696 6886
rect 261772 598 261984 626
rect 261772 480 261800 598
rect 261956 490 261984 598
rect 262140 490 262168 29174
rect 262416 29102 262444 32028
rect 263428 29170 263456 32028
rect 263416 29164 263468 29170
rect 263416 29106 263468 29112
rect 262404 29096 262456 29102
rect 262404 29038 262456 29044
rect 263508 29096 263560 29102
rect 263508 29038 263560 29044
rect 263520 3330 263548 29038
rect 264532 29034 264560 32028
rect 265544 29238 265572 32028
rect 266268 29504 266320 29510
rect 266268 29446 266320 29452
rect 265532 29232 265584 29238
rect 265532 29174 265584 29180
rect 264888 29164 264940 29170
rect 264888 29106 264940 29112
rect 264520 29028 264572 29034
rect 264520 28970 264572 28976
rect 264900 3534 264928 29106
rect 266280 3534 266308 29446
rect 266648 29102 266676 32028
rect 267556 29300 267608 29306
rect 267556 29242 267608 29248
rect 266636 29096 266688 29102
rect 266636 29038 266688 29044
rect 267568 3534 267596 29242
rect 267660 29170 267688 32028
rect 268764 29510 268792 32028
rect 268752 29504 268804 29510
rect 268752 29446 268804 29452
rect 269776 29306 269804 32028
rect 269764 29300 269816 29306
rect 269764 29242 269816 29248
rect 270408 29232 270460 29238
rect 270408 29174 270460 29180
rect 267648 29164 267700 29170
rect 267648 29106 267700 29112
rect 269028 29096 269080 29102
rect 269028 29038 269080 29044
rect 268936 29028 268988 29034
rect 268936 28970 268988 28976
rect 268948 6914 268976 28970
rect 268856 6886 268976 6914
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 264888 3528 264940 3534
rect 264888 3470 264940 3476
rect 265348 3528 265400 3534
rect 265348 3470 265400 3476
rect 266268 3528 266320 3534
rect 266268 3470 266320 3476
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 267556 3528 267608 3534
rect 267556 3470 267608 3476
rect 267740 3528 267792 3534
rect 267740 3470 267792 3476
rect 262956 3324 263008 3330
rect 262956 3266 263008 3272
rect 263508 3324 263560 3330
rect 263508 3266 263560 3272
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 261956 462 262168 490
rect 262968 480 262996 3266
rect 264164 480 264192 3470
rect 265360 480 265388 3470
rect 266556 480 266584 3470
rect 267752 480 267780 3470
rect 268856 480 268884 6886
rect 269040 3534 269068 29038
rect 269028 3528 269080 3534
rect 269028 3470 269080 3476
rect 270052 598 270264 626
rect 270052 480 270080 598
rect 270236 490 270264 598
rect 270420 490 270448 29174
rect 270788 29102 270816 32028
rect 271788 29164 271840 29170
rect 271788 29106 271840 29112
rect 270776 29096 270828 29102
rect 270776 29038 270828 29044
rect 271800 3330 271828 29106
rect 271892 29034 271920 32028
rect 272904 29238 272932 32028
rect 272892 29232 272944 29238
rect 272892 29174 272944 29180
rect 274008 29170 274036 32028
rect 273996 29164 274048 29170
rect 273996 29106 274048 29112
rect 274548 29164 274600 29170
rect 274548 29106 274600 29112
rect 273904 29096 273956 29102
rect 273904 29038 273956 29044
rect 271880 29028 271932 29034
rect 271880 28970 271932 28976
rect 273628 3528 273680 3534
rect 273628 3470 273680 3476
rect 272432 3460 272484 3466
rect 272432 3402 272484 3408
rect 271236 3324 271288 3330
rect 271236 3266 271288 3272
rect 271788 3324 271840 3330
rect 271788 3266 271840 3272
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270236 462 270448 490
rect 271248 480 271276 3266
rect 272444 480 272472 3402
rect 273640 480 273668 3470
rect 273916 3466 273944 29038
rect 274560 3534 274588 29106
rect 275020 29102 275048 32028
rect 276124 29170 276152 32028
rect 276112 29164 276164 29170
rect 276112 29106 276164 29112
rect 275008 29096 275060 29102
rect 275008 29038 275060 29044
rect 277136 16574 277164 32028
rect 278240 30326 278268 32028
rect 277308 30320 277360 30326
rect 277308 30262 277360 30268
rect 278228 30320 278280 30326
rect 278228 30262 278280 30268
rect 277216 29164 277268 29170
rect 277216 29106 277268 29112
rect 277044 16546 277164 16574
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 276020 3528 276072 3534
rect 276020 3470 276072 3476
rect 273904 3460 273956 3466
rect 273904 3402 273956 3408
rect 274824 3052 274876 3058
rect 274824 2994 274876 3000
rect 274836 480 274864 2994
rect 276032 480 276060 3470
rect 277044 3058 277072 16546
rect 277228 6914 277256 29106
rect 277136 6886 277256 6914
rect 277032 3052 277084 3058
rect 277032 2994 277084 3000
rect 277136 480 277164 6886
rect 277320 3534 277348 30262
rect 279252 29170 279280 32028
rect 279240 29164 279292 29170
rect 279240 29106 279292 29112
rect 280356 29102 280384 32028
rect 278688 29096 278740 29102
rect 278688 29038 278740 29044
rect 280344 29096 280396 29102
rect 280344 29038 280396 29044
rect 277308 3528 277360 3534
rect 277308 3470 277360 3476
rect 278332 598 278544 626
rect 278332 480 278360 598
rect 278516 490 278544 598
rect 278700 490 278728 29038
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 279516 3460 279568 3466
rect 279516 3402 279568 3408
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 278516 462 278728 490
rect 279528 480 279556 3402
rect 280724 480 280752 3470
rect 281368 3466 281396 32028
rect 282472 29170 282500 32028
rect 281448 29164 281500 29170
rect 281448 29106 281500 29112
rect 282460 29164 282512 29170
rect 282460 29106 282512 29112
rect 281460 3534 281488 29106
rect 283484 29034 283512 32028
rect 282828 29028 282880 29034
rect 282828 28970 282880 28976
rect 283472 29028 283524 29034
rect 283472 28970 283524 28976
rect 282840 3534 282868 28970
rect 284588 3534 284616 32028
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 281908 3528 281960 3534
rect 281908 3470 281960 3476
rect 282828 3528 282880 3534
rect 282828 3470 282880 3476
rect 283104 3528 283156 3534
rect 283104 3470 283156 3476
rect 284576 3528 284628 3534
rect 284576 3470 284628 3476
rect 285404 3528 285456 3534
rect 285404 3470 285456 3476
rect 281356 3460 281408 3466
rect 281356 3402 281408 3408
rect 281920 480 281948 3470
rect 283116 480 283144 3470
rect 284300 3052 284352 3058
rect 284300 2994 284352 3000
rect 284312 480 284340 2994
rect 285416 480 285444 3470
rect 285600 3058 285628 32028
rect 286612 3534 286640 32028
rect 287716 30326 287744 32028
rect 286968 30320 287020 30326
rect 286968 30262 287020 30268
rect 287704 30320 287756 30326
rect 287704 30262 287756 30268
rect 286600 3528 286652 3534
rect 286600 3470 286652 3476
rect 285588 3052 285640 3058
rect 285588 2994 285640 3000
rect 286612 598 286824 626
rect 286612 480 286640 598
rect 286796 490 286824 598
rect 286980 490 287008 30262
rect 288728 29186 288756 32028
rect 289832 29186 289860 32028
rect 288360 29158 288756 29186
rect 289740 29158 289860 29186
rect 290844 29170 290872 32028
rect 289912 29164 289964 29170
rect 288360 3330 288388 29158
rect 289740 3534 289768 29158
rect 289912 29106 289964 29112
rect 290832 29164 290884 29170
rect 290832 29106 290884 29112
rect 289924 16574 289952 29106
rect 289924 16546 290228 16574
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 287796 3324 287848 3330
rect 287796 3266 287848 3272
rect 288348 3324 288400 3330
rect 288348 3266 288400 3272
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 286796 462 287008 490
rect 287808 480 287836 3266
rect 289004 480 289032 3470
rect 290200 480 290228 16546
rect 291948 3534 291976 32028
rect 292960 6914 292988 32028
rect 294064 29186 294092 32028
rect 293880 29158 294092 29186
rect 293880 6914 293908 29158
rect 295076 6914 295104 32028
rect 296180 6914 296208 32028
rect 297192 29170 297220 32028
rect 296720 29164 296772 29170
rect 296720 29106 296772 29112
rect 297180 29164 297232 29170
rect 297180 29106 297232 29112
rect 296732 16574 296760 29106
rect 298296 16574 298324 32028
rect 299308 26234 299336 32028
rect 300320 29170 300348 32028
rect 299572 29164 299624 29170
rect 299572 29106 299624 29112
rect 300308 29164 300360 29170
rect 300308 29106 300360 29112
rect 299308 26206 299428 26234
rect 296732 16546 297312 16574
rect 298296 16546 298508 16574
rect 292592 6886 292988 6914
rect 293696 6886 293908 6914
rect 294892 6886 295104 6914
rect 296088 6886 296208 6914
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 291936 3528 291988 3534
rect 291936 3470 291988 3476
rect 291396 480 291424 3470
rect 292592 480 292620 6886
rect 293696 480 293724 6886
rect 294892 480 294920 6886
rect 296088 480 296116 6886
rect 297284 480 297312 16546
rect 298480 480 298508 16546
rect 299400 3210 299428 26206
rect 299584 11762 299612 29106
rect 299572 11756 299624 11762
rect 299572 11698 299624 11704
rect 300768 11756 300820 11762
rect 300768 11698 300820 11704
rect 299400 3182 299704 3210
rect 299676 480 299704 3182
rect 300780 480 300808 11698
rect 301424 3534 301452 32028
rect 301412 3528 301464 3534
rect 301412 3470 301464 3476
rect 301964 3528 302016 3534
rect 301964 3470 302016 3476
rect 301976 480 302004 3470
rect 302436 3058 302464 32028
rect 303540 3534 303568 32028
rect 304552 26234 304580 32028
rect 305656 29170 305684 32028
rect 306668 29170 306696 32028
rect 305644 29164 305696 29170
rect 305644 29106 305696 29112
rect 306288 29164 306340 29170
rect 306288 29106 306340 29112
rect 306656 29164 306708 29170
rect 306656 29106 306708 29112
rect 307668 29164 307720 29170
rect 307668 29106 307720 29112
rect 304552 26206 304948 26234
rect 304920 3534 304948 26206
rect 303528 3528 303580 3534
rect 303528 3470 303580 3476
rect 304356 3528 304408 3534
rect 304356 3470 304408 3476
rect 304908 3528 304960 3534
rect 304908 3470 304960 3476
rect 305552 3528 305604 3534
rect 305552 3470 305604 3476
rect 302424 3052 302476 3058
rect 302424 2994 302476 3000
rect 303160 3052 303212 3058
rect 303160 2994 303212 3000
rect 303172 480 303200 2994
rect 304368 480 304396 3470
rect 305564 480 305592 3470
rect 306300 2802 306328 29106
rect 307680 3482 307708 29106
rect 307772 3602 307800 32028
rect 308784 29186 308812 32028
rect 308784 29158 309180 29186
rect 309888 29170 309916 32028
rect 310900 29170 310928 32028
rect 309152 16574 309180 29158
rect 309876 29164 309928 29170
rect 309876 29106 309928 29112
rect 310428 29164 310480 29170
rect 310428 29106 310480 29112
rect 310888 29164 310940 29170
rect 310888 29106 310940 29112
rect 311808 29164 311860 29170
rect 311808 29106 311860 29112
rect 309152 16546 309824 16574
rect 307760 3596 307812 3602
rect 307760 3538 307812 3544
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 307680 3454 307984 3482
rect 306300 2774 306420 2802
rect 306392 490 306420 2774
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 3454
rect 309060 480 309088 3538
rect 309796 490 309824 16546
rect 310440 3534 310468 29106
rect 311820 3534 311848 29106
rect 312004 29102 312032 32028
rect 311992 29096 312044 29102
rect 311992 29038 312044 29044
rect 313016 26234 313044 32028
rect 313280 29096 313332 29102
rect 313280 29038 313332 29044
rect 313016 26206 313228 26234
rect 310428 3528 310480 3534
rect 310428 3470 310480 3476
rect 311440 3528 311492 3534
rect 311440 3470 311492 3476
rect 311808 3528 311860 3534
rect 311808 3470 311860 3476
rect 312636 3528 312688 3534
rect 312636 3470 312688 3476
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 3470
rect 312648 480 312676 3470
rect 313200 2990 313228 26206
rect 313292 16574 313320 29038
rect 314120 29034 314148 32028
rect 315132 30326 315160 32028
rect 315120 30320 315172 30326
rect 315120 30262 315172 30268
rect 316144 29170 316172 32028
rect 316224 30320 316276 30326
rect 316224 30262 316276 30268
rect 316132 29164 316184 29170
rect 316132 29106 316184 29112
rect 314108 29028 314160 29034
rect 314108 28970 314160 28976
rect 314568 29028 314620 29034
rect 314568 28970 314620 28976
rect 313292 16546 313872 16574
rect 313188 2984 313240 2990
rect 313188 2926 313240 2932
rect 313844 480 313872 16546
rect 314580 4146 314608 28970
rect 316236 16574 316264 30262
rect 316236 16546 317184 16574
rect 314568 4140 314620 4146
rect 314568 4082 314620 4088
rect 316224 4140 316276 4146
rect 316224 4082 316276 4088
rect 315028 2984 315080 2990
rect 315028 2926 315080 2932
rect 315040 480 315068 2926
rect 316236 480 316264 4082
rect 317156 2938 317184 16546
rect 317248 3058 317276 32028
rect 318260 29170 318288 32028
rect 317328 29164 317380 29170
rect 317328 29106 317380 29112
rect 318248 29164 318300 29170
rect 318248 29106 318300 29112
rect 318708 29164 318760 29170
rect 318708 29106 318760 29112
rect 317340 3330 317368 29106
rect 318720 3534 318748 29106
rect 319364 29102 319392 32028
rect 320376 29170 320404 32028
rect 320364 29164 320416 29170
rect 320364 29106 320416 29112
rect 321284 29164 321336 29170
rect 321284 29106 321336 29112
rect 319352 29096 319404 29102
rect 319352 29038 319404 29044
rect 321296 3534 321324 29106
rect 321480 26234 321508 32028
rect 321560 29096 321612 29102
rect 321560 29038 321612 29044
rect 321388 26206 321508 26234
rect 318708 3528 318760 3534
rect 318708 3470 318760 3476
rect 320916 3528 320968 3534
rect 320916 3470 320968 3476
rect 321284 3528 321336 3534
rect 321284 3470 321336 3476
rect 317328 3324 317380 3330
rect 317328 3266 317380 3272
rect 318524 3324 318576 3330
rect 318524 3266 318576 3272
rect 317236 3052 317288 3058
rect 317236 2994 317288 3000
rect 317156 2910 317368 2938
rect 317340 480 317368 2910
rect 318536 480 318564 3266
rect 319720 3052 319772 3058
rect 319720 2994 319772 3000
rect 319732 480 319760 2994
rect 320928 480 320956 3470
rect 321388 3194 321416 26206
rect 321572 16574 321600 29038
rect 322492 26234 322520 32028
rect 323596 29170 323624 32028
rect 323584 29164 323636 29170
rect 323584 29106 323636 29112
rect 324228 29164 324280 29170
rect 324228 29106 324280 29112
rect 322492 26206 322888 26234
rect 321572 16546 322152 16574
rect 321376 3188 321428 3194
rect 321376 3130 321428 3136
rect 322124 480 322152 16546
rect 322860 3058 322888 26206
rect 324240 3670 324268 29106
rect 324608 29102 324636 32028
rect 324596 29096 324648 29102
rect 324596 29038 324648 29044
rect 325608 29096 325660 29102
rect 325608 29038 325660 29044
rect 325620 4146 325648 29038
rect 325712 29034 325740 32028
rect 325700 29028 325752 29034
rect 325700 28970 325752 28976
rect 326724 26234 326752 32028
rect 327828 29170 327856 32028
rect 328840 29170 328868 32028
rect 329852 29170 329880 32028
rect 327816 29164 327868 29170
rect 327816 29106 327868 29112
rect 328368 29164 328420 29170
rect 328368 29106 328420 29112
rect 328828 29164 328880 29170
rect 328828 29106 328880 29112
rect 329748 29164 329800 29170
rect 329748 29106 329800 29112
rect 329840 29164 329892 29170
rect 329840 29106 329892 29112
rect 327724 29028 327776 29034
rect 327724 28970 327776 28976
rect 326724 26206 327028 26234
rect 325608 4140 325660 4146
rect 325608 4082 325660 4088
rect 324228 3664 324280 3670
rect 324228 3606 324280 3612
rect 326804 3664 326856 3670
rect 326804 3606 326856 3612
rect 323308 3528 323360 3534
rect 323308 3470 323360 3476
rect 322848 3052 322900 3058
rect 322848 2994 322900 3000
rect 323320 480 323348 3470
rect 324412 3188 324464 3194
rect 324412 3130 324464 3136
rect 324424 480 324452 3130
rect 325608 3052 325660 3058
rect 325608 2994 325660 3000
rect 325620 480 325648 2994
rect 326816 480 326844 3606
rect 327000 3602 327028 26206
rect 326988 3596 327040 3602
rect 326988 3538 327040 3544
rect 327736 3534 327764 28970
rect 328000 4140 328052 4146
rect 328000 4082 328052 4088
rect 327724 3528 327776 3534
rect 327724 3470 327776 3476
rect 328012 480 328040 4082
rect 328380 3466 328408 29106
rect 329196 3528 329248 3534
rect 329196 3470 329248 3476
rect 328368 3460 328420 3466
rect 328368 3402 328420 3408
rect 329208 480 329236 3470
rect 329760 3194 329788 29106
rect 330956 26234 330984 32028
rect 331968 29170 331996 32028
rect 333072 29170 333100 32028
rect 334084 29170 334112 32028
rect 331128 29164 331180 29170
rect 331128 29106 331180 29112
rect 331956 29164 332008 29170
rect 331956 29106 332008 29112
rect 332508 29164 332560 29170
rect 332508 29106 332560 29112
rect 333060 29164 333112 29170
rect 333060 29106 333112 29112
rect 333888 29164 333940 29170
rect 333888 29106 333940 29112
rect 334072 29164 334124 29170
rect 334072 29106 334124 29112
rect 335084 29164 335136 29170
rect 335084 29106 335136 29112
rect 330956 26206 331076 26234
rect 330392 3596 330444 3602
rect 330392 3538 330444 3544
rect 329748 3188 329800 3194
rect 329748 3130 329800 3136
rect 330404 480 330432 3538
rect 331048 3398 331076 26206
rect 331140 3534 331168 29106
rect 332520 3670 332548 29106
rect 333900 4010 333928 29106
rect 333888 4004 333940 4010
rect 333888 3946 333940 3952
rect 332508 3664 332560 3670
rect 332508 3606 332560 3612
rect 335096 3534 335124 29106
rect 335188 26234 335216 32028
rect 336200 29170 336228 32028
rect 337304 29170 337332 32028
rect 338316 29170 338344 32028
rect 336188 29164 336240 29170
rect 336188 29106 336240 29112
rect 336648 29164 336700 29170
rect 336648 29106 336700 29112
rect 337292 29164 337344 29170
rect 337292 29106 337344 29112
rect 338028 29164 338080 29170
rect 338028 29106 338080 29112
rect 338304 29164 338356 29170
rect 338304 29106 338356 29112
rect 339316 29164 339368 29170
rect 339316 29106 339368 29112
rect 335188 26206 335308 26234
rect 335280 3602 335308 26206
rect 336280 3664 336332 3670
rect 336280 3606 336332 3612
rect 335268 3596 335320 3602
rect 335268 3538 335320 3544
rect 331128 3528 331180 3534
rect 331128 3470 331180 3476
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 335084 3528 335136 3534
rect 335084 3470 335136 3476
rect 331588 3460 331640 3466
rect 331588 3402 331640 3408
rect 331036 3392 331088 3398
rect 331036 3334 331088 3340
rect 331600 480 331628 3402
rect 332692 3188 332744 3194
rect 332692 3130 332744 3136
rect 332704 480 332732 3130
rect 333900 480 333928 3470
rect 335084 3392 335136 3398
rect 335084 3334 335136 3340
rect 335096 480 335124 3334
rect 336292 480 336320 3606
rect 336660 3262 336688 29106
rect 337476 4004 337528 4010
rect 337476 3946 337528 3952
rect 336648 3256 336700 3262
rect 336648 3198 336700 3204
rect 337488 480 337516 3946
rect 338040 3466 338068 29106
rect 338672 3528 338724 3534
rect 338672 3470 338724 3476
rect 338028 3460 338080 3466
rect 338028 3402 338080 3408
rect 338684 480 338712 3470
rect 339328 3330 339356 29106
rect 339420 3534 339448 32028
rect 340432 26234 340460 32028
rect 341536 29170 341564 32028
rect 342548 29170 342576 32028
rect 341524 29164 341576 29170
rect 341524 29106 341576 29112
rect 342168 29164 342220 29170
rect 342168 29106 342220 29112
rect 342536 29164 342588 29170
rect 342536 29106 342588 29112
rect 343548 29164 343600 29170
rect 343548 29106 343600 29112
rect 340432 26206 340828 26234
rect 340800 4078 340828 26206
rect 342180 4146 342208 29106
rect 342168 4140 342220 4146
rect 342168 4082 342220 4088
rect 340788 4072 340840 4078
rect 340788 4014 340840 4020
rect 339868 3596 339920 3602
rect 339868 3538 339920 3544
rect 339408 3528 339460 3534
rect 339408 3470 339460 3476
rect 339316 3324 339368 3330
rect 339316 3266 339368 3272
rect 339880 480 339908 3538
rect 343560 3466 343588 29106
rect 343652 29034 343680 32028
rect 344664 29152 344692 32028
rect 345676 29170 345704 32028
rect 346780 29170 346808 32028
rect 345664 29164 345716 29170
rect 344664 29124 344968 29152
rect 343640 29028 343692 29034
rect 343640 28970 343692 28976
rect 344836 29028 344888 29034
rect 344836 28970 344888 28976
rect 344848 3534 344876 28970
rect 344940 3806 344968 29124
rect 345664 29106 345716 29112
rect 346308 29164 346360 29170
rect 346308 29106 346360 29112
rect 346768 29164 346820 29170
rect 346768 29106 346820 29112
rect 347688 29164 347740 29170
rect 347688 29106 347740 29112
rect 345756 4072 345808 4078
rect 345756 4014 345808 4020
rect 344928 3800 344980 3806
rect 344928 3742 344980 3748
rect 344560 3528 344612 3534
rect 344560 3470 344612 3476
rect 344836 3528 344888 3534
rect 344836 3470 344888 3476
rect 342168 3460 342220 3466
rect 342168 3402 342220 3408
rect 343548 3460 343600 3466
rect 343548 3402 343600 3408
rect 340972 3256 341024 3262
rect 340972 3198 341024 3204
rect 340984 480 341012 3198
rect 342180 480 342208 3402
rect 343364 3324 343416 3330
rect 343364 3266 343416 3272
rect 343376 480 343404 3266
rect 344572 480 344600 3470
rect 345768 480 345796 4014
rect 346320 3262 346348 29106
rect 346952 4140 347004 4146
rect 346952 4082 347004 4088
rect 346308 3256 346360 3262
rect 346308 3198 346360 3204
rect 346964 480 346992 4082
rect 347700 3330 347728 29106
rect 347792 29102 347820 32028
rect 348896 29186 348924 32028
rect 348896 29158 349108 29186
rect 347780 29096 347832 29102
rect 347780 29038 347832 29044
rect 348976 29096 349028 29102
rect 348976 29038 349028 29044
rect 348988 3466 349016 29038
rect 348056 3460 348108 3466
rect 348056 3402 348108 3408
rect 348976 3460 349028 3466
rect 348976 3402 349028 3408
rect 347688 3324 347740 3330
rect 347688 3266 347740 3272
rect 348068 480 348096 3402
rect 349080 2922 349108 29158
rect 349908 29034 349936 32028
rect 351012 29170 351040 32028
rect 352024 29170 352052 32028
rect 351000 29164 351052 29170
rect 351000 29106 351052 29112
rect 351828 29164 351880 29170
rect 351828 29106 351880 29112
rect 352012 29164 352064 29170
rect 352012 29106 352064 29112
rect 349896 29028 349948 29034
rect 349896 28970 349948 28976
rect 350448 29028 350500 29034
rect 350448 28970 350500 28976
rect 350460 4146 350488 28970
rect 350448 4140 350500 4146
rect 350448 4082 350500 4088
rect 351840 3806 351868 29106
rect 350448 3800 350500 3806
rect 350448 3742 350500 3748
rect 351828 3800 351880 3806
rect 351828 3742 351880 3748
rect 349252 3528 349304 3534
rect 349252 3470 349304 3476
rect 349068 2916 349120 2922
rect 349068 2858 349120 2864
rect 349264 480 349292 3470
rect 350460 480 350488 3742
rect 353128 3602 353156 32028
rect 354140 29170 354168 32028
rect 353208 29164 353260 29170
rect 353208 29106 353260 29112
rect 354128 29164 354180 29170
rect 354128 29106 354180 29112
rect 354588 29164 354640 29170
rect 354588 29106 354640 29112
rect 353220 4010 353248 29106
rect 353208 4004 353260 4010
rect 353208 3946 353260 3952
rect 354600 3738 354628 29106
rect 355244 29102 355272 32028
rect 356256 29170 356284 32028
rect 356244 29164 356296 29170
rect 356244 29106 356296 29112
rect 357256 29164 357308 29170
rect 357256 29106 357308 29112
rect 355232 29096 355284 29102
rect 355232 29038 355284 29044
rect 355968 29096 356020 29102
rect 355968 29038 356020 29044
rect 354588 3732 354640 3738
rect 354588 3674 354640 3680
rect 353116 3596 353168 3602
rect 353116 3538 353168 3544
rect 354036 3460 354088 3466
rect 354036 3402 354088 3408
rect 352840 3324 352892 3330
rect 352840 3266 352892 3272
rect 351644 3256 351696 3262
rect 351644 3198 351696 3204
rect 351656 480 351684 3198
rect 352852 480 352880 3266
rect 354048 480 354076 3402
rect 355980 3330 356008 29038
rect 356336 4140 356388 4146
rect 356336 4082 356388 4088
rect 355968 3324 356020 3330
rect 355968 3266 356020 3272
rect 355232 2916 355284 2922
rect 355232 2858 355284 2864
rect 355244 480 355272 2858
rect 356348 480 356376 4082
rect 357268 3534 357296 29106
rect 357360 3670 357388 32028
rect 358372 26234 358400 32028
rect 359384 29170 359412 32028
rect 360488 29170 360516 32028
rect 359372 29164 359424 29170
rect 359372 29106 359424 29112
rect 360108 29164 360160 29170
rect 360108 29106 360160 29112
rect 360476 29164 360528 29170
rect 360476 29106 360528 29112
rect 361396 29164 361448 29170
rect 361396 29106 361448 29112
rect 358372 26206 358768 26234
rect 358740 4146 358768 26206
rect 358728 4140 358780 4146
rect 358728 4082 358780 4088
rect 358728 4004 358780 4010
rect 358728 3946 358780 3952
rect 357532 3800 357584 3806
rect 357532 3742 357584 3748
rect 357348 3664 357400 3670
rect 357348 3606 357400 3612
rect 357256 3528 357308 3534
rect 357256 3470 357308 3476
rect 357544 480 357572 3742
rect 358740 480 358768 3946
rect 359924 3596 359976 3602
rect 359924 3538 359976 3544
rect 359936 480 359964 3538
rect 360120 3126 360148 29106
rect 361408 3806 361436 29106
rect 361396 3800 361448 3806
rect 361396 3742 361448 3748
rect 361500 3738 361528 32028
rect 362604 26234 362632 32028
rect 363616 29170 363644 32028
rect 364720 29170 364748 32028
rect 365732 29170 365760 32028
rect 363604 29164 363656 29170
rect 363604 29106 363656 29112
rect 364248 29164 364300 29170
rect 364248 29106 364300 29112
rect 364708 29164 364760 29170
rect 364708 29106 364760 29112
rect 365628 29164 365680 29170
rect 365628 29106 365680 29112
rect 365720 29164 365772 29170
rect 365720 29106 365772 29112
rect 362604 26206 362908 26234
rect 361120 3732 361172 3738
rect 361120 3674 361172 3680
rect 361488 3732 361540 3738
rect 361488 3674 361540 3680
rect 360108 3120 360160 3126
rect 360108 3062 360160 3068
rect 361132 480 361160 3674
rect 362880 3602 362908 26206
rect 362868 3596 362920 3602
rect 362868 3538 362920 3544
rect 364260 3534 364288 29106
rect 364616 3664 364668 3670
rect 364616 3606 364668 3612
rect 363512 3528 363564 3534
rect 363512 3470 363564 3476
rect 364248 3528 364300 3534
rect 364248 3470 364300 3476
rect 362316 3324 362368 3330
rect 362316 3266 362368 3272
rect 362328 480 362356 3266
rect 363524 480 363552 3470
rect 364628 480 364656 3606
rect 365640 2922 365668 29106
rect 366836 26234 366864 32028
rect 367848 29170 367876 32028
rect 368952 29170 368980 32028
rect 369964 29170 369992 32028
rect 367008 29164 367060 29170
rect 367008 29106 367060 29112
rect 367836 29164 367888 29170
rect 367836 29106 367888 29112
rect 368388 29164 368440 29170
rect 368388 29106 368440 29112
rect 368940 29164 368992 29170
rect 368940 29106 368992 29112
rect 369768 29164 369820 29170
rect 369768 29106 369820 29112
rect 369952 29164 370004 29170
rect 369952 29106 370004 29112
rect 370964 29164 371016 29170
rect 370964 29106 371016 29112
rect 366836 26206 366956 26234
rect 365812 4140 365864 4146
rect 365812 4082 365864 4088
rect 365628 2916 365680 2922
rect 365628 2858 365680 2864
rect 365824 480 365852 4082
rect 366928 3466 366956 26206
rect 367020 3874 367048 29106
rect 367008 3868 367060 3874
rect 367008 3810 367060 3816
rect 368204 3800 368256 3806
rect 368204 3742 368256 3748
rect 366916 3460 366968 3466
rect 366916 3402 366968 3408
rect 367008 3120 367060 3126
rect 367008 3062 367060 3068
rect 367020 480 367048 3062
rect 368216 480 368244 3742
rect 368400 3126 368428 29106
rect 369780 4010 369808 29106
rect 369768 4004 369820 4010
rect 369768 3946 369820 3952
rect 369400 3732 369452 3738
rect 369400 3674 369452 3680
rect 368388 3120 368440 3126
rect 368388 3062 368440 3068
rect 369412 480 369440 3674
rect 370976 3670 371004 29106
rect 371068 26234 371096 32028
rect 372080 29170 372108 32028
rect 373184 29170 373212 32028
rect 374196 29170 374224 32028
rect 372068 29164 372120 29170
rect 372068 29106 372120 29112
rect 372528 29164 372580 29170
rect 372528 29106 372580 29112
rect 373172 29164 373224 29170
rect 373172 29106 373224 29112
rect 373908 29164 373960 29170
rect 373908 29106 373960 29112
rect 374184 29164 374236 29170
rect 374184 29106 374236 29112
rect 371068 26206 371188 26234
rect 370964 3664 371016 3670
rect 370964 3606 371016 3612
rect 371160 3602 371188 26206
rect 372540 3738 372568 29106
rect 373920 3942 373948 29106
rect 373908 3936 373960 3942
rect 373908 3878 373960 3884
rect 374092 3868 374144 3874
rect 374092 3810 374144 3816
rect 372528 3732 372580 3738
rect 372528 3674 372580 3680
rect 370596 3596 370648 3602
rect 370596 3538 370648 3544
rect 371148 3596 371200 3602
rect 371148 3538 371200 3544
rect 370608 480 370636 3538
rect 371700 3528 371752 3534
rect 371700 3470 371752 3476
rect 371712 480 371740 3470
rect 372896 2916 372948 2922
rect 372896 2858 372948 2864
rect 372908 480 372936 2858
rect 374104 480 374132 3810
rect 375208 3534 375236 32028
rect 375288 29164 375340 29170
rect 375288 29106 375340 29112
rect 375300 4078 375328 29106
rect 376312 26234 376340 32028
rect 377324 29170 377352 32028
rect 378428 29170 378456 32028
rect 377312 29164 377364 29170
rect 377312 29106 377364 29112
rect 378048 29164 378100 29170
rect 378048 29106 378100 29112
rect 378416 29164 378468 29170
rect 378416 29106 378468 29112
rect 379244 29164 379296 29170
rect 379244 29106 379296 29112
rect 376312 26206 376708 26234
rect 375288 4072 375340 4078
rect 375288 4014 375340 4020
rect 376680 3874 376708 26206
rect 377680 4004 377732 4010
rect 377680 3946 377732 3952
rect 376668 3868 376720 3874
rect 376668 3810 376720 3816
rect 375196 3528 375248 3534
rect 375196 3470 375248 3476
rect 375288 3460 375340 3466
rect 375288 3402 375340 3408
rect 375300 480 375328 3402
rect 376484 3120 376536 3126
rect 376484 3062 376536 3068
rect 376496 480 376524 3062
rect 377692 480 377720 3946
rect 378060 3806 378088 29106
rect 378048 3800 378100 3806
rect 378048 3742 378100 3748
rect 379256 3670 379284 29106
rect 379440 26234 379468 32028
rect 379348 26206 379468 26234
rect 380544 26234 380572 32028
rect 381556 29170 381584 32028
rect 382660 29170 382688 32028
rect 381544 29164 381596 29170
rect 381544 29106 381596 29112
rect 382188 29164 382240 29170
rect 382188 29106 382240 29112
rect 382648 29164 382700 29170
rect 382648 29106 382700 29112
rect 383568 29164 383620 29170
rect 383568 29106 383620 29112
rect 380544 26206 380848 26234
rect 378876 3664 378928 3670
rect 378876 3606 378928 3612
rect 379244 3664 379296 3670
rect 379244 3606 379296 3612
rect 378888 480 378916 3606
rect 379348 3466 379376 26206
rect 380820 3602 380848 26206
rect 382200 4146 382228 29106
rect 382188 4140 382240 4146
rect 382188 4082 382240 4088
rect 383476 4072 383528 4078
rect 383476 4014 383528 4020
rect 382372 3936 382424 3942
rect 382372 3878 382424 3884
rect 381176 3732 381228 3738
rect 381176 3674 381228 3680
rect 379980 3596 380032 3602
rect 379980 3538 380032 3544
rect 380808 3596 380860 3602
rect 380808 3538 380860 3544
rect 379336 3460 379388 3466
rect 379336 3402 379388 3408
rect 379992 480 380020 3538
rect 381188 480 381216 3674
rect 382384 480 382412 3878
rect 383488 3482 383516 4014
rect 383580 4010 383608 29106
rect 383672 29102 383700 32028
rect 384776 29186 384804 32028
rect 384776 29158 384988 29186
rect 383660 29096 383712 29102
rect 383660 29038 383712 29044
rect 384856 29096 384908 29102
rect 384856 29038 384908 29044
rect 384868 4078 384896 29038
rect 384856 4072 384908 4078
rect 384856 4014 384908 4020
rect 383568 4004 383620 4010
rect 383568 3946 383620 3952
rect 384960 3738 384988 29158
rect 385788 29034 385816 32028
rect 386892 29170 386920 32028
rect 387904 29170 387932 32028
rect 386880 29164 386932 29170
rect 386880 29106 386932 29112
rect 387708 29164 387760 29170
rect 387708 29106 387760 29112
rect 387892 29164 387944 29170
rect 387892 29106 387944 29112
rect 388904 29164 388956 29170
rect 388904 29106 388956 29112
rect 385776 29028 385828 29034
rect 385776 28970 385828 28976
rect 386328 29028 386380 29034
rect 386328 28970 386380 28976
rect 386340 3874 386368 28970
rect 387720 3942 387748 29106
rect 387708 3936 387760 3942
rect 387708 3878 387760 3884
rect 385960 3868 386012 3874
rect 385960 3810 386012 3816
rect 386328 3868 386380 3874
rect 386328 3810 386380 3816
rect 384948 3732 385000 3738
rect 384948 3674 385000 3680
rect 384764 3528 384816 3534
rect 383488 3454 383608 3482
rect 384764 3470 384816 3476
rect 383580 480 383608 3454
rect 384776 480 384804 3470
rect 385972 480 386000 3810
rect 387156 3800 387208 3806
rect 387156 3742 387208 3748
rect 387168 480 387196 3742
rect 388260 3664 388312 3670
rect 388260 3606 388312 3612
rect 388272 480 388300 3606
rect 388916 3534 388944 29106
rect 389008 26234 389036 32028
rect 390020 29170 390048 32028
rect 391032 29170 391060 32028
rect 392136 29170 392164 32028
rect 390008 29164 390060 29170
rect 390008 29106 390060 29112
rect 390468 29164 390520 29170
rect 390468 29106 390520 29112
rect 391020 29164 391072 29170
rect 391020 29106 391072 29112
rect 391848 29164 391900 29170
rect 391848 29106 391900 29112
rect 392124 29164 392176 29170
rect 392124 29106 392176 29112
rect 393044 29164 393096 29170
rect 393044 29106 393096 29112
rect 389008 26206 389128 26234
rect 389100 3806 389128 26206
rect 389088 3800 389140 3806
rect 389088 3742 389140 3748
rect 388904 3528 388956 3534
rect 388904 3470 388956 3476
rect 389456 3460 389508 3466
rect 389456 3402 389508 3408
rect 389468 480 389496 3402
rect 390480 3398 390508 29106
rect 391860 6914 391888 29106
rect 391768 6886 391888 6914
rect 390652 3596 390704 3602
rect 390652 3538 390704 3544
rect 390468 3392 390520 3398
rect 390468 3334 390520 3340
rect 390664 480 390692 3538
rect 391768 3330 391796 6886
rect 391848 4140 391900 4146
rect 391848 4082 391900 4088
rect 391756 3324 391808 3330
rect 391756 3266 391808 3272
rect 391860 480 391888 4082
rect 393056 4010 393084 29106
rect 393148 26234 393176 32028
rect 394252 26234 394280 32028
rect 395264 29170 395292 32028
rect 396368 29170 396396 32028
rect 395252 29164 395304 29170
rect 395252 29106 395304 29112
rect 395988 29164 396040 29170
rect 395988 29106 396040 29112
rect 396356 29164 396408 29170
rect 396356 29106 396408 29112
rect 397276 29164 397328 29170
rect 397276 29106 397328 29112
rect 393148 26206 393268 26234
rect 394252 26206 394648 26234
rect 392952 4004 393004 4010
rect 392952 3946 393004 3952
rect 393044 4004 393096 4010
rect 393044 3946 393096 3952
rect 392964 1986 392992 3946
rect 393240 3670 393268 26206
rect 394620 4078 394648 26206
rect 394240 4072 394292 4078
rect 394240 4014 394292 4020
rect 394608 4072 394660 4078
rect 394608 4014 394660 4020
rect 393228 3664 393280 3670
rect 393228 3606 393280 3612
rect 392964 1958 393084 1986
rect 393056 480 393084 1958
rect 394252 480 394280 4014
rect 395344 3732 395396 3738
rect 395344 3674 395396 3680
rect 395356 480 395384 3674
rect 396000 3466 396028 29106
rect 397288 4146 397316 29106
rect 397276 4140 397328 4146
rect 397276 4082 397328 4088
rect 397380 3874 397408 32028
rect 398484 26234 398512 32028
rect 399496 29170 399524 32028
rect 400600 29170 400628 32028
rect 399484 29164 399536 29170
rect 399484 29106 399536 29112
rect 400128 29164 400180 29170
rect 400128 29106 400180 29112
rect 400588 29164 400640 29170
rect 400588 29106 400640 29112
rect 401508 29164 401560 29170
rect 401508 29106 401560 29112
rect 398484 26206 398788 26234
rect 398760 3942 398788 26206
rect 400140 6914 400168 29106
rect 400048 6886 400168 6914
rect 397736 3936 397788 3942
rect 397736 3878 397788 3884
rect 398748 3936 398800 3942
rect 398748 3878 398800 3884
rect 400048 3890 400076 6886
rect 396540 3868 396592 3874
rect 396540 3810 396592 3816
rect 397368 3868 397420 3874
rect 397368 3810 397420 3816
rect 395988 3460 396040 3466
rect 395988 3402 396040 3408
rect 396552 480 396580 3810
rect 397748 480 397776 3878
rect 400048 3862 400352 3890
rect 400324 3806 400352 3862
rect 400312 3800 400364 3806
rect 400312 3742 400364 3748
rect 400128 3732 400180 3738
rect 400128 3674 400180 3680
rect 398932 3528 398984 3534
rect 398932 3470 398984 3476
rect 398944 480 398972 3470
rect 400140 480 400168 3674
rect 401520 3602 401548 29106
rect 401612 29034 401640 32028
rect 402716 29152 402744 32028
rect 403728 29170 403756 32028
rect 404740 29170 404768 32028
rect 403716 29164 403768 29170
rect 402716 29124 402928 29152
rect 401600 29028 401652 29034
rect 401600 28970 401652 28976
rect 402796 29028 402848 29034
rect 402796 28970 402848 28976
rect 401508 3596 401560 3602
rect 401508 3538 401560 3544
rect 402808 3534 402836 28970
rect 402900 3874 402928 29124
rect 403716 29106 403768 29112
rect 404268 29164 404320 29170
rect 404268 29106 404320 29112
rect 404728 29164 404780 29170
rect 404728 29106 404780 29112
rect 405648 29164 405700 29170
rect 405648 29106 405700 29112
rect 404280 4010 404308 29106
rect 403624 4004 403676 4010
rect 403624 3946 403676 3952
rect 404268 4004 404320 4010
rect 404268 3946 404320 3952
rect 402888 3868 402940 3874
rect 402888 3810 402940 3816
rect 402796 3528 402848 3534
rect 402796 3470 402848 3476
rect 401324 3392 401376 3398
rect 401324 3334 401376 3340
rect 401336 480 401364 3334
rect 402520 3324 402572 3330
rect 402520 3266 402572 3272
rect 402532 480 402560 3266
rect 403636 480 403664 3946
rect 404820 3664 404872 3670
rect 404820 3606 404872 3612
rect 404832 480 404860 3606
rect 405660 3262 405688 29106
rect 405844 29102 405872 32028
rect 406856 29186 406884 32028
rect 406856 29158 407068 29186
rect 407960 29170 407988 32028
rect 408972 29170 409000 32028
rect 410076 29170 410104 32028
rect 405832 29096 405884 29102
rect 405832 29038 405884 29044
rect 406936 29096 406988 29102
rect 406936 29038 406988 29044
rect 406016 4072 406068 4078
rect 406016 4014 406068 4020
rect 405648 3256 405700 3262
rect 405648 3198 405700 3204
rect 406028 480 406056 4014
rect 406948 3330 406976 29038
rect 407040 3670 407068 29158
rect 407948 29164 408000 29170
rect 407948 29106 408000 29112
rect 408408 29164 408460 29170
rect 408408 29106 408460 29112
rect 408960 29164 409012 29170
rect 408960 29106 409012 29112
rect 409788 29164 409840 29170
rect 409788 29106 409840 29112
rect 410064 29164 410116 29170
rect 410064 29106 410116 29112
rect 408420 6914 408448 29106
rect 408328 6886 408448 6914
rect 407028 3664 407080 3670
rect 407028 3606 407080 3612
rect 407212 3460 407264 3466
rect 407212 3402 407264 3408
rect 406936 3324 406988 3330
rect 406936 3266 406988 3272
rect 407224 480 407252 3402
rect 408328 3398 408356 6886
rect 408408 4140 408460 4146
rect 408408 4082 408460 4088
rect 408316 3392 408368 3398
rect 408316 3334 408368 3340
rect 408420 480 408448 4082
rect 409800 3738 409828 29106
rect 410800 3936 410852 3942
rect 410800 3878 410852 3884
rect 409604 3732 409656 3738
rect 409604 3674 409656 3680
rect 409788 3732 409840 3738
rect 409788 3674 409840 3680
rect 409616 480 409644 3674
rect 410812 480 410840 3878
rect 411088 3466 411116 32028
rect 411168 29164 411220 29170
rect 411168 29106 411220 29112
rect 411180 4078 411208 29106
rect 412192 26234 412220 32028
rect 413204 29102 413232 32028
rect 414308 29170 414336 32028
rect 414296 29164 414348 29170
rect 414296 29106 414348 29112
rect 415124 29164 415176 29170
rect 415124 29106 415176 29112
rect 413192 29096 413244 29102
rect 413192 29038 413244 29044
rect 413928 29096 413980 29102
rect 413928 29038 413980 29044
rect 412192 26206 412588 26234
rect 411168 4072 411220 4078
rect 411168 4014 411220 4020
rect 412560 3806 412588 26206
rect 413940 4146 413968 29038
rect 413928 4140 413980 4146
rect 413928 4082 413980 4088
rect 411904 3800 411956 3806
rect 411904 3742 411956 3748
rect 412548 3800 412600 3806
rect 412548 3742 412600 3748
rect 411076 3460 411128 3466
rect 411076 3402 411128 3408
rect 411916 480 411944 3742
rect 413100 3596 413152 3602
rect 413100 3538 413152 3544
rect 413112 480 413140 3538
rect 415136 3534 415164 29106
rect 415320 26234 415348 32028
rect 415228 26206 415348 26234
rect 416424 26234 416452 32028
rect 417436 29170 417464 32028
rect 418540 29170 418568 32028
rect 419552 29170 419580 32028
rect 417424 29164 417476 29170
rect 417424 29106 417476 29112
rect 418068 29164 418120 29170
rect 418068 29106 418120 29112
rect 418528 29164 418580 29170
rect 418528 29106 418580 29112
rect 419448 29164 419500 29170
rect 419448 29106 419500 29112
rect 419540 29164 419592 29170
rect 419540 29106 419592 29112
rect 416424 26206 416728 26234
rect 415228 3602 415256 26206
rect 416700 6914 416728 26206
rect 416608 6886 416728 6914
rect 416608 3942 416636 6886
rect 418080 4010 418108 29106
rect 416688 4004 416740 4010
rect 416688 3946 416740 3952
rect 418068 4004 418120 4010
rect 418068 3946 418120 3952
rect 416596 3936 416648 3942
rect 416596 3878 416648 3884
rect 415492 3868 415544 3874
rect 415492 3810 415544 3816
rect 415216 3596 415268 3602
rect 415216 3538 415268 3544
rect 414296 3528 414348 3534
rect 414296 3470 414348 3476
rect 415124 3528 415176 3534
rect 415124 3470 415176 3476
rect 414308 480 414336 3470
rect 415504 480 415532 3810
rect 416700 480 416728 3946
rect 418988 3324 419040 3330
rect 418988 3266 419040 3272
rect 417884 3256 417936 3262
rect 417884 3198 417936 3204
rect 417896 480 417924 3198
rect 419000 480 419028 3266
rect 419460 3194 419488 29106
rect 420564 26234 420592 32028
rect 421668 29170 421696 32028
rect 422680 29170 422708 32028
rect 423784 29170 423812 32028
rect 420828 29164 420880 29170
rect 420828 29106 420880 29112
rect 421656 29164 421708 29170
rect 421656 29106 421708 29112
rect 422208 29164 422260 29170
rect 422208 29106 422260 29112
rect 422668 29164 422720 29170
rect 422668 29106 422720 29112
rect 423588 29164 423640 29170
rect 423588 29106 423640 29112
rect 423772 29164 423824 29170
rect 423772 29106 423824 29112
rect 420564 26206 420776 26234
rect 420748 3670 420776 26206
rect 420184 3664 420236 3670
rect 420184 3606 420236 3612
rect 420736 3664 420788 3670
rect 420736 3606 420788 3612
rect 419448 3188 419500 3194
rect 419448 3130 419500 3136
rect 420196 480 420224 3606
rect 420840 3262 420868 29106
rect 422220 3874 422248 29106
rect 422208 3868 422260 3874
rect 422208 3810 422260 3816
rect 423600 3738 423628 29106
rect 424796 26234 424824 32028
rect 425900 29170 425928 32028
rect 426912 29170 426940 32028
rect 428016 29170 428044 32028
rect 424968 29164 425020 29170
rect 424968 29106 425020 29112
rect 425888 29164 425940 29170
rect 425888 29106 425940 29112
rect 426348 29164 426400 29170
rect 426348 29106 426400 29112
rect 426900 29164 426952 29170
rect 426900 29106 426952 29112
rect 427728 29164 427780 29170
rect 427728 29106 427780 29112
rect 428004 29164 428056 29170
rect 428004 29106 428056 29112
rect 428924 29164 428976 29170
rect 428924 29106 428976 29112
rect 424796 26206 424916 26234
rect 423772 4072 423824 4078
rect 423772 4014 423824 4020
rect 422576 3732 422628 3738
rect 422576 3674 422628 3680
rect 423588 3732 423640 3738
rect 423588 3674 423640 3680
rect 421380 3392 421432 3398
rect 421380 3334 421432 3340
rect 420828 3256 420880 3262
rect 420828 3198 420880 3204
rect 421392 480 421420 3334
rect 422588 480 422616 3674
rect 423784 480 423812 4014
rect 424888 3398 424916 26206
rect 424980 4078 425008 29106
rect 424968 4072 425020 4078
rect 424968 4014 425020 4020
rect 426164 3800 426216 3806
rect 426164 3742 426216 3748
rect 424968 3460 425020 3466
rect 424968 3402 425020 3408
rect 424876 3392 424928 3398
rect 424876 3334 424928 3340
rect 424980 480 425008 3402
rect 426176 480 426204 3742
rect 426360 3330 426388 29106
rect 427268 4140 427320 4146
rect 427268 4082 427320 4088
rect 426348 3324 426400 3330
rect 426348 3266 426400 3272
rect 427280 480 427308 4082
rect 427740 3126 427768 29106
rect 428936 3806 428964 29106
rect 429028 26234 429056 32028
rect 430132 26234 430160 32028
rect 431144 29102 431172 32028
rect 432248 29102 432276 32028
rect 431132 29096 431184 29102
rect 431132 29038 431184 29044
rect 431868 29096 431920 29102
rect 431868 29038 431920 29044
rect 432236 29096 432288 29102
rect 432236 29038 432288 29044
rect 433064 29096 433116 29102
rect 433064 29038 433116 29044
rect 429028 26206 429148 26234
rect 430132 26206 430528 26234
rect 428924 3800 428976 3806
rect 428924 3742 428976 3748
rect 429120 3534 429148 26206
rect 430500 4146 430528 26206
rect 430488 4140 430540 4146
rect 430488 4082 430540 4088
rect 430856 3936 430908 3942
rect 430856 3878 430908 3884
rect 429660 3596 429712 3602
rect 429660 3538 429712 3544
rect 428464 3528 428516 3534
rect 428464 3470 428516 3476
rect 429108 3528 429160 3534
rect 429108 3470 429160 3476
rect 427728 3120 427780 3126
rect 427728 3062 427780 3068
rect 428476 480 428504 3470
rect 429672 480 429700 3538
rect 430868 480 430896 3878
rect 431880 3058 431908 29038
rect 433076 4010 433104 29038
rect 433260 26234 433288 32028
rect 433168 26206 433288 26234
rect 434272 26234 434300 32028
rect 435376 29170 435404 32028
rect 436388 29170 436416 32028
rect 437492 29170 437520 32028
rect 435364 29164 435416 29170
rect 435364 29106 435416 29112
rect 436008 29164 436060 29170
rect 436008 29106 436060 29112
rect 436376 29164 436428 29170
rect 436376 29106 436428 29112
rect 437388 29164 437440 29170
rect 437388 29106 437440 29112
rect 437480 29164 437532 29170
rect 437480 29106 437532 29112
rect 434272 26206 434668 26234
rect 432052 4004 432104 4010
rect 432052 3946 432104 3952
rect 433064 4004 433116 4010
rect 433064 3946 433116 3952
rect 431868 3052 431920 3058
rect 431868 2994 431920 3000
rect 432064 480 432092 3946
rect 433168 3602 433196 26206
rect 433156 3596 433208 3602
rect 433156 3538 433208 3544
rect 434640 3466 434668 26206
rect 436020 3942 436048 29106
rect 436008 3936 436060 3942
rect 436008 3878 436060 3884
rect 437400 3874 437428 29106
rect 438504 26234 438532 32028
rect 439608 29170 439636 32028
rect 440620 29170 440648 32028
rect 441724 29170 441752 32028
rect 438768 29164 438820 29170
rect 438768 29106 438820 29112
rect 439596 29164 439648 29170
rect 439596 29106 439648 29112
rect 440148 29164 440200 29170
rect 440148 29106 440200 29112
rect 440608 29164 440660 29170
rect 440608 29106 440660 29112
rect 441528 29164 441580 29170
rect 441528 29106 441580 29112
rect 441712 29164 441764 29170
rect 441712 29106 441764 29112
rect 438504 26206 438716 26234
rect 436744 3868 436796 3874
rect 436744 3810 436796 3816
rect 437388 3868 437440 3874
rect 437388 3810 437440 3816
rect 435548 3664 435600 3670
rect 435548 3606 435600 3612
rect 434628 3460 434680 3466
rect 434628 3402 434680 3408
rect 434444 3256 434496 3262
rect 434444 3198 434496 3204
rect 433248 3188 433300 3194
rect 433248 3130 433300 3136
rect 433260 480 433288 3130
rect 434456 480 434484 3198
rect 435560 480 435588 3606
rect 436756 480 436784 3810
rect 437940 3732 437992 3738
rect 437940 3674 437992 3680
rect 437952 480 437980 3674
rect 438688 3670 438716 26206
rect 438676 3664 438728 3670
rect 438676 3606 438728 3612
rect 438780 3194 438808 29106
rect 440160 4078 440188 29106
rect 441540 6914 441568 29106
rect 442736 26234 442764 32028
rect 443840 29170 443868 32028
rect 444852 29170 444880 32028
rect 445956 29170 445984 32028
rect 442908 29164 442960 29170
rect 442908 29106 442960 29112
rect 443828 29164 443880 29170
rect 443828 29106 443880 29112
rect 444288 29164 444340 29170
rect 444288 29106 444340 29112
rect 444840 29164 444892 29170
rect 444840 29106 444892 29112
rect 445668 29164 445720 29170
rect 445668 29106 445720 29112
rect 445944 29164 445996 29170
rect 445944 29106 445996 29112
rect 446864 29164 446916 29170
rect 446864 29106 446916 29112
rect 442736 26206 442856 26234
rect 441448 6886 441568 6914
rect 439136 4072 439188 4078
rect 439136 4014 439188 4020
rect 440148 4072 440200 4078
rect 440148 4014 440200 4020
rect 438768 3188 438820 3194
rect 438768 3130 438820 3136
rect 439148 480 439176 4014
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 440344 480 440372 3334
rect 441448 3262 441476 6886
rect 442828 3738 442856 26206
rect 442816 3732 442868 3738
rect 442816 3674 442868 3680
rect 441528 3324 441580 3330
rect 441528 3266 441580 3272
rect 441436 3256 441488 3262
rect 441436 3198 441488 3204
rect 441540 480 441568 3266
rect 442920 3126 442948 29106
rect 444300 3806 444328 29106
rect 443828 3800 443880 3806
rect 443828 3742 443880 3748
rect 444288 3800 444340 3806
rect 444288 3742 444340 3748
rect 442632 3120 442684 3126
rect 442632 3062 442684 3068
rect 442908 3120 442960 3126
rect 442908 3062 442960 3068
rect 442644 480 442672 3062
rect 443840 480 443868 3742
rect 445024 3528 445076 3534
rect 445024 3470 445076 3476
rect 445036 480 445064 3470
rect 445680 3330 445708 29106
rect 446220 4140 446272 4146
rect 446220 4082 446272 4088
rect 445668 3324 445720 3330
rect 445668 3266 445720 3272
rect 446232 480 446260 4082
rect 446876 3534 446904 29106
rect 446968 26234 446996 32028
rect 448072 26234 448100 32028
rect 449084 29170 449112 32028
rect 450096 29170 450124 32028
rect 449072 29164 449124 29170
rect 449072 29106 449124 29112
rect 449808 29164 449860 29170
rect 449808 29106 449860 29112
rect 450084 29164 450136 29170
rect 450084 29106 450136 29112
rect 451096 29164 451148 29170
rect 451096 29106 451148 29112
rect 446968 26206 447088 26234
rect 448072 26206 448468 26234
rect 446864 3528 446916 3534
rect 446864 3470 446916 3476
rect 447060 3466 447088 26206
rect 447048 3460 447100 3466
rect 447048 3402 447100 3408
rect 448440 3058 448468 26206
rect 449820 6914 449848 29106
rect 449728 6886 449848 6914
rect 448612 4004 448664 4010
rect 448612 3946 448664 3952
rect 447416 3052 447468 3058
rect 447416 2994 447468 3000
rect 448428 3052 448480 3058
rect 448428 2994 448480 3000
rect 447428 480 447456 2994
rect 448624 480 448652 3946
rect 449728 2854 449756 6886
rect 451108 3602 451136 29106
rect 451200 4010 451228 32028
rect 452212 26234 452240 32028
rect 453316 29170 453344 32028
rect 454328 29170 454356 32028
rect 455432 29170 455460 32028
rect 453304 29164 453356 29170
rect 453304 29106 453356 29112
rect 453948 29164 454000 29170
rect 453948 29106 454000 29112
rect 454316 29164 454368 29170
rect 454316 29106 454368 29112
rect 455328 29164 455380 29170
rect 455328 29106 455380 29112
rect 455420 29164 455472 29170
rect 455420 29106 455472 29112
rect 452212 26206 452608 26234
rect 451188 4004 451240 4010
rect 451188 3946 451240 3952
rect 452580 3942 452608 26206
rect 452108 3936 452160 3942
rect 452108 3878 452160 3884
rect 452568 3936 452620 3942
rect 452568 3878 452620 3884
rect 449808 3596 449860 3602
rect 449808 3538 449860 3544
rect 451096 3596 451148 3602
rect 451096 3538 451148 3544
rect 449716 2848 449768 2854
rect 449716 2790 449768 2796
rect 449820 480 449848 3538
rect 450912 3392 450964 3398
rect 450912 3334 450964 3340
rect 450924 480 450952 3334
rect 452120 480 452148 3878
rect 453304 3868 453356 3874
rect 453304 3810 453356 3816
rect 453316 480 453344 3810
rect 453960 3398 453988 29106
rect 455340 4146 455368 29106
rect 456444 26234 456472 32028
rect 457548 29170 457576 32028
rect 458560 29170 458588 32028
rect 456708 29164 456760 29170
rect 456708 29106 456760 29112
rect 457536 29164 457588 29170
rect 457536 29106 457588 29112
rect 458088 29164 458140 29170
rect 458088 29106 458140 29112
rect 458548 29164 458600 29170
rect 458548 29106 458600 29112
rect 459468 29164 459520 29170
rect 459468 29106 459520 29112
rect 456444 26206 456656 26234
rect 455328 4140 455380 4146
rect 455328 4082 455380 4088
rect 456628 3874 456656 26206
rect 456616 3868 456668 3874
rect 456616 3810 456668 3816
rect 455696 3664 455748 3670
rect 455696 3606 455748 3612
rect 453948 3392 454000 3398
rect 453948 3334 454000 3340
rect 454500 3188 454552 3194
rect 454500 3130 454552 3136
rect 454512 480 454540 3130
rect 455708 480 455736 3606
rect 456720 2922 456748 29106
rect 458100 6914 458128 29106
rect 458008 6886 458128 6914
rect 456892 4072 456944 4078
rect 456892 4014 456944 4020
rect 456708 2916 456760 2922
rect 456708 2858 456760 2864
rect 456904 480 456932 4014
rect 458008 3194 458036 6886
rect 458088 3256 458140 3262
rect 458088 3198 458140 3204
rect 457996 3188 458048 3194
rect 457996 3130 458048 3136
rect 458100 480 458128 3198
rect 459480 3126 459508 29106
rect 459664 29034 459692 32028
rect 460676 29152 460704 32028
rect 461780 29170 461808 32028
rect 462792 29170 462820 32028
rect 463804 29170 463832 32028
rect 461768 29164 461820 29170
rect 460676 29124 460888 29152
rect 459652 29028 459704 29034
rect 459652 28970 459704 28976
rect 460756 29028 460808 29034
rect 460756 28970 460808 28976
rect 460768 4078 460796 28970
rect 460756 4072 460808 4078
rect 460756 4014 460808 4020
rect 460388 3732 460440 3738
rect 460388 3674 460440 3680
rect 459192 3120 459244 3126
rect 459192 3062 459244 3068
rect 459468 3120 459520 3126
rect 459468 3062 459520 3068
rect 459204 480 459232 3062
rect 460400 480 460428 3674
rect 460860 3670 460888 29124
rect 461768 29106 461820 29112
rect 462228 29164 462280 29170
rect 462228 29106 462280 29112
rect 462780 29164 462832 29170
rect 462780 29106 462832 29112
rect 463608 29164 463660 29170
rect 463608 29106 463660 29112
rect 463792 29164 463844 29170
rect 463792 29106 463844 29112
rect 462240 3806 462268 29106
rect 461584 3800 461636 3806
rect 461584 3742 461636 3748
rect 462228 3800 462280 3806
rect 462228 3742 462280 3748
rect 460848 3664 460900 3670
rect 460848 3606 460900 3612
rect 461596 480 461624 3742
rect 462780 3324 462832 3330
rect 462780 3266 462832 3272
rect 462792 480 462820 3266
rect 463620 2990 463648 29106
rect 464908 3534 464936 32028
rect 465920 29170 465948 32028
rect 467024 29170 467052 32028
rect 468036 29170 468064 32028
rect 464988 29164 465040 29170
rect 464988 29106 465040 29112
rect 465908 29164 465960 29170
rect 465908 29106 465960 29112
rect 466368 29164 466420 29170
rect 466368 29106 466420 29112
rect 467012 29164 467064 29170
rect 467012 29106 467064 29112
rect 467748 29164 467800 29170
rect 467748 29106 467800 29112
rect 468024 29164 468076 29170
rect 468024 29106 468076 29112
rect 469036 29164 469088 29170
rect 469036 29106 469088 29112
rect 463976 3528 464028 3534
rect 463976 3470 464028 3476
rect 464896 3528 464948 3534
rect 464896 3470 464948 3476
rect 463608 2984 463660 2990
rect 463608 2926 463660 2932
rect 463988 480 464016 3470
rect 465000 3262 465028 29106
rect 466380 3738 466408 29106
rect 467760 4962 467788 29106
rect 467748 4956 467800 4962
rect 467748 4898 467800 4904
rect 466368 3732 466420 3738
rect 466368 3674 466420 3680
rect 469048 3602 469076 29106
rect 468668 3596 468720 3602
rect 468668 3538 468720 3544
rect 469036 3596 469088 3602
rect 469036 3538 469088 3544
rect 465172 3460 465224 3466
rect 465172 3402 465224 3408
rect 464988 3256 465040 3262
rect 464988 3198 465040 3204
rect 465184 480 465212 3402
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467472 2848 467524 2854
rect 467472 2790 467524 2796
rect 467484 480 467512 2790
rect 468680 480 468708 3538
rect 469140 3466 469168 32028
rect 470152 30258 470180 32028
rect 470140 30252 470192 30258
rect 470140 30194 470192 30200
rect 471256 29170 471284 32028
rect 471336 30252 471388 30258
rect 471336 30194 471388 30200
rect 471244 29164 471296 29170
rect 471244 29106 471296 29112
rect 471348 5166 471376 30194
rect 472268 29170 472296 32028
rect 473372 29170 473400 32028
rect 471888 29164 471940 29170
rect 471888 29106 471940 29112
rect 472256 29164 472308 29170
rect 472256 29106 472308 29112
rect 473268 29164 473320 29170
rect 473268 29106 473320 29112
rect 473360 29164 473412 29170
rect 473360 29106 473412 29112
rect 471336 5160 471388 5166
rect 471336 5102 471388 5108
rect 469864 4004 469916 4010
rect 469864 3946 469916 3952
rect 469128 3460 469180 3466
rect 469128 3402 469180 3408
rect 469876 480 469904 3946
rect 471060 3936 471112 3942
rect 471060 3878 471112 3884
rect 471072 480 471100 3878
rect 471900 3058 471928 29106
rect 472256 3392 472308 3398
rect 472256 3334 472308 3340
rect 471888 3052 471940 3058
rect 471888 2994 471940 3000
rect 472268 480 472296 3334
rect 473280 3330 473308 29106
rect 474384 26234 474412 32028
rect 475488 29170 475516 32028
rect 476500 29170 476528 32028
rect 477604 29170 477632 32028
rect 475384 29164 475436 29170
rect 475384 29106 475436 29112
rect 475476 29164 475528 29170
rect 475476 29106 475528 29112
rect 476028 29164 476080 29170
rect 476028 29106 476080 29112
rect 476488 29164 476540 29170
rect 476488 29106 476540 29112
rect 477408 29164 477460 29170
rect 477408 29106 477460 29112
rect 477592 29164 477644 29170
rect 477592 29106 477644 29112
rect 474384 26206 474688 26234
rect 473452 4140 473504 4146
rect 473452 4082 473504 4088
rect 473268 3324 473320 3330
rect 473268 3266 473320 3272
rect 473464 480 473492 4082
rect 474660 3398 474688 26206
rect 475396 5302 475424 29106
rect 475384 5296 475436 5302
rect 475384 5238 475436 5244
rect 476040 4010 476068 29106
rect 477420 5098 477448 29106
rect 478616 26234 478644 32028
rect 479628 29170 479656 32028
rect 480732 29170 480760 32028
rect 481744 29170 481772 32028
rect 478788 29164 478840 29170
rect 478788 29106 478840 29112
rect 479616 29164 479668 29170
rect 479616 29106 479668 29112
rect 480168 29164 480220 29170
rect 480168 29106 480220 29112
rect 480720 29164 480772 29170
rect 480720 29106 480772 29112
rect 481548 29164 481600 29170
rect 481548 29106 481600 29112
rect 481732 29164 481784 29170
rect 481732 29106 481784 29112
rect 478616 26206 478736 26234
rect 477408 5092 477460 5098
rect 477408 5034 477460 5040
rect 476028 4004 476080 4010
rect 476028 3946 476080 3952
rect 478708 3942 478736 26206
rect 478696 3936 478748 3942
rect 478696 3878 478748 3884
rect 475752 3868 475804 3874
rect 475752 3810 475804 3816
rect 474648 3392 474700 3398
rect 474648 3334 474700 3340
rect 474556 2916 474608 2922
rect 474556 2858 474608 2864
rect 474568 480 474596 2858
rect 475764 480 475792 3810
rect 476948 3188 477000 3194
rect 476948 3130 477000 3136
rect 476960 480 476988 3130
rect 478800 3126 478828 29106
rect 480180 4826 480208 29106
rect 480168 4820 480220 4826
rect 480168 4762 480220 4768
rect 481560 4146 481588 29106
rect 482848 4894 482876 32028
rect 483860 29170 483888 32028
rect 484964 29170 484992 32028
rect 485976 29170 486004 32028
rect 482928 29164 482980 29170
rect 482928 29106 482980 29112
rect 483848 29164 483900 29170
rect 483848 29106 483900 29112
rect 484308 29164 484360 29170
rect 484308 29106 484360 29112
rect 484952 29164 485004 29170
rect 484952 29106 485004 29112
rect 485688 29164 485740 29170
rect 485688 29106 485740 29112
rect 485964 29164 486016 29170
rect 485964 29106 486016 29112
rect 486976 29164 487028 29170
rect 486976 29106 487028 29112
rect 482836 4888 482888 4894
rect 482836 4830 482888 4836
rect 481548 4140 481600 4146
rect 481548 4082 481600 4088
rect 479340 4072 479392 4078
rect 479340 4014 479392 4020
rect 478144 3120 478196 3126
rect 478144 3062 478196 3068
rect 478788 3120 478840 3126
rect 478788 3062 478840 3068
rect 478156 480 478184 3062
rect 479352 480 479380 4014
rect 481732 3800 481784 3806
rect 481732 3742 481784 3748
rect 480536 3664 480588 3670
rect 480536 3606 480588 3612
rect 480548 480 480576 3606
rect 481744 480 481772 3742
rect 482940 3194 482968 29106
rect 484320 3670 484348 29106
rect 484308 3664 484360 3670
rect 484308 3606 484360 3612
rect 485228 3528 485280 3534
rect 485228 3470 485280 3476
rect 484032 3256 484084 3262
rect 484032 3198 484084 3204
rect 482928 3188 482980 3194
rect 482928 3130 482980 3136
rect 482836 2984 482888 2990
rect 482836 2926 482888 2932
rect 482848 480 482876 2926
rect 484044 480 484072 3198
rect 485240 480 485268 3470
rect 485700 3262 485728 29106
rect 486988 5030 487016 29106
rect 486976 5024 487028 5030
rect 486976 4966 487028 4972
rect 487080 4078 487108 32028
rect 488092 26234 488120 32028
rect 489196 29170 489224 32028
rect 490208 29170 490236 32028
rect 491312 29170 491340 32028
rect 489184 29164 489236 29170
rect 489184 29106 489236 29112
rect 489828 29164 489880 29170
rect 489828 29106 489880 29112
rect 490196 29164 490248 29170
rect 490196 29106 490248 29112
rect 491208 29164 491260 29170
rect 491208 29106 491260 29112
rect 491300 29164 491352 29170
rect 491300 29106 491352 29112
rect 488092 26206 488488 26234
rect 487620 4956 487672 4962
rect 487620 4898 487672 4904
rect 487068 4072 487120 4078
rect 487068 4014 487120 4020
rect 486424 3732 486476 3738
rect 486424 3674 486476 3680
rect 485688 3256 485740 3262
rect 485688 3198 485740 3204
rect 486436 480 486464 3674
rect 487632 480 487660 4898
rect 488460 3738 488488 26206
rect 489840 4962 489868 29106
rect 491116 5160 491168 5166
rect 491116 5102 491168 5108
rect 489828 4956 489880 4962
rect 489828 4898 489880 4904
rect 488448 3732 488500 3738
rect 488448 3674 488500 3680
rect 488816 3596 488868 3602
rect 488816 3538 488868 3544
rect 488828 480 488856 3538
rect 489920 3460 489972 3466
rect 489920 3402 489972 3408
rect 489932 480 489960 3402
rect 491128 480 491156 5102
rect 491220 3874 491248 29106
rect 492324 29102 492352 32028
rect 493336 29170 493364 32028
rect 494440 29170 494468 32028
rect 495452 29170 495480 32028
rect 492588 29164 492640 29170
rect 492588 29106 492640 29112
rect 493324 29164 493376 29170
rect 493324 29106 493376 29112
rect 493968 29164 494020 29170
rect 493968 29106 494020 29112
rect 494428 29164 494480 29170
rect 494428 29106 494480 29112
rect 495348 29164 495400 29170
rect 495348 29106 495400 29112
rect 495440 29164 495492 29170
rect 495440 29106 495492 29112
rect 492312 29096 492364 29102
rect 492312 29038 492364 29044
rect 491208 3868 491260 3874
rect 491208 3810 491260 3816
rect 492600 3806 492628 29106
rect 493416 29096 493468 29102
rect 493416 29038 493468 29044
rect 493428 5234 493456 29038
rect 493416 5228 493468 5234
rect 493416 5170 493468 5176
rect 492588 3800 492640 3806
rect 492588 3742 492640 3748
rect 493980 3534 494008 29106
rect 494704 5296 494756 5302
rect 494704 5238 494756 5244
rect 493968 3528 494020 3534
rect 493968 3470 494020 3476
rect 493508 3324 493560 3330
rect 493508 3266 493560 3272
rect 492312 3052 492364 3058
rect 492312 2994 492364 3000
rect 492324 480 492352 2994
rect 493520 480 493548 3266
rect 494716 480 494744 5238
rect 495360 3602 495388 29106
rect 496556 26234 496584 32028
rect 497568 29170 497596 32028
rect 498672 29646 498700 32028
rect 498660 29640 498712 29646
rect 498660 29582 498712 29588
rect 499684 29170 499712 32028
rect 497464 29164 497516 29170
rect 497464 29106 497516 29112
rect 497556 29164 497608 29170
rect 497556 29106 497608 29112
rect 498108 29164 498160 29170
rect 498108 29106 498160 29112
rect 499672 29164 499724 29170
rect 499672 29106 499724 29112
rect 500684 29164 500736 29170
rect 500684 29106 500736 29112
rect 496556 26206 496768 26234
rect 495348 3596 495400 3602
rect 495348 3538 495400 3544
rect 496740 3398 496768 26206
rect 497476 5166 497504 29106
rect 497464 5160 497516 5166
rect 497464 5102 497516 5108
rect 497096 4004 497148 4010
rect 497096 3946 497148 3952
rect 495900 3392 495952 3398
rect 495900 3334 495952 3340
rect 496728 3392 496780 3398
rect 496728 3334 496780 3340
rect 495912 480 495940 3334
rect 497108 480 497136 3946
rect 498120 3466 498148 29106
rect 498200 5092 498252 5098
rect 498200 5034 498252 5040
rect 498108 3460 498160 3466
rect 498108 3402 498160 3408
rect 498212 480 498240 5034
rect 500592 3936 500644 3942
rect 500592 3878 500644 3884
rect 499396 3120 499448 3126
rect 499396 3062 499448 3068
rect 499408 480 499436 3062
rect 500604 480 500632 3878
rect 500696 3126 500724 29106
rect 500788 26234 500816 32028
rect 501800 29170 501828 32028
rect 502904 29170 502932 32028
rect 503916 29170 503944 32028
rect 501788 29164 501840 29170
rect 501788 29106 501840 29112
rect 502248 29164 502300 29170
rect 502248 29106 502300 29112
rect 502892 29164 502944 29170
rect 502892 29106 502944 29112
rect 503628 29164 503680 29170
rect 503628 29106 503680 29112
rect 503904 29164 503956 29170
rect 503904 29106 503956 29112
rect 504824 29164 504876 29170
rect 504824 29106 504876 29112
rect 500788 26206 500908 26234
rect 500880 3330 500908 26206
rect 502260 5098 502288 29106
rect 502248 5092 502300 5098
rect 502248 5034 502300 5040
rect 501788 4820 501840 4826
rect 501788 4762 501840 4768
rect 500868 3324 500920 3330
rect 500868 3266 500920 3272
rect 500684 3120 500736 3126
rect 500684 3062 500736 3068
rect 501800 480 501828 4762
rect 503640 4146 503668 29106
rect 502984 4140 503036 4146
rect 502984 4082 503036 4088
rect 503628 4140 503680 4146
rect 503628 4082 503680 4088
rect 502996 480 503024 4082
rect 504836 3194 504864 29106
rect 505020 26234 505048 32028
rect 504928 26206 505048 26234
rect 506032 26234 506060 32028
rect 507136 29170 507164 32028
rect 508148 29714 508176 32028
rect 508136 29708 508188 29714
rect 508136 29650 508188 29656
rect 507124 29164 507176 29170
rect 507124 29106 507176 29112
rect 507768 29164 507820 29170
rect 507768 29106 507820 29112
rect 506032 26206 506428 26234
rect 504928 4826 504956 26206
rect 505376 4888 505428 4894
rect 505376 4830 505428 4836
rect 504916 4820 504968 4826
rect 504916 4762 504968 4768
rect 504180 3188 504232 3194
rect 504180 3130 504232 3136
rect 504824 3188 504876 3194
rect 504824 3130 504876 3136
rect 504192 480 504220 3130
rect 505388 480 505416 4830
rect 506400 4010 506428 26206
rect 506388 4004 506440 4010
rect 506388 3946 506440 3952
rect 506480 3664 506532 3670
rect 506480 3606 506532 3612
rect 506492 480 506520 3606
rect 507780 3262 507808 29106
rect 508872 5024 508924 5030
rect 508872 4966 508924 4972
rect 507676 3256 507728 3262
rect 507676 3198 507728 3204
rect 507768 3256 507820 3262
rect 507768 3198 507820 3204
rect 507688 480 507716 3198
rect 508884 480 508912 4966
rect 509160 3942 509188 32028
rect 510264 26234 510292 32028
rect 511276 29170 511304 32028
rect 511356 29708 511408 29714
rect 511356 29650 511408 29656
rect 511264 29164 511316 29170
rect 511264 29106 511316 29112
rect 510264 26206 510568 26234
rect 510068 4072 510120 4078
rect 510068 4014 510120 4020
rect 509148 3936 509200 3942
rect 509148 3878 509200 3884
rect 510080 480 510108 4014
rect 510540 3670 510568 26206
rect 511368 5302 511396 29650
rect 512380 29170 512408 32028
rect 513392 29170 513420 32028
rect 514496 29714 514524 32028
rect 514484 29708 514536 29714
rect 514484 29650 514536 29656
rect 515508 29170 515536 32028
rect 516612 29170 516640 32028
rect 517624 29170 517652 32028
rect 511908 29164 511960 29170
rect 511908 29106 511960 29112
rect 512368 29164 512420 29170
rect 512368 29106 512420 29112
rect 513288 29164 513340 29170
rect 513288 29106 513340 29112
rect 513380 29164 513432 29170
rect 513380 29106 513432 29112
rect 514668 29164 514720 29170
rect 514668 29106 514720 29112
rect 515496 29164 515548 29170
rect 515496 29106 515548 29112
rect 516048 29164 516100 29170
rect 516048 29106 516100 29112
rect 516600 29164 516652 29170
rect 516600 29106 516652 29112
rect 517428 29164 517480 29170
rect 517428 29106 517480 29112
rect 517612 29164 517664 29170
rect 517612 29106 517664 29112
rect 518624 29164 518676 29170
rect 518624 29106 518676 29112
rect 511356 5296 511408 5302
rect 511356 5238 511408 5244
rect 511920 5030 511948 29106
rect 511908 5024 511960 5030
rect 511908 4966 511960 4972
rect 512460 4956 512512 4962
rect 512460 4898 512512 4904
rect 511264 3732 511316 3738
rect 511264 3674 511316 3680
rect 510528 3664 510580 3670
rect 510528 3606 510580 3612
rect 511276 480 511304 3674
rect 512472 480 512500 4898
rect 513300 4078 513328 29106
rect 513288 4072 513340 4078
rect 513288 4014 513340 4020
rect 513564 3868 513616 3874
rect 513564 3810 513616 3816
rect 513576 480 513604 3810
rect 514680 3738 514708 29106
rect 515956 5228 516008 5234
rect 515956 5170 516008 5176
rect 514760 3800 514812 3806
rect 514760 3742 514812 3748
rect 514668 3732 514720 3738
rect 514668 3674 514720 3680
rect 514772 480 514800 3742
rect 515968 480 515996 5170
rect 516060 3806 516088 29106
rect 517440 3874 517468 29106
rect 518636 4962 518664 29106
rect 518728 26234 518756 32028
rect 519740 29170 519768 32028
rect 520844 29170 520872 32028
rect 520924 29640 520976 29646
rect 520924 29582 520976 29588
rect 519728 29164 519780 29170
rect 519728 29106 519780 29112
rect 520188 29164 520240 29170
rect 520188 29106 520240 29112
rect 520832 29164 520884 29170
rect 520832 29106 520884 29112
rect 518728 26206 518848 26234
rect 518624 4956 518676 4962
rect 518624 4898 518676 4904
rect 517428 3868 517480 3874
rect 517428 3810 517480 3816
rect 516048 3800 516100 3806
rect 516048 3742 516100 3748
rect 518820 3602 518848 26206
rect 519544 5160 519596 5166
rect 519544 5102 519596 5108
rect 518348 3596 518400 3602
rect 518348 3538 518400 3544
rect 518808 3596 518860 3602
rect 518808 3538 518860 3544
rect 517152 3528 517204 3534
rect 517152 3470 517204 3476
rect 517164 480 517192 3470
rect 518360 480 518388 3538
rect 519556 480 519584 5102
rect 520200 3534 520228 29106
rect 520936 4214 520964 29582
rect 521856 29170 521884 32028
rect 521568 29164 521620 29170
rect 521568 29106 521620 29112
rect 521844 29164 521896 29170
rect 521844 29106 521896 29112
rect 521580 4894 521608 29106
rect 521568 4888 521620 4894
rect 521568 4830 521620 4836
rect 520924 4208 520976 4214
rect 520924 4150 520976 4156
rect 520188 3528 520240 3534
rect 520188 3470 520240 3476
rect 522868 3466 522896 32028
rect 523972 29986 524000 32028
rect 523960 29980 524012 29986
rect 523960 29922 524012 29928
rect 524984 29170 525012 32028
rect 525064 29708 525116 29714
rect 525064 29650 525116 29656
rect 522948 29164 523000 29170
rect 522948 29106 523000 29112
rect 524972 29164 525024 29170
rect 524972 29106 525024 29112
rect 521844 3460 521896 3466
rect 521844 3402 521896 3408
rect 522856 3460 522908 3466
rect 522856 3402 522908 3408
rect 520740 3392 520792 3398
rect 520740 3334 520792 3340
rect 520752 480 520780 3334
rect 521856 480 521884 3402
rect 522960 2854 522988 29106
rect 525076 5166 525104 29650
rect 525708 29164 525760 29170
rect 525708 29106 525760 29112
rect 525064 5160 525116 5166
rect 525064 5102 525116 5108
rect 523040 4208 523092 4214
rect 523040 4150 523092 4156
rect 522948 2848 523000 2854
rect 522948 2790 523000 2796
rect 523052 480 523080 4150
rect 525432 3324 525484 3330
rect 525432 3266 525484 3272
rect 524236 3120 524288 3126
rect 524236 3062 524288 3068
rect 524248 480 524276 3062
rect 525444 480 525472 3266
rect 525720 3058 525748 29106
rect 526088 29102 526116 32028
rect 526076 29096 526128 29102
rect 526076 29038 526128 29044
rect 526904 29096 526956 29102
rect 526904 29038 526956 29044
rect 526628 5092 526680 5098
rect 526628 5034 526680 5040
rect 525708 3052 525760 3058
rect 525708 2994 525760 3000
rect 526640 480 526668 5034
rect 526916 2990 526944 29038
rect 527100 26234 527128 32028
rect 527008 26206 527128 26234
rect 528204 26234 528232 32028
rect 529216 29034 529244 32028
rect 529296 29980 529348 29986
rect 529296 29922 529348 29928
rect 529204 29028 529256 29034
rect 529204 28970 529256 28976
rect 528204 26206 528508 26234
rect 527008 6186 527036 26206
rect 526996 6180 527048 6186
rect 526996 6122 527048 6128
rect 527824 4140 527876 4146
rect 527824 4082 527876 4088
rect 526904 2984 526956 2990
rect 526904 2926 526956 2932
rect 527836 480 527864 4082
rect 528480 3330 528508 26206
rect 529308 5098 529336 29922
rect 530320 29850 530348 32028
rect 530308 29844 530360 29850
rect 530308 29786 530360 29792
rect 531332 29170 531360 32028
rect 531320 29164 531372 29170
rect 531320 29106 531372 29112
rect 529848 29028 529900 29034
rect 529848 28970 529900 28976
rect 529296 5092 529348 5098
rect 529296 5034 529348 5040
rect 528468 3324 528520 3330
rect 528468 3266 528520 3272
rect 529020 3188 529072 3194
rect 529020 3130 529072 3136
rect 529032 480 529060 3130
rect 529860 2922 529888 28970
rect 532436 26234 532464 32028
rect 533448 29170 533476 32028
rect 534552 29170 534580 32028
rect 535564 29170 535592 32028
rect 536668 29782 536696 32028
rect 536656 29776 536708 29782
rect 536656 29718 536708 29724
rect 537680 29170 537708 32028
rect 538692 29170 538720 32028
rect 539796 29714 539824 32028
rect 539784 29708 539836 29714
rect 539784 29650 539836 29656
rect 532608 29164 532660 29170
rect 532608 29106 532660 29112
rect 533436 29164 533488 29170
rect 533436 29106 533488 29112
rect 533988 29164 534040 29170
rect 533988 29106 534040 29112
rect 534540 29164 534592 29170
rect 534540 29106 534592 29112
rect 535368 29164 535420 29170
rect 535368 29106 535420 29112
rect 535552 29164 535604 29170
rect 535552 29106 535604 29112
rect 536748 29164 536800 29170
rect 536748 29106 536800 29112
rect 537668 29164 537720 29170
rect 537668 29106 537720 29112
rect 538128 29164 538180 29170
rect 538128 29106 538180 29112
rect 538680 29164 538732 29170
rect 538680 29106 538732 29112
rect 539508 29164 539560 29170
rect 539508 29106 539560 29112
rect 532436 26206 532556 26234
rect 530124 4820 530176 4826
rect 530124 4762 530176 4768
rect 529848 2916 529900 2922
rect 529848 2858 529900 2864
rect 530136 480 530164 4762
rect 532528 4010 532556 26206
rect 531320 4004 531372 4010
rect 531320 3946 531372 3952
rect 532516 4004 532568 4010
rect 532516 3946 532568 3952
rect 531332 480 531360 3946
rect 532516 3256 532568 3262
rect 532516 3198 532568 3204
rect 532528 480 532556 3198
rect 532620 3126 532648 29106
rect 533712 5296 533764 5302
rect 533712 5238 533764 5244
rect 532608 3120 532660 3126
rect 532608 3062 532660 3068
rect 533724 480 533752 5238
rect 534000 4826 534028 29106
rect 533988 4820 534040 4826
rect 533988 4762 534040 4768
rect 534908 3936 534960 3942
rect 534908 3878 534960 3884
rect 534920 480 534948 3878
rect 535380 3398 535408 29106
rect 536104 3664 536156 3670
rect 536104 3606 536156 3612
rect 535368 3392 535420 3398
rect 535368 3334 535420 3340
rect 536116 480 536144 3606
rect 536760 3194 536788 29106
rect 537208 5024 537260 5030
rect 537208 4966 537260 4972
rect 536748 3188 536800 3194
rect 536748 3130 536800 3136
rect 537220 480 537248 4966
rect 538140 4146 538168 29106
rect 538128 4140 538180 4146
rect 538128 4082 538180 4088
rect 538404 4072 538456 4078
rect 538404 4014 538456 4020
rect 538416 480 538444 4014
rect 539520 3262 539548 29106
rect 540808 26234 540836 32028
rect 541912 26234 541940 32028
rect 542924 29578 542952 32028
rect 542912 29572 542964 29578
rect 542912 29514 542964 29520
rect 544028 29170 544056 32028
rect 544016 29164 544068 29170
rect 544016 29106 544068 29112
rect 544936 29164 544988 29170
rect 544936 29106 544988 29112
rect 540808 26206 540928 26234
rect 541912 26206 542308 26234
rect 540796 5160 540848 5166
rect 540796 5102 540848 5108
rect 539600 3732 539652 3738
rect 539600 3674 539652 3680
rect 539508 3256 539560 3262
rect 539508 3198 539560 3204
rect 539612 480 539640 3674
rect 540808 480 540836 5102
rect 540900 3670 540928 26206
rect 542280 3942 542308 26206
rect 544384 4956 544436 4962
rect 544384 4898 544436 4904
rect 542268 3936 542320 3942
rect 542268 3878 542320 3884
rect 543188 3868 543240 3874
rect 543188 3810 543240 3816
rect 541992 3800 542044 3806
rect 541992 3742 542044 3748
rect 540888 3664 540940 3670
rect 540888 3606 540940 3612
rect 542004 480 542032 3742
rect 543200 480 543228 3810
rect 544396 480 544424 4898
rect 544948 4078 544976 29106
rect 544936 4072 544988 4078
rect 544936 4014 544988 4020
rect 545040 3874 545068 32028
rect 546144 29918 546172 32028
rect 546132 29912 546184 29918
rect 546132 29854 546184 29860
rect 547156 29102 547184 32028
rect 548260 29170 548288 32028
rect 548248 29164 548300 29170
rect 548248 29106 548300 29112
rect 549168 29164 549220 29170
rect 549168 29106 549220 29112
rect 547144 29096 547196 29102
rect 547144 29038 547196 29044
rect 547788 29096 547840 29102
rect 547788 29038 547840 29044
rect 545028 3868 545080 3874
rect 545028 3810 545080 3816
rect 547800 3738 547828 29038
rect 547880 4888 547932 4894
rect 547880 4830 547932 4836
rect 547788 3732 547840 3738
rect 547788 3674 547840 3680
rect 545488 3596 545540 3602
rect 545488 3538 545540 3544
rect 545500 480 545528 3538
rect 546684 3528 546736 3534
rect 546684 3470 546736 3476
rect 546696 480 546724 3470
rect 547892 480 547920 4830
rect 549180 3806 549208 29106
rect 549272 29102 549300 32028
rect 550376 29186 550404 32028
rect 551402 32014 551968 32042
rect 550376 29158 550588 29186
rect 549260 29096 549312 29102
rect 549260 29038 549312 29044
rect 550456 29096 550508 29102
rect 550456 29038 550508 29044
rect 549168 3800 549220 3806
rect 549168 3742 549220 3748
rect 550468 3466 550496 29038
rect 550560 3602 550588 29158
rect 551468 5092 551520 5098
rect 551468 5034 551520 5040
rect 550548 3596 550600 3602
rect 550548 3538 550600 3544
rect 550272 3460 550324 3466
rect 550272 3402 550324 3408
rect 550456 3460 550508 3466
rect 550456 3402 550508 3408
rect 549076 2848 549128 2854
rect 549076 2790 549128 2796
rect 549088 480 549116 2790
rect 550284 480 550312 3402
rect 551480 480 551508 5034
rect 551940 3534 551968 32014
rect 552676 20670 552704 674970
rect 552756 672988 552808 672994
rect 552756 672930 552808 672936
rect 552768 458182 552796 672930
rect 554042 670848 554098 670857
rect 554042 670783 554098 670792
rect 552846 669760 552902 669769
rect 552846 669695 552902 669704
rect 552860 538218 552888 669695
rect 552848 538212 552900 538218
rect 552848 538154 552900 538160
rect 552756 458176 552808 458182
rect 552756 458118 552808 458124
rect 554056 60722 554084 670783
rect 554148 485790 554176 675446
rect 558276 675436 558328 675442
rect 558276 675378 558328 675384
rect 555516 673804 555568 673810
rect 555516 673746 555568 673752
rect 554228 673124 554280 673130
rect 554228 673066 554280 673072
rect 554240 511970 554268 673066
rect 555422 672208 555478 672217
rect 555422 672143 555478 672152
rect 554228 511964 554280 511970
rect 554228 511906 554280 511912
rect 554136 485784 554188 485790
rect 554136 485726 554188 485732
rect 554044 60716 554096 60722
rect 554044 60658 554096 60664
rect 552664 20664 552716 20670
rect 552664 20606 552716 20612
rect 555436 6866 555464 672143
rect 555528 233238 555556 673746
rect 556988 673260 557040 673266
rect 556988 673202 557040 673208
rect 556896 672648 556948 672654
rect 556896 672590 556948 672596
rect 556802 670168 556858 670177
rect 556802 670103 556858 670112
rect 555516 233232 555568 233238
rect 555516 233174 555568 233180
rect 556816 33114 556844 670103
rect 556908 313274 556936 672590
rect 557000 564398 557028 673202
rect 557080 672036 557132 672042
rect 557080 671978 557132 671984
rect 557092 632058 557120 671978
rect 558184 670880 558236 670886
rect 558184 670822 558236 670828
rect 557080 632052 557132 632058
rect 557080 631994 557132 632000
rect 556988 564392 557040 564398
rect 556988 564334 557040 564340
rect 556896 313268 556948 313274
rect 556896 313210 556948 313216
rect 558196 113150 558224 670822
rect 558288 405686 558316 675378
rect 576216 675368 576268 675374
rect 576216 675310 576268 675316
rect 574836 675300 574888 675306
rect 574836 675242 574888 675248
rect 565084 675096 565136 675102
rect 565084 675038 565136 675044
rect 561036 673940 561088 673946
rect 561036 673882 561088 673888
rect 558368 673396 558420 673402
rect 558368 673338 558420 673344
rect 558380 618254 558408 673338
rect 560942 672344 560998 672353
rect 560942 672279 560998 672288
rect 558368 618248 558420 618254
rect 558368 618190 558420 618196
rect 558276 405680 558328 405686
rect 558276 405622 558328 405628
rect 558184 113144 558236 113150
rect 558184 113086 558236 113092
rect 560956 46918 560984 672279
rect 561048 273222 561076 673882
rect 562324 672172 562376 672178
rect 562324 672114 562376 672120
rect 561036 273216 561088 273222
rect 561036 273158 561088 273164
rect 562336 86970 562364 672114
rect 562416 671220 562468 671226
rect 562416 671162 562468 671168
rect 562428 325650 562456 671162
rect 562416 325644 562468 325650
rect 562416 325586 562468 325592
rect 565096 126954 565124 675038
rect 572076 674484 572128 674490
rect 572076 674426 572128 674432
rect 571984 674416 572036 674422
rect 571984 674358 572036 674364
rect 570604 674348 570656 674354
rect 570604 674290 570656 674296
rect 565176 674144 565228 674150
rect 565176 674086 565228 674092
rect 565188 379506 565216 674086
rect 569224 672240 569276 672246
rect 569224 672182 569276 672188
rect 566648 671628 566700 671634
rect 566648 671570 566700 671576
rect 566464 670744 566516 670750
rect 566464 670686 566516 670692
rect 565176 379500 565228 379506
rect 565176 379442 565228 379448
rect 565084 126948 565136 126954
rect 565084 126890 565136 126896
rect 566476 100706 566504 670686
rect 566554 670304 566610 670313
rect 566554 670239 566610 670248
rect 566568 167006 566596 670239
rect 566660 592006 566688 671570
rect 566648 592000 566700 592006
rect 566648 591942 566700 591948
rect 566556 167000 566608 167006
rect 566556 166942 566608 166948
rect 569236 139398 569264 672182
rect 569500 671832 569552 671838
rect 569500 671774 569552 671780
rect 569408 671696 569460 671702
rect 569408 671638 569460 671644
rect 569314 670440 569370 670449
rect 569314 670375 569370 670384
rect 569328 206990 569356 670375
rect 569420 578202 569448 671638
rect 569512 644434 569540 671774
rect 569500 644428 569552 644434
rect 569500 644370 569552 644376
rect 569408 578196 569460 578202
rect 569408 578138 569460 578144
rect 570616 431934 570644 674290
rect 570604 431928 570656 431934
rect 570604 431870 570656 431876
rect 571996 419490 572024 674358
rect 572088 471986 572116 674426
rect 573364 670948 573416 670954
rect 573364 670890 573416 670896
rect 572076 471980 572128 471986
rect 572076 471922 572128 471928
rect 571984 419484 572036 419490
rect 571984 419426 572036 419432
rect 569316 206984 569368 206990
rect 569316 206926 569368 206932
rect 573376 193186 573404 670890
rect 574744 670812 574796 670818
rect 574744 670754 574796 670760
rect 573454 670576 573510 670585
rect 573454 670511 573510 670520
rect 573468 245614 573496 670511
rect 573456 245608 573508 245614
rect 573456 245550 573508 245556
rect 573364 193180 573416 193186
rect 573364 193122 573416 193128
rect 574756 153202 574784 670754
rect 574848 299470 574876 675242
rect 576124 674892 576176 674898
rect 576124 674834 576176 674840
rect 574836 299464 574888 299470
rect 574836 299406 574888 299412
rect 574744 153196 574796 153202
rect 574744 153138 574796 153144
rect 569224 139392 569276 139398
rect 569224 139334 569276 139340
rect 566464 100700 566516 100706
rect 566464 100642 566516 100648
rect 562324 86964 562376 86970
rect 562324 86906 562376 86912
rect 576136 73166 576164 674834
rect 576228 353258 576256 675310
rect 579528 673328 579580 673334
rect 579528 673270 579580 673276
rect 578884 672308 578936 672314
rect 578884 672250 578936 672256
rect 576216 353252 576268 353258
rect 576216 353194 576268 353200
rect 578896 179217 578924 672250
rect 578976 671492 579028 671498
rect 578976 671434 579028 671440
rect 578988 524521 579016 671434
rect 579540 670721 579568 673270
rect 580264 672784 580316 672790
rect 580264 672726 580316 672732
rect 579526 670712 579582 670721
rect 579526 670647 579582 670656
rect 580172 644428 580224 644434
rect 580172 644370 580224 644376
rect 580184 644065 580212 644370
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 579712 632052 579764 632058
rect 579712 631994 579764 632000
rect 579724 630873 579752 631994
rect 579710 630864 579766 630873
rect 579710 630799 579766 630808
rect 579804 618248 579856 618254
rect 579804 618190 579856 618196
rect 579816 617545 579844 618190
rect 579802 617536 579858 617545
rect 579802 617471 579858 617480
rect 580172 592000 580224 592006
rect 580172 591942 580224 591948
rect 580184 591025 580212 591942
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580172 578196 580224 578202
rect 580172 578138 580224 578144
rect 580184 577697 580212 578138
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 578974 524512 579030 524521
rect 578974 524447 579030 524456
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 579712 419484 579764 419490
rect 579712 419426 579764 419432
rect 579724 418305 579752 419426
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 579804 405680 579856 405686
rect 579804 405622 579856 405628
rect 579816 404977 579844 405622
rect 579802 404968 579858 404977
rect 579802 404903 579858 404912
rect 579804 379500 579856 379506
rect 579804 379442 579856 379448
rect 579816 378457 579844 379442
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580276 219065 580304 672726
rect 580356 671968 580408 671974
rect 580356 671910 580408 671916
rect 580368 258913 580396 671910
rect 580448 671560 580500 671566
rect 580448 671502 580500 671508
rect 580460 365129 580488 671502
rect 580446 365120 580502 365129
rect 580446 365055 580502 365064
rect 580354 258904 580410 258913
rect 580354 258839 580410 258848
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 578882 179208 578938 179217
rect 578882 179143 578938 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 576124 73160 576176 73166
rect 576124 73102 576176 73108
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 560944 46912 560996 46918
rect 560944 46854 560996 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 556804 33108 556856 33114
rect 580170 33079 580172 33088
rect 556804 33050 556856 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 556804 29912 556856 29918
rect 556804 29854 556856 29860
rect 555424 6860 555476 6866
rect 555424 6802 555476 6808
rect 554964 6180 555016 6186
rect 554964 6122 555016 6128
rect 551928 3528 551980 3534
rect 551928 3470 551980 3476
rect 552664 3052 552716 3058
rect 552664 2994 552716 3000
rect 552676 480 552704 2994
rect 553768 2984 553820 2990
rect 553768 2926 553820 2932
rect 553780 480 553808 2926
rect 554976 480 555004 6122
rect 556816 4894 556844 29854
rect 557540 29844 557592 29850
rect 557540 29786 557592 29792
rect 557552 16574 557580 29786
rect 564532 29776 564584 29782
rect 564532 29718 564584 29724
rect 564544 16574 564572 29718
rect 568580 29708 568632 29714
rect 568580 29650 568632 29656
rect 568592 16574 568620 29650
rect 572812 29640 572864 29646
rect 572812 29582 572864 29588
rect 557552 16546 558592 16574
rect 564544 16546 565216 16574
rect 568592 16546 568712 16574
rect 556804 4888 556856 4894
rect 556804 4830 556856 4836
rect 556160 3324 556212 3330
rect 556160 3266 556212 3272
rect 556172 480 556200 3266
rect 557356 2916 557408 2922
rect 557356 2858 557408 2864
rect 557368 480 557396 2858
rect 558564 480 558592 16546
rect 562048 4820 562100 4826
rect 562048 4762 562100 4768
rect 560852 4004 560904 4010
rect 560852 3946 560904 3952
rect 559748 3120 559800 3126
rect 559748 3062 559800 3068
rect 559760 480 559788 3062
rect 560864 480 560892 3946
rect 562060 480 562088 4762
rect 563244 3392 563296 3398
rect 563244 3334 563296 3340
rect 563256 480 563284 3334
rect 564440 3188 564492 3194
rect 564440 3130 564492 3136
rect 564452 480 564480 3130
rect 565188 490 565216 16546
rect 566832 4140 566884 4146
rect 566832 4082 566884 4088
rect 565464 598 565676 626
rect 565464 490 565492 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 462 565492 490
rect 565648 480 565676 598
rect 566844 480 566872 4082
rect 568028 3256 568080 3262
rect 568028 3198 568080 3204
rect 568040 480 568068 3198
rect 568684 490 568712 16546
rect 572824 6914 572852 29582
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 572732 6886 572852 6914
rect 571524 3936 571576 3942
rect 571524 3878 571576 3884
rect 570328 3664 570380 3670
rect 570328 3606 570380 3612
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 3606
rect 571536 480 571564 3878
rect 572732 480 572760 6886
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 576308 4888 576360 4894
rect 576308 4830 576360 4836
rect 573916 4072 573968 4078
rect 573916 4014 573968 4020
rect 573928 480 573956 4014
rect 575112 3868 575164 3874
rect 575112 3810 575164 3816
rect 575124 480 575152 3810
rect 576320 480 576348 4830
rect 578608 3800 578660 3806
rect 578608 3742 578660 3748
rect 577412 3732 577464 3738
rect 577412 3674 577464 3680
rect 577424 480 577452 3674
rect 578620 480 578648 3742
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583392 3528 583444 3534
rect 583392 3470 583444 3476
rect 583404 480 583432 3470
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 4802 673784 4858 673840
rect 3330 671200 3386 671256
rect 3330 658180 3332 658200
rect 3332 658180 3384 658200
rect 3384 658180 3386 658200
rect 3330 658144 3386 658180
rect 3330 632032 3386 632088
rect 3330 619112 3386 619168
rect 3054 606056 3110 606112
rect 3330 579944 3386 580000
rect 3146 566888 3202 566944
rect 2962 553832 3018 553888
rect 3146 527856 3202 527912
rect 2962 501744 3018 501800
rect 3238 475632 3294 475688
rect 3054 462576 3110 462632
rect 3330 449520 3386 449576
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 2962 410488 3018 410544
rect 3330 397432 3386 397488
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 2962 267144 3018 267200
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 3606 514800 3662 514856
rect 3514 254088 3570 254144
rect 3514 241032 3570 241088
rect 3514 188808 3570 188864
rect 3422 149776 3478 149832
rect 3422 136720 3478 136776
rect 3146 110608 3202 110664
rect 3514 97552 3570 97608
rect 3146 84632 3202 84688
rect 3422 71612 3424 71632
rect 3424 71612 3476 71632
rect 3476 71612 3478 71632
rect 3422 71576 3478 71612
rect 11702 669976 11758 670032
rect 10414 669704 10470 669760
rect 2778 58520 2834 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 15842 673648 15898 673704
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 18602 669840 18658 669896
rect 29642 670656 29698 670712
rect 34242 672152 34298 672208
rect 47858 672288 47914 672344
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 535918 673784 535974 673840
rect 545026 673648 545082 673704
rect 39026 671336 39082 671392
rect 57334 671336 57390 671392
rect 89074 671336 89130 671392
rect 102874 671336 102930 671392
rect 116490 671336 116546 671392
rect 189630 671336 189686 671392
rect 394146 671336 394202 671392
rect 531226 671336 531282 671392
rect 540334 671336 540390 671392
rect 549350 671336 549406 671392
rect 554042 670792 554098 670848
rect 552846 669704 552902 669760
rect 555422 672152 555478 672208
rect 556802 670112 556858 670168
rect 560942 672288 560998 672344
rect 566554 670248 566610 670304
rect 569314 670384 569370 670440
rect 573454 670520 573510 670576
rect 579526 670656 579582 670712
rect 580170 644000 580226 644056
rect 579710 630808 579766 630864
rect 579802 617480 579858 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 537784 580226 537840
rect 578974 524456 579030 524512
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 431568 580226 431624
rect 579710 418240 579766 418296
rect 579802 404912 579858 404968
rect 579802 378392 579858 378448
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 580446 365064 580502 365120
rect 580354 258848 580410 258904
rect 580262 219000 580318 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 578882 179152 578938 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 4797 673842 4863 673845
rect 535913 673842 535979 673845
rect 4797 673840 535979 673842
rect 4797 673784 4802 673840
rect 4858 673784 535918 673840
rect 535974 673784 535979 673840
rect 4797 673782 535979 673784
rect 4797 673779 4863 673782
rect 535913 673779 535979 673782
rect 15837 673706 15903 673709
rect 545021 673706 545087 673709
rect 15837 673704 545087 673706
rect 15837 673648 15842 673704
rect 15898 673648 545026 673704
rect 545082 673648 545087 673704
rect 15837 673646 545087 673648
rect 15837 673643 15903 673646
rect 545021 673643 545087 673646
rect 47853 672346 47919 672349
rect 560937 672346 561003 672349
rect 47853 672344 561003 672346
rect 47853 672288 47858 672344
rect 47914 672288 560942 672344
rect 560998 672288 561003 672344
rect 47853 672286 561003 672288
rect 47853 672283 47919 672286
rect 560937 672283 561003 672286
rect 34237 672210 34303 672213
rect 555417 672210 555483 672213
rect 34237 672208 555483 672210
rect 34237 672152 34242 672208
rect 34298 672152 555422 672208
rect 555478 672152 555483 672208
rect 34237 672150 555483 672152
rect 34237 672147 34303 672150
rect 555417 672147 555483 672150
rect 39021 671396 39087 671397
rect 39021 671392 39068 671396
rect 39132 671394 39138 671396
rect 57329 671394 57395 671397
rect 89069 671396 89135 671397
rect 102869 671396 102935 671397
rect 116485 671396 116551 671397
rect -960 671258 480 671348
rect 39021 671336 39026 671392
rect 39021 671332 39068 671336
rect 39132 671334 39178 671394
rect 57329 671392 64890 671394
rect 57329 671336 57334 671392
rect 57390 671336 64890 671392
rect 57329 671334 64890 671336
rect 39132 671332 39138 671334
rect 39021 671331 39087 671332
rect 57329 671331 57395 671334
rect 3325 671258 3391 671261
rect -960 671256 3391 671258
rect -960 671200 3330 671256
rect 3386 671200 3391 671256
rect -960 671198 3391 671200
rect -960 671108 480 671198
rect 3325 671195 3391 671198
rect 64830 670850 64890 671334
rect 89069 671392 89116 671396
rect 89180 671394 89186 671396
rect 89069 671336 89074 671392
rect 89069 671332 89116 671336
rect 89180 671334 89226 671394
rect 102869 671392 102916 671396
rect 102980 671394 102986 671396
rect 102869 671336 102874 671392
rect 89180 671332 89186 671334
rect 102869 671332 102916 671336
rect 102980 671334 103026 671394
rect 116485 671392 116532 671396
rect 116596 671394 116602 671396
rect 189625 671394 189691 671397
rect 199694 671394 199700 671396
rect 116485 671336 116490 671392
rect 102980 671332 102986 671334
rect 116485 671332 116532 671336
rect 116596 671334 116642 671394
rect 189625 671392 199700 671394
rect 189625 671336 189630 671392
rect 189686 671336 199700 671392
rect 189625 671334 199700 671336
rect 116596 671332 116602 671334
rect 89069 671331 89135 671332
rect 102869 671331 102935 671332
rect 116485 671331 116551 671332
rect 189625 671331 189691 671334
rect 199694 671332 199700 671334
rect 199764 671332 199770 671396
rect 394141 671394 394207 671397
rect 393270 671392 394207 671394
rect 393270 671336 394146 671392
rect 394202 671336 394207 671392
rect 393270 671334 394207 671336
rect 199878 670924 199884 670988
rect 199948 670986 199954 670988
rect 393270 670986 393330 671334
rect 394141 671331 394207 671334
rect 529974 671332 529980 671396
rect 530044 671394 530050 671396
rect 531221 671394 531287 671397
rect 540329 671396 540395 671397
rect 549345 671396 549411 671397
rect 540278 671394 540284 671396
rect 530044 671392 531287 671394
rect 530044 671336 531226 671392
rect 531282 671336 531287 671392
rect 530044 671334 531287 671336
rect 540238 671334 540284 671394
rect 540348 671392 540395 671396
rect 549294 671394 549300 671396
rect 540390 671336 540395 671392
rect 530044 671332 530050 671334
rect 531221 671331 531287 671334
rect 540278 671332 540284 671334
rect 540348 671332 540395 671336
rect 549254 671334 549300 671394
rect 549364 671392 549411 671396
rect 549406 671336 549411 671392
rect 549294 671332 549300 671334
rect 549364 671332 549411 671336
rect 540329 671331 540395 671332
rect 549345 671331 549411 671332
rect 199948 670926 393330 670986
rect 199948 670924 199954 670926
rect 554037 670850 554103 670853
rect 64830 670848 554103 670850
rect 64830 670792 554042 670848
rect 554098 670792 554103 670848
rect 64830 670790 554103 670792
rect 554037 670787 554103 670790
rect 29637 670714 29703 670717
rect 529974 670714 529980 670716
rect 29637 670712 529980 670714
rect 29637 670656 29642 670712
rect 29698 670656 529980 670712
rect 29637 670654 529980 670656
rect 29637 670651 29703 670654
rect 529974 670652 529980 670654
rect 530044 670652 530050 670716
rect 579521 670714 579587 670717
rect 583520 670714 584960 670804
rect 579521 670712 584960 670714
rect 579521 670656 579526 670712
rect 579582 670656 584960 670712
rect 579521 670654 584960 670656
rect 579521 670651 579587 670654
rect 116526 670516 116532 670580
rect 116596 670578 116602 670580
rect 573449 670578 573515 670581
rect 116596 670576 573515 670578
rect 116596 670520 573454 670576
rect 573510 670520 573515 670576
rect 583520 670564 584960 670654
rect 116596 670518 573515 670520
rect 116596 670516 116602 670518
rect 573449 670515 573515 670518
rect 102910 670380 102916 670444
rect 102980 670442 102986 670444
rect 569309 670442 569375 670445
rect 102980 670440 569375 670442
rect 102980 670384 569314 670440
rect 569370 670384 569375 670440
rect 102980 670382 569375 670384
rect 102980 670380 102986 670382
rect 569309 670379 569375 670382
rect 89110 670244 89116 670308
rect 89180 670306 89186 670308
rect 566549 670306 566615 670309
rect 89180 670304 566615 670306
rect 89180 670248 566554 670304
rect 566610 670248 566615 670304
rect 89180 670246 566615 670248
rect 89180 670244 89186 670246
rect 566549 670243 566615 670246
rect 39062 670108 39068 670172
rect 39132 670170 39138 670172
rect 556797 670170 556863 670173
rect 39132 670168 556863 670170
rect 39132 670112 556802 670168
rect 556858 670112 556863 670168
rect 39132 670110 556863 670112
rect 39132 670108 39138 670110
rect 556797 670107 556863 670110
rect 11697 670034 11763 670037
rect 540278 670034 540284 670036
rect 11697 670032 540284 670034
rect 11697 669976 11702 670032
rect 11758 669976 540284 670032
rect 11697 669974 540284 669976
rect 11697 669971 11763 669974
rect 540278 669972 540284 669974
rect 540348 669972 540354 670036
rect 18597 669898 18663 669901
rect 549294 669898 549300 669900
rect 18597 669896 549300 669898
rect 18597 669840 18602 669896
rect 18658 669840 549300 669896
rect 18597 669838 549300 669840
rect 18597 669835 18663 669838
rect 549294 669836 549300 669838
rect 549364 669836 549370 669900
rect 10409 669762 10475 669765
rect 199878 669762 199884 669764
rect 10409 669760 199884 669762
rect 10409 669704 10414 669760
rect 10470 669704 199884 669760
rect 10409 669702 199884 669704
rect 10409 669699 10475 669702
rect 199878 669700 199884 669702
rect 199948 669700 199954 669764
rect 200062 669700 200068 669764
rect 200132 669762 200138 669764
rect 552841 669762 552907 669765
rect 200132 669760 552907 669762
rect 200132 669704 552846 669760
rect 552902 669704 552907 669760
rect 200132 669702 552907 669704
rect 200132 669700 200138 669702
rect 552841 669699 552907 669702
rect -960 658202 480 658292
rect 3325 658202 3391 658205
rect -960 658200 3391 658202
rect -960 658144 3330 658200
rect 3386 658144 3391 658200
rect -960 658142 3391 658144
rect -960 658052 480 658142
rect 3325 658139 3391 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3325 632090 3391 632093
rect -960 632088 3391 632090
rect -960 632032 3330 632088
rect 3386 632032 3391 632088
rect -960 632030 3391 632032
rect -960 631940 480 632030
rect 3325 632027 3391 632030
rect 579705 630866 579771 630869
rect 583520 630866 584960 630956
rect 579705 630864 584960 630866
rect 579705 630808 579710 630864
rect 579766 630808 584960 630864
rect 579705 630806 584960 630808
rect 579705 630803 579771 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3325 619170 3391 619173
rect -960 619168 3391 619170
rect -960 619112 3330 619168
rect 3386 619112 3391 619168
rect -960 619110 3391 619112
rect -960 619020 480 619110
rect 3325 619107 3391 619110
rect 579797 617538 579863 617541
rect 583520 617538 584960 617628
rect 579797 617536 584960 617538
rect 579797 617480 579802 617536
rect 579858 617480 584960 617536
rect 579797 617478 584960 617480
rect 579797 617475 579863 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3049 606114 3115 606117
rect -960 606112 3115 606114
rect -960 606056 3054 606112
rect 3110 606056 3115 606112
rect -960 606054 3115 606056
rect -960 605964 480 606054
rect 3049 606051 3115 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3141 566946 3207 566949
rect -960 566944 3207 566946
rect -960 566888 3146 566944
rect 3202 566888 3207 566944
rect -960 566886 3207 566888
rect -960 566796 480 566886
rect 3141 566883 3207 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 2957 553890 3023 553893
rect -960 553888 3023 553890
rect -960 553832 2962 553888
rect 3018 553832 3023 553888
rect -960 553830 3023 553832
rect -960 553740 480 553830
rect 2957 553827 3023 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3141 527914 3207 527917
rect -960 527912 3207 527914
rect -960 527856 3146 527912
rect 3202 527856 3207 527912
rect -960 527854 3207 527856
rect -960 527764 480 527854
rect 3141 527851 3207 527854
rect 578969 524514 579035 524517
rect 583520 524514 584960 524604
rect 578969 524512 584960 524514
rect 578969 524456 578974 524512
rect 579030 524456 584960 524512
rect 578969 524454 584960 524456
rect 578969 524451 579035 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2957 501802 3023 501805
rect -960 501800 3023 501802
rect -960 501744 2962 501800
rect 3018 501744 3023 501800
rect -960 501742 3023 501744
rect -960 501652 480 501742
rect 2957 501739 3023 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3233 475690 3299 475693
rect -960 475688 3299 475690
rect -960 475632 3238 475688
rect 3294 475632 3299 475688
rect -960 475630 3299 475632
rect -960 475540 480 475630
rect 3233 475627 3299 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3049 462634 3115 462637
rect -960 462632 3115 462634
rect -960 462576 3054 462632
rect 3110 462576 3115 462632
rect -960 462574 3115 462576
rect -960 462484 480 462574
rect 3049 462571 3115 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 579797 404970 579863 404973
rect 583520 404970 584960 405060
rect 579797 404968 584960 404970
rect 579797 404912 579802 404968
rect 579858 404912 584960 404968
rect 579797 404910 584960 404912
rect 579797 404907 579863 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580441 365122 580507 365125
rect 583520 365122 584960 365212
rect 580441 365120 584960 365122
rect 580441 365064 580446 365120
rect 580502 365064 584960 365120
rect 580441 365062 584960 365064
rect 580441 365059 580507 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 580349 258906 580415 258909
rect 583520 258906 584960 258996
rect 580349 258904 584960 258906
rect 580349 258848 580354 258904
rect 580410 258848 584960 258904
rect 580349 258846 584960 258848
rect 580349 258843 580415 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 578877 179210 578943 179213
rect 583520 179210 584960 179300
rect 578877 179208 584960 179210
rect 578877 179152 578882 179208
rect 578938 179152 584960 179208
rect 578877 179150 584960 179152
rect 578877 179147 578943 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2773 58578 2839 58581
rect -960 58576 2839 58578
rect -960 58520 2778 58576
rect 2834 58520 2839 58576
rect -960 58518 2839 58520
rect -960 58428 480 58518
rect 2773 58515 2839 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 39068 671392 39132 671396
rect 39068 671336 39082 671392
rect 39082 671336 39132 671392
rect 39068 671332 39132 671336
rect 89116 671392 89180 671396
rect 89116 671336 89130 671392
rect 89130 671336 89180 671392
rect 89116 671332 89180 671336
rect 102916 671392 102980 671396
rect 102916 671336 102930 671392
rect 102930 671336 102980 671392
rect 102916 671332 102980 671336
rect 116532 671392 116596 671396
rect 116532 671336 116546 671392
rect 116546 671336 116596 671392
rect 116532 671332 116596 671336
rect 199700 671332 199764 671396
rect 199884 670924 199948 670988
rect 529980 671332 530044 671396
rect 540284 671392 540348 671396
rect 540284 671336 540334 671392
rect 540334 671336 540348 671392
rect 540284 671332 540348 671336
rect 549300 671392 549364 671396
rect 549300 671336 549350 671392
rect 549350 671336 549364 671392
rect 549300 671332 549364 671336
rect 529980 670652 530044 670716
rect 116532 670516 116596 670580
rect 102916 670380 102980 670444
rect 89116 670244 89180 670308
rect 39068 670108 39132 670172
rect 540284 669972 540348 670036
rect 549300 669836 549364 669900
rect 199884 669700 199948 669764
rect 200068 669700 200132 669764
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 674000 31574 680058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 674000 38414 686898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 674000 42134 690618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 674000 45854 694338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 674000 49574 698058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 674000 56414 705242
rect 59514 674000 60134 707162
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 674000 63854 676338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 674000 67574 680058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 674000 74414 686898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 674000 78134 690618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 674000 81854 694338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 674000 85574 698058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 674000 92414 705242
rect 95514 674000 96134 707162
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 674000 99854 676338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 674000 103574 680058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 674000 110414 686898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 674000 114134 690618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 674000 117854 694338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 674000 121574 698058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 674000 128414 705242
rect 131514 674000 132134 707162
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 674000 135854 676338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 674000 139574 680058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 674000 146414 686898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 674000 150134 690618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 674000 153854 694338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 674000 157574 698058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 674000 164414 705242
rect 167514 674000 168134 707162
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 674000 171854 676338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 674000 175574 680058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 674000 182414 686898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 674000 186134 690618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 674000 189854 694338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 674000 193574 698058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 674000 200414 705242
rect 203514 674000 204134 707162
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 674000 207854 676338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 674000 211574 680058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 674000 218414 686898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 674000 222134 690618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 674000 225854 694338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 674000 229574 698058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 674000 236414 705242
rect 239514 674000 240134 707162
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 674000 243854 676338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 674000 247574 680058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 674000 254414 686898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 674000 258134 690618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 674000 261854 694338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 674000 265574 698058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 674000 272414 705242
rect 275514 674000 276134 707162
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 674000 279854 676338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 674000 283574 680058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 674000 290414 686898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 674000 294134 690618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 674000 297854 694338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 674000 301574 698058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 674000 308414 705242
rect 311514 674000 312134 707162
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 674000 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 674000 319574 680058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 674000 326414 686898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 674000 330134 690618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 674000 333854 694338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 674000 337574 698058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 674000 344414 705242
rect 347514 674000 348134 707162
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 674000 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 674000 355574 680058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 674000 362414 686898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 674000 366134 690618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 674000 369854 694338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 674000 373574 698058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 674000 380414 705242
rect 383514 674000 384134 707162
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 674000 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 674000 391574 680058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 674000 398414 686898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 674000 402134 690618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 674000 405854 694338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 674000 409574 698058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 674000 416414 705242
rect 419514 674000 420134 707162
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 674000 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 674000 427574 680058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 674000 434414 686898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 674000 438134 690618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 674000 441854 694338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 674000 445574 698058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 674000 452414 705242
rect 455514 674000 456134 707162
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 674000 459854 676338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 674000 463574 680058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 674000 470414 686898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 674000 474134 690618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 674000 477854 694338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 674000 481574 698058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 674000 488414 705242
rect 491514 674000 492134 707162
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 674000 495854 676338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 674000 499574 680058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 674000 506414 686898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 674000 510134 690618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 674000 513854 694338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 674000 517574 698058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 674000 524414 705242
rect 527514 674000 528134 707162
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 674000 531854 676338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 674000 535574 680058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 674000 542414 686898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 674000 546134 690618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 674000 549854 694338
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 674000 553574 698058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 39067 671396 39133 671397
rect 39067 671332 39068 671396
rect 39132 671332 39133 671396
rect 39067 671331 39133 671332
rect 89115 671396 89181 671397
rect 89115 671332 89116 671396
rect 89180 671332 89181 671396
rect 89115 671331 89181 671332
rect 102915 671396 102981 671397
rect 102915 671332 102916 671396
rect 102980 671332 102981 671396
rect 102915 671331 102981 671332
rect 116531 671396 116597 671397
rect 116531 671332 116532 671396
rect 116596 671332 116597 671396
rect 116531 671331 116597 671332
rect 199699 671396 199765 671397
rect 199699 671332 199700 671396
rect 199764 671332 199765 671396
rect 199699 671331 199765 671332
rect 529979 671396 530045 671397
rect 529979 671332 529980 671396
rect 530044 671332 530045 671396
rect 529979 671331 530045 671332
rect 540283 671396 540349 671397
rect 540283 671332 540284 671396
rect 540348 671332 540349 671396
rect 540283 671331 540349 671332
rect 549299 671396 549365 671397
rect 549299 671332 549300 671396
rect 549364 671332 549365 671396
rect 549299 671331 549365 671332
rect 39070 670173 39130 671331
rect 89118 670309 89178 671331
rect 102918 670445 102978 671331
rect 116534 670581 116594 671331
rect 116531 670580 116597 670581
rect 116531 670516 116532 670580
rect 116596 670516 116597 670580
rect 116531 670515 116597 670516
rect 102915 670444 102981 670445
rect 102915 670380 102916 670444
rect 102980 670380 102981 670444
rect 102915 670379 102981 670380
rect 89115 670308 89181 670309
rect 89115 670244 89116 670308
rect 89180 670244 89181 670308
rect 89115 670243 89181 670244
rect 39067 670172 39133 670173
rect 39067 670108 39068 670172
rect 39132 670108 39133 670172
rect 39067 670107 39133 670108
rect 199702 669490 199762 671331
rect 199883 670988 199949 670989
rect 199883 670924 199884 670988
rect 199948 670924 199949 670988
rect 199883 670923 199949 670924
rect 199886 669765 199946 670923
rect 529982 670717 530042 671331
rect 529979 670716 530045 670717
rect 529979 670652 529980 670716
rect 530044 670652 530045 670716
rect 529979 670651 530045 670652
rect 540286 670037 540346 671331
rect 540283 670036 540349 670037
rect 540283 669972 540284 670036
rect 540348 669972 540349 670036
rect 540283 669971 540349 669972
rect 549302 669901 549362 671331
rect 549299 669900 549365 669901
rect 549299 669836 549300 669900
rect 549364 669836 549365 669900
rect 549299 669835 549365 669836
rect 199883 669764 199949 669765
rect 199883 669700 199884 669764
rect 199948 669700 199949 669764
rect 199883 669699 199949 669700
rect 200067 669764 200133 669765
rect 200067 669700 200068 669764
rect 200132 669700 200133 669764
rect 200067 669699 200133 669700
rect 200070 669490 200130 669699
rect 51568 669454 51888 669486
rect 51568 669218 51610 669454
rect 51846 669218 51888 669454
rect 51568 669134 51888 669218
rect 51568 668898 51610 669134
rect 51846 668898 51888 669134
rect 51568 668866 51888 668898
rect 82288 669454 82608 669486
rect 82288 669218 82330 669454
rect 82566 669218 82608 669454
rect 82288 669134 82608 669218
rect 82288 668898 82330 669134
rect 82566 668898 82608 669134
rect 82288 668866 82608 668898
rect 113008 669454 113328 669486
rect 113008 669218 113050 669454
rect 113286 669218 113328 669454
rect 113008 669134 113328 669218
rect 113008 668898 113050 669134
rect 113286 668898 113328 669134
rect 113008 668866 113328 668898
rect 143728 669454 144048 669486
rect 143728 669218 143770 669454
rect 144006 669218 144048 669454
rect 143728 669134 144048 669218
rect 143728 668898 143770 669134
rect 144006 668898 144048 669134
rect 143728 668866 144048 668898
rect 174448 669454 174768 669486
rect 174448 669218 174490 669454
rect 174726 669218 174768 669454
rect 199702 669430 200130 669490
rect 205168 669454 205488 669486
rect 174448 669134 174768 669218
rect 174448 668898 174490 669134
rect 174726 668898 174768 669134
rect 174448 668866 174768 668898
rect 205168 669218 205210 669454
rect 205446 669218 205488 669454
rect 205168 669134 205488 669218
rect 205168 668898 205210 669134
rect 205446 668898 205488 669134
rect 205168 668866 205488 668898
rect 235888 669454 236208 669486
rect 235888 669218 235930 669454
rect 236166 669218 236208 669454
rect 235888 669134 236208 669218
rect 235888 668898 235930 669134
rect 236166 668898 236208 669134
rect 235888 668866 236208 668898
rect 266608 669454 266928 669486
rect 266608 669218 266650 669454
rect 266886 669218 266928 669454
rect 266608 669134 266928 669218
rect 266608 668898 266650 669134
rect 266886 668898 266928 669134
rect 266608 668866 266928 668898
rect 297328 669454 297648 669486
rect 297328 669218 297370 669454
rect 297606 669218 297648 669454
rect 297328 669134 297648 669218
rect 297328 668898 297370 669134
rect 297606 668898 297648 669134
rect 297328 668866 297648 668898
rect 328048 669454 328368 669486
rect 328048 669218 328090 669454
rect 328326 669218 328368 669454
rect 328048 669134 328368 669218
rect 328048 668898 328090 669134
rect 328326 668898 328368 669134
rect 328048 668866 328368 668898
rect 358768 669454 359088 669486
rect 358768 669218 358810 669454
rect 359046 669218 359088 669454
rect 358768 669134 359088 669218
rect 358768 668898 358810 669134
rect 359046 668898 359088 669134
rect 358768 668866 359088 668898
rect 389488 669454 389808 669486
rect 389488 669218 389530 669454
rect 389766 669218 389808 669454
rect 389488 669134 389808 669218
rect 389488 668898 389530 669134
rect 389766 668898 389808 669134
rect 389488 668866 389808 668898
rect 420208 669454 420528 669486
rect 420208 669218 420250 669454
rect 420486 669218 420528 669454
rect 420208 669134 420528 669218
rect 420208 668898 420250 669134
rect 420486 668898 420528 669134
rect 420208 668866 420528 668898
rect 450928 669454 451248 669486
rect 450928 669218 450970 669454
rect 451206 669218 451248 669454
rect 450928 669134 451248 669218
rect 450928 668898 450970 669134
rect 451206 668898 451248 669134
rect 450928 668866 451248 668898
rect 481648 669454 481968 669486
rect 481648 669218 481690 669454
rect 481926 669218 481968 669454
rect 481648 669134 481968 669218
rect 481648 668898 481690 669134
rect 481926 668898 481968 669134
rect 481648 668866 481968 668898
rect 512368 669454 512688 669486
rect 512368 669218 512410 669454
rect 512646 669218 512688 669454
rect 512368 669134 512688 669218
rect 512368 668898 512410 669134
rect 512646 668898 512688 669134
rect 512368 668866 512688 668898
rect 543088 669454 543408 669486
rect 543088 669218 543130 669454
rect 543366 669218 543408 669454
rect 543088 669134 543408 669218
rect 543088 668898 543130 669134
rect 543366 668898 543408 669134
rect 543088 668866 543408 668898
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 36208 651454 36528 651486
rect 36208 651218 36250 651454
rect 36486 651218 36528 651454
rect 36208 651134 36528 651218
rect 36208 650898 36250 651134
rect 36486 650898 36528 651134
rect 36208 650866 36528 650898
rect 66928 651454 67248 651486
rect 66928 651218 66970 651454
rect 67206 651218 67248 651454
rect 66928 651134 67248 651218
rect 66928 650898 66970 651134
rect 67206 650898 67248 651134
rect 66928 650866 67248 650898
rect 97648 651454 97968 651486
rect 97648 651218 97690 651454
rect 97926 651218 97968 651454
rect 97648 651134 97968 651218
rect 97648 650898 97690 651134
rect 97926 650898 97968 651134
rect 97648 650866 97968 650898
rect 128368 651454 128688 651486
rect 128368 651218 128410 651454
rect 128646 651218 128688 651454
rect 128368 651134 128688 651218
rect 128368 650898 128410 651134
rect 128646 650898 128688 651134
rect 128368 650866 128688 650898
rect 159088 651454 159408 651486
rect 159088 651218 159130 651454
rect 159366 651218 159408 651454
rect 159088 651134 159408 651218
rect 159088 650898 159130 651134
rect 159366 650898 159408 651134
rect 159088 650866 159408 650898
rect 189808 651454 190128 651486
rect 189808 651218 189850 651454
rect 190086 651218 190128 651454
rect 189808 651134 190128 651218
rect 189808 650898 189850 651134
rect 190086 650898 190128 651134
rect 189808 650866 190128 650898
rect 220528 651454 220848 651486
rect 220528 651218 220570 651454
rect 220806 651218 220848 651454
rect 220528 651134 220848 651218
rect 220528 650898 220570 651134
rect 220806 650898 220848 651134
rect 220528 650866 220848 650898
rect 251248 651454 251568 651486
rect 251248 651218 251290 651454
rect 251526 651218 251568 651454
rect 251248 651134 251568 651218
rect 251248 650898 251290 651134
rect 251526 650898 251568 651134
rect 251248 650866 251568 650898
rect 281968 651454 282288 651486
rect 281968 651218 282010 651454
rect 282246 651218 282288 651454
rect 281968 651134 282288 651218
rect 281968 650898 282010 651134
rect 282246 650898 282288 651134
rect 281968 650866 282288 650898
rect 312688 651454 313008 651486
rect 312688 651218 312730 651454
rect 312966 651218 313008 651454
rect 312688 651134 313008 651218
rect 312688 650898 312730 651134
rect 312966 650898 313008 651134
rect 312688 650866 313008 650898
rect 343408 651454 343728 651486
rect 343408 651218 343450 651454
rect 343686 651218 343728 651454
rect 343408 651134 343728 651218
rect 343408 650898 343450 651134
rect 343686 650898 343728 651134
rect 343408 650866 343728 650898
rect 374128 651454 374448 651486
rect 374128 651218 374170 651454
rect 374406 651218 374448 651454
rect 374128 651134 374448 651218
rect 374128 650898 374170 651134
rect 374406 650898 374448 651134
rect 374128 650866 374448 650898
rect 404848 651454 405168 651486
rect 404848 651218 404890 651454
rect 405126 651218 405168 651454
rect 404848 651134 405168 651218
rect 404848 650898 404890 651134
rect 405126 650898 405168 651134
rect 404848 650866 405168 650898
rect 435568 651454 435888 651486
rect 435568 651218 435610 651454
rect 435846 651218 435888 651454
rect 435568 651134 435888 651218
rect 435568 650898 435610 651134
rect 435846 650898 435888 651134
rect 435568 650866 435888 650898
rect 466288 651454 466608 651486
rect 466288 651218 466330 651454
rect 466566 651218 466608 651454
rect 466288 651134 466608 651218
rect 466288 650898 466330 651134
rect 466566 650898 466608 651134
rect 466288 650866 466608 650898
rect 497008 651454 497328 651486
rect 497008 651218 497050 651454
rect 497286 651218 497328 651454
rect 497008 651134 497328 651218
rect 497008 650898 497050 651134
rect 497286 650898 497328 651134
rect 497008 650866 497328 650898
rect 527728 651454 528048 651486
rect 527728 651218 527770 651454
rect 528006 651218 528048 651454
rect 527728 651134 528048 651218
rect 527728 650898 527770 651134
rect 528006 650898 528048 651134
rect 527728 650866 528048 650898
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 51568 633454 51888 633486
rect 51568 633218 51610 633454
rect 51846 633218 51888 633454
rect 51568 633134 51888 633218
rect 51568 632898 51610 633134
rect 51846 632898 51888 633134
rect 51568 632866 51888 632898
rect 82288 633454 82608 633486
rect 82288 633218 82330 633454
rect 82566 633218 82608 633454
rect 82288 633134 82608 633218
rect 82288 632898 82330 633134
rect 82566 632898 82608 633134
rect 82288 632866 82608 632898
rect 113008 633454 113328 633486
rect 113008 633218 113050 633454
rect 113286 633218 113328 633454
rect 113008 633134 113328 633218
rect 113008 632898 113050 633134
rect 113286 632898 113328 633134
rect 113008 632866 113328 632898
rect 143728 633454 144048 633486
rect 143728 633218 143770 633454
rect 144006 633218 144048 633454
rect 143728 633134 144048 633218
rect 143728 632898 143770 633134
rect 144006 632898 144048 633134
rect 143728 632866 144048 632898
rect 174448 633454 174768 633486
rect 174448 633218 174490 633454
rect 174726 633218 174768 633454
rect 174448 633134 174768 633218
rect 174448 632898 174490 633134
rect 174726 632898 174768 633134
rect 174448 632866 174768 632898
rect 205168 633454 205488 633486
rect 205168 633218 205210 633454
rect 205446 633218 205488 633454
rect 205168 633134 205488 633218
rect 205168 632898 205210 633134
rect 205446 632898 205488 633134
rect 205168 632866 205488 632898
rect 235888 633454 236208 633486
rect 235888 633218 235930 633454
rect 236166 633218 236208 633454
rect 235888 633134 236208 633218
rect 235888 632898 235930 633134
rect 236166 632898 236208 633134
rect 235888 632866 236208 632898
rect 266608 633454 266928 633486
rect 266608 633218 266650 633454
rect 266886 633218 266928 633454
rect 266608 633134 266928 633218
rect 266608 632898 266650 633134
rect 266886 632898 266928 633134
rect 266608 632866 266928 632898
rect 297328 633454 297648 633486
rect 297328 633218 297370 633454
rect 297606 633218 297648 633454
rect 297328 633134 297648 633218
rect 297328 632898 297370 633134
rect 297606 632898 297648 633134
rect 297328 632866 297648 632898
rect 328048 633454 328368 633486
rect 328048 633218 328090 633454
rect 328326 633218 328368 633454
rect 328048 633134 328368 633218
rect 328048 632898 328090 633134
rect 328326 632898 328368 633134
rect 328048 632866 328368 632898
rect 358768 633454 359088 633486
rect 358768 633218 358810 633454
rect 359046 633218 359088 633454
rect 358768 633134 359088 633218
rect 358768 632898 358810 633134
rect 359046 632898 359088 633134
rect 358768 632866 359088 632898
rect 389488 633454 389808 633486
rect 389488 633218 389530 633454
rect 389766 633218 389808 633454
rect 389488 633134 389808 633218
rect 389488 632898 389530 633134
rect 389766 632898 389808 633134
rect 389488 632866 389808 632898
rect 420208 633454 420528 633486
rect 420208 633218 420250 633454
rect 420486 633218 420528 633454
rect 420208 633134 420528 633218
rect 420208 632898 420250 633134
rect 420486 632898 420528 633134
rect 420208 632866 420528 632898
rect 450928 633454 451248 633486
rect 450928 633218 450970 633454
rect 451206 633218 451248 633454
rect 450928 633134 451248 633218
rect 450928 632898 450970 633134
rect 451206 632898 451248 633134
rect 450928 632866 451248 632898
rect 481648 633454 481968 633486
rect 481648 633218 481690 633454
rect 481926 633218 481968 633454
rect 481648 633134 481968 633218
rect 481648 632898 481690 633134
rect 481926 632898 481968 633134
rect 481648 632866 481968 632898
rect 512368 633454 512688 633486
rect 512368 633218 512410 633454
rect 512646 633218 512688 633454
rect 512368 633134 512688 633218
rect 512368 632898 512410 633134
rect 512646 632898 512688 633134
rect 512368 632866 512688 632898
rect 543088 633454 543408 633486
rect 543088 633218 543130 633454
rect 543366 633218 543408 633454
rect 543088 633134 543408 633218
rect 543088 632898 543130 633134
rect 543366 632898 543408 633134
rect 543088 632866 543408 632898
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 36208 615454 36528 615486
rect 36208 615218 36250 615454
rect 36486 615218 36528 615454
rect 36208 615134 36528 615218
rect 36208 614898 36250 615134
rect 36486 614898 36528 615134
rect 36208 614866 36528 614898
rect 66928 615454 67248 615486
rect 66928 615218 66970 615454
rect 67206 615218 67248 615454
rect 66928 615134 67248 615218
rect 66928 614898 66970 615134
rect 67206 614898 67248 615134
rect 66928 614866 67248 614898
rect 97648 615454 97968 615486
rect 97648 615218 97690 615454
rect 97926 615218 97968 615454
rect 97648 615134 97968 615218
rect 97648 614898 97690 615134
rect 97926 614898 97968 615134
rect 97648 614866 97968 614898
rect 128368 615454 128688 615486
rect 128368 615218 128410 615454
rect 128646 615218 128688 615454
rect 128368 615134 128688 615218
rect 128368 614898 128410 615134
rect 128646 614898 128688 615134
rect 128368 614866 128688 614898
rect 159088 615454 159408 615486
rect 159088 615218 159130 615454
rect 159366 615218 159408 615454
rect 159088 615134 159408 615218
rect 159088 614898 159130 615134
rect 159366 614898 159408 615134
rect 159088 614866 159408 614898
rect 189808 615454 190128 615486
rect 189808 615218 189850 615454
rect 190086 615218 190128 615454
rect 189808 615134 190128 615218
rect 189808 614898 189850 615134
rect 190086 614898 190128 615134
rect 189808 614866 190128 614898
rect 220528 615454 220848 615486
rect 220528 615218 220570 615454
rect 220806 615218 220848 615454
rect 220528 615134 220848 615218
rect 220528 614898 220570 615134
rect 220806 614898 220848 615134
rect 220528 614866 220848 614898
rect 251248 615454 251568 615486
rect 251248 615218 251290 615454
rect 251526 615218 251568 615454
rect 251248 615134 251568 615218
rect 251248 614898 251290 615134
rect 251526 614898 251568 615134
rect 251248 614866 251568 614898
rect 281968 615454 282288 615486
rect 281968 615218 282010 615454
rect 282246 615218 282288 615454
rect 281968 615134 282288 615218
rect 281968 614898 282010 615134
rect 282246 614898 282288 615134
rect 281968 614866 282288 614898
rect 312688 615454 313008 615486
rect 312688 615218 312730 615454
rect 312966 615218 313008 615454
rect 312688 615134 313008 615218
rect 312688 614898 312730 615134
rect 312966 614898 313008 615134
rect 312688 614866 313008 614898
rect 343408 615454 343728 615486
rect 343408 615218 343450 615454
rect 343686 615218 343728 615454
rect 343408 615134 343728 615218
rect 343408 614898 343450 615134
rect 343686 614898 343728 615134
rect 343408 614866 343728 614898
rect 374128 615454 374448 615486
rect 374128 615218 374170 615454
rect 374406 615218 374448 615454
rect 374128 615134 374448 615218
rect 374128 614898 374170 615134
rect 374406 614898 374448 615134
rect 374128 614866 374448 614898
rect 404848 615454 405168 615486
rect 404848 615218 404890 615454
rect 405126 615218 405168 615454
rect 404848 615134 405168 615218
rect 404848 614898 404890 615134
rect 405126 614898 405168 615134
rect 404848 614866 405168 614898
rect 435568 615454 435888 615486
rect 435568 615218 435610 615454
rect 435846 615218 435888 615454
rect 435568 615134 435888 615218
rect 435568 614898 435610 615134
rect 435846 614898 435888 615134
rect 435568 614866 435888 614898
rect 466288 615454 466608 615486
rect 466288 615218 466330 615454
rect 466566 615218 466608 615454
rect 466288 615134 466608 615218
rect 466288 614898 466330 615134
rect 466566 614898 466608 615134
rect 466288 614866 466608 614898
rect 497008 615454 497328 615486
rect 497008 615218 497050 615454
rect 497286 615218 497328 615454
rect 497008 615134 497328 615218
rect 497008 614898 497050 615134
rect 497286 614898 497328 615134
rect 497008 614866 497328 614898
rect 527728 615454 528048 615486
rect 527728 615218 527770 615454
rect 528006 615218 528048 615454
rect 527728 615134 528048 615218
rect 527728 614898 527770 615134
rect 528006 614898 528048 615134
rect 527728 614866 528048 614898
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 51568 597454 51888 597486
rect 51568 597218 51610 597454
rect 51846 597218 51888 597454
rect 51568 597134 51888 597218
rect 51568 596898 51610 597134
rect 51846 596898 51888 597134
rect 51568 596866 51888 596898
rect 82288 597454 82608 597486
rect 82288 597218 82330 597454
rect 82566 597218 82608 597454
rect 82288 597134 82608 597218
rect 82288 596898 82330 597134
rect 82566 596898 82608 597134
rect 82288 596866 82608 596898
rect 113008 597454 113328 597486
rect 113008 597218 113050 597454
rect 113286 597218 113328 597454
rect 113008 597134 113328 597218
rect 113008 596898 113050 597134
rect 113286 596898 113328 597134
rect 113008 596866 113328 596898
rect 143728 597454 144048 597486
rect 143728 597218 143770 597454
rect 144006 597218 144048 597454
rect 143728 597134 144048 597218
rect 143728 596898 143770 597134
rect 144006 596898 144048 597134
rect 143728 596866 144048 596898
rect 174448 597454 174768 597486
rect 174448 597218 174490 597454
rect 174726 597218 174768 597454
rect 174448 597134 174768 597218
rect 174448 596898 174490 597134
rect 174726 596898 174768 597134
rect 174448 596866 174768 596898
rect 205168 597454 205488 597486
rect 205168 597218 205210 597454
rect 205446 597218 205488 597454
rect 205168 597134 205488 597218
rect 205168 596898 205210 597134
rect 205446 596898 205488 597134
rect 205168 596866 205488 596898
rect 235888 597454 236208 597486
rect 235888 597218 235930 597454
rect 236166 597218 236208 597454
rect 235888 597134 236208 597218
rect 235888 596898 235930 597134
rect 236166 596898 236208 597134
rect 235888 596866 236208 596898
rect 266608 597454 266928 597486
rect 266608 597218 266650 597454
rect 266886 597218 266928 597454
rect 266608 597134 266928 597218
rect 266608 596898 266650 597134
rect 266886 596898 266928 597134
rect 266608 596866 266928 596898
rect 297328 597454 297648 597486
rect 297328 597218 297370 597454
rect 297606 597218 297648 597454
rect 297328 597134 297648 597218
rect 297328 596898 297370 597134
rect 297606 596898 297648 597134
rect 297328 596866 297648 596898
rect 328048 597454 328368 597486
rect 328048 597218 328090 597454
rect 328326 597218 328368 597454
rect 328048 597134 328368 597218
rect 328048 596898 328090 597134
rect 328326 596898 328368 597134
rect 328048 596866 328368 596898
rect 358768 597454 359088 597486
rect 358768 597218 358810 597454
rect 359046 597218 359088 597454
rect 358768 597134 359088 597218
rect 358768 596898 358810 597134
rect 359046 596898 359088 597134
rect 358768 596866 359088 596898
rect 389488 597454 389808 597486
rect 389488 597218 389530 597454
rect 389766 597218 389808 597454
rect 389488 597134 389808 597218
rect 389488 596898 389530 597134
rect 389766 596898 389808 597134
rect 389488 596866 389808 596898
rect 420208 597454 420528 597486
rect 420208 597218 420250 597454
rect 420486 597218 420528 597454
rect 420208 597134 420528 597218
rect 420208 596898 420250 597134
rect 420486 596898 420528 597134
rect 420208 596866 420528 596898
rect 450928 597454 451248 597486
rect 450928 597218 450970 597454
rect 451206 597218 451248 597454
rect 450928 597134 451248 597218
rect 450928 596898 450970 597134
rect 451206 596898 451248 597134
rect 450928 596866 451248 596898
rect 481648 597454 481968 597486
rect 481648 597218 481690 597454
rect 481926 597218 481968 597454
rect 481648 597134 481968 597218
rect 481648 596898 481690 597134
rect 481926 596898 481968 597134
rect 481648 596866 481968 596898
rect 512368 597454 512688 597486
rect 512368 597218 512410 597454
rect 512646 597218 512688 597454
rect 512368 597134 512688 597218
rect 512368 596898 512410 597134
rect 512646 596898 512688 597134
rect 512368 596866 512688 596898
rect 543088 597454 543408 597486
rect 543088 597218 543130 597454
rect 543366 597218 543408 597454
rect 543088 597134 543408 597218
rect 543088 596898 543130 597134
rect 543366 596898 543408 597134
rect 543088 596866 543408 596898
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 36208 579454 36528 579486
rect 36208 579218 36250 579454
rect 36486 579218 36528 579454
rect 36208 579134 36528 579218
rect 36208 578898 36250 579134
rect 36486 578898 36528 579134
rect 36208 578866 36528 578898
rect 66928 579454 67248 579486
rect 66928 579218 66970 579454
rect 67206 579218 67248 579454
rect 66928 579134 67248 579218
rect 66928 578898 66970 579134
rect 67206 578898 67248 579134
rect 66928 578866 67248 578898
rect 97648 579454 97968 579486
rect 97648 579218 97690 579454
rect 97926 579218 97968 579454
rect 97648 579134 97968 579218
rect 97648 578898 97690 579134
rect 97926 578898 97968 579134
rect 97648 578866 97968 578898
rect 128368 579454 128688 579486
rect 128368 579218 128410 579454
rect 128646 579218 128688 579454
rect 128368 579134 128688 579218
rect 128368 578898 128410 579134
rect 128646 578898 128688 579134
rect 128368 578866 128688 578898
rect 159088 579454 159408 579486
rect 159088 579218 159130 579454
rect 159366 579218 159408 579454
rect 159088 579134 159408 579218
rect 159088 578898 159130 579134
rect 159366 578898 159408 579134
rect 159088 578866 159408 578898
rect 189808 579454 190128 579486
rect 189808 579218 189850 579454
rect 190086 579218 190128 579454
rect 189808 579134 190128 579218
rect 189808 578898 189850 579134
rect 190086 578898 190128 579134
rect 189808 578866 190128 578898
rect 220528 579454 220848 579486
rect 220528 579218 220570 579454
rect 220806 579218 220848 579454
rect 220528 579134 220848 579218
rect 220528 578898 220570 579134
rect 220806 578898 220848 579134
rect 220528 578866 220848 578898
rect 251248 579454 251568 579486
rect 251248 579218 251290 579454
rect 251526 579218 251568 579454
rect 251248 579134 251568 579218
rect 251248 578898 251290 579134
rect 251526 578898 251568 579134
rect 251248 578866 251568 578898
rect 281968 579454 282288 579486
rect 281968 579218 282010 579454
rect 282246 579218 282288 579454
rect 281968 579134 282288 579218
rect 281968 578898 282010 579134
rect 282246 578898 282288 579134
rect 281968 578866 282288 578898
rect 312688 579454 313008 579486
rect 312688 579218 312730 579454
rect 312966 579218 313008 579454
rect 312688 579134 313008 579218
rect 312688 578898 312730 579134
rect 312966 578898 313008 579134
rect 312688 578866 313008 578898
rect 343408 579454 343728 579486
rect 343408 579218 343450 579454
rect 343686 579218 343728 579454
rect 343408 579134 343728 579218
rect 343408 578898 343450 579134
rect 343686 578898 343728 579134
rect 343408 578866 343728 578898
rect 374128 579454 374448 579486
rect 374128 579218 374170 579454
rect 374406 579218 374448 579454
rect 374128 579134 374448 579218
rect 374128 578898 374170 579134
rect 374406 578898 374448 579134
rect 374128 578866 374448 578898
rect 404848 579454 405168 579486
rect 404848 579218 404890 579454
rect 405126 579218 405168 579454
rect 404848 579134 405168 579218
rect 404848 578898 404890 579134
rect 405126 578898 405168 579134
rect 404848 578866 405168 578898
rect 435568 579454 435888 579486
rect 435568 579218 435610 579454
rect 435846 579218 435888 579454
rect 435568 579134 435888 579218
rect 435568 578898 435610 579134
rect 435846 578898 435888 579134
rect 435568 578866 435888 578898
rect 466288 579454 466608 579486
rect 466288 579218 466330 579454
rect 466566 579218 466608 579454
rect 466288 579134 466608 579218
rect 466288 578898 466330 579134
rect 466566 578898 466608 579134
rect 466288 578866 466608 578898
rect 497008 579454 497328 579486
rect 497008 579218 497050 579454
rect 497286 579218 497328 579454
rect 497008 579134 497328 579218
rect 497008 578898 497050 579134
rect 497286 578898 497328 579134
rect 497008 578866 497328 578898
rect 527728 579454 528048 579486
rect 527728 579218 527770 579454
rect 528006 579218 528048 579454
rect 527728 579134 528048 579218
rect 527728 578898 527770 579134
rect 528006 578898 528048 579134
rect 527728 578866 528048 578898
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 51568 561454 51888 561486
rect 51568 561218 51610 561454
rect 51846 561218 51888 561454
rect 51568 561134 51888 561218
rect 51568 560898 51610 561134
rect 51846 560898 51888 561134
rect 51568 560866 51888 560898
rect 82288 561454 82608 561486
rect 82288 561218 82330 561454
rect 82566 561218 82608 561454
rect 82288 561134 82608 561218
rect 82288 560898 82330 561134
rect 82566 560898 82608 561134
rect 82288 560866 82608 560898
rect 113008 561454 113328 561486
rect 113008 561218 113050 561454
rect 113286 561218 113328 561454
rect 113008 561134 113328 561218
rect 113008 560898 113050 561134
rect 113286 560898 113328 561134
rect 113008 560866 113328 560898
rect 143728 561454 144048 561486
rect 143728 561218 143770 561454
rect 144006 561218 144048 561454
rect 143728 561134 144048 561218
rect 143728 560898 143770 561134
rect 144006 560898 144048 561134
rect 143728 560866 144048 560898
rect 174448 561454 174768 561486
rect 174448 561218 174490 561454
rect 174726 561218 174768 561454
rect 174448 561134 174768 561218
rect 174448 560898 174490 561134
rect 174726 560898 174768 561134
rect 174448 560866 174768 560898
rect 205168 561454 205488 561486
rect 205168 561218 205210 561454
rect 205446 561218 205488 561454
rect 205168 561134 205488 561218
rect 205168 560898 205210 561134
rect 205446 560898 205488 561134
rect 205168 560866 205488 560898
rect 235888 561454 236208 561486
rect 235888 561218 235930 561454
rect 236166 561218 236208 561454
rect 235888 561134 236208 561218
rect 235888 560898 235930 561134
rect 236166 560898 236208 561134
rect 235888 560866 236208 560898
rect 266608 561454 266928 561486
rect 266608 561218 266650 561454
rect 266886 561218 266928 561454
rect 266608 561134 266928 561218
rect 266608 560898 266650 561134
rect 266886 560898 266928 561134
rect 266608 560866 266928 560898
rect 297328 561454 297648 561486
rect 297328 561218 297370 561454
rect 297606 561218 297648 561454
rect 297328 561134 297648 561218
rect 297328 560898 297370 561134
rect 297606 560898 297648 561134
rect 297328 560866 297648 560898
rect 328048 561454 328368 561486
rect 328048 561218 328090 561454
rect 328326 561218 328368 561454
rect 328048 561134 328368 561218
rect 328048 560898 328090 561134
rect 328326 560898 328368 561134
rect 328048 560866 328368 560898
rect 358768 561454 359088 561486
rect 358768 561218 358810 561454
rect 359046 561218 359088 561454
rect 358768 561134 359088 561218
rect 358768 560898 358810 561134
rect 359046 560898 359088 561134
rect 358768 560866 359088 560898
rect 389488 561454 389808 561486
rect 389488 561218 389530 561454
rect 389766 561218 389808 561454
rect 389488 561134 389808 561218
rect 389488 560898 389530 561134
rect 389766 560898 389808 561134
rect 389488 560866 389808 560898
rect 420208 561454 420528 561486
rect 420208 561218 420250 561454
rect 420486 561218 420528 561454
rect 420208 561134 420528 561218
rect 420208 560898 420250 561134
rect 420486 560898 420528 561134
rect 420208 560866 420528 560898
rect 450928 561454 451248 561486
rect 450928 561218 450970 561454
rect 451206 561218 451248 561454
rect 450928 561134 451248 561218
rect 450928 560898 450970 561134
rect 451206 560898 451248 561134
rect 450928 560866 451248 560898
rect 481648 561454 481968 561486
rect 481648 561218 481690 561454
rect 481926 561218 481968 561454
rect 481648 561134 481968 561218
rect 481648 560898 481690 561134
rect 481926 560898 481968 561134
rect 481648 560866 481968 560898
rect 512368 561454 512688 561486
rect 512368 561218 512410 561454
rect 512646 561218 512688 561454
rect 512368 561134 512688 561218
rect 512368 560898 512410 561134
rect 512646 560898 512688 561134
rect 512368 560866 512688 560898
rect 543088 561454 543408 561486
rect 543088 561218 543130 561454
rect 543366 561218 543408 561454
rect 543088 561134 543408 561218
rect 543088 560898 543130 561134
rect 543366 560898 543408 561134
rect 543088 560866 543408 560898
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 36208 543454 36528 543486
rect 36208 543218 36250 543454
rect 36486 543218 36528 543454
rect 36208 543134 36528 543218
rect 36208 542898 36250 543134
rect 36486 542898 36528 543134
rect 36208 542866 36528 542898
rect 66928 543454 67248 543486
rect 66928 543218 66970 543454
rect 67206 543218 67248 543454
rect 66928 543134 67248 543218
rect 66928 542898 66970 543134
rect 67206 542898 67248 543134
rect 66928 542866 67248 542898
rect 97648 543454 97968 543486
rect 97648 543218 97690 543454
rect 97926 543218 97968 543454
rect 97648 543134 97968 543218
rect 97648 542898 97690 543134
rect 97926 542898 97968 543134
rect 97648 542866 97968 542898
rect 128368 543454 128688 543486
rect 128368 543218 128410 543454
rect 128646 543218 128688 543454
rect 128368 543134 128688 543218
rect 128368 542898 128410 543134
rect 128646 542898 128688 543134
rect 128368 542866 128688 542898
rect 159088 543454 159408 543486
rect 159088 543218 159130 543454
rect 159366 543218 159408 543454
rect 159088 543134 159408 543218
rect 159088 542898 159130 543134
rect 159366 542898 159408 543134
rect 159088 542866 159408 542898
rect 189808 543454 190128 543486
rect 189808 543218 189850 543454
rect 190086 543218 190128 543454
rect 189808 543134 190128 543218
rect 189808 542898 189850 543134
rect 190086 542898 190128 543134
rect 189808 542866 190128 542898
rect 220528 543454 220848 543486
rect 220528 543218 220570 543454
rect 220806 543218 220848 543454
rect 220528 543134 220848 543218
rect 220528 542898 220570 543134
rect 220806 542898 220848 543134
rect 220528 542866 220848 542898
rect 251248 543454 251568 543486
rect 251248 543218 251290 543454
rect 251526 543218 251568 543454
rect 251248 543134 251568 543218
rect 251248 542898 251290 543134
rect 251526 542898 251568 543134
rect 251248 542866 251568 542898
rect 281968 543454 282288 543486
rect 281968 543218 282010 543454
rect 282246 543218 282288 543454
rect 281968 543134 282288 543218
rect 281968 542898 282010 543134
rect 282246 542898 282288 543134
rect 281968 542866 282288 542898
rect 312688 543454 313008 543486
rect 312688 543218 312730 543454
rect 312966 543218 313008 543454
rect 312688 543134 313008 543218
rect 312688 542898 312730 543134
rect 312966 542898 313008 543134
rect 312688 542866 313008 542898
rect 343408 543454 343728 543486
rect 343408 543218 343450 543454
rect 343686 543218 343728 543454
rect 343408 543134 343728 543218
rect 343408 542898 343450 543134
rect 343686 542898 343728 543134
rect 343408 542866 343728 542898
rect 374128 543454 374448 543486
rect 374128 543218 374170 543454
rect 374406 543218 374448 543454
rect 374128 543134 374448 543218
rect 374128 542898 374170 543134
rect 374406 542898 374448 543134
rect 374128 542866 374448 542898
rect 404848 543454 405168 543486
rect 404848 543218 404890 543454
rect 405126 543218 405168 543454
rect 404848 543134 405168 543218
rect 404848 542898 404890 543134
rect 405126 542898 405168 543134
rect 404848 542866 405168 542898
rect 435568 543454 435888 543486
rect 435568 543218 435610 543454
rect 435846 543218 435888 543454
rect 435568 543134 435888 543218
rect 435568 542898 435610 543134
rect 435846 542898 435888 543134
rect 435568 542866 435888 542898
rect 466288 543454 466608 543486
rect 466288 543218 466330 543454
rect 466566 543218 466608 543454
rect 466288 543134 466608 543218
rect 466288 542898 466330 543134
rect 466566 542898 466608 543134
rect 466288 542866 466608 542898
rect 497008 543454 497328 543486
rect 497008 543218 497050 543454
rect 497286 543218 497328 543454
rect 497008 543134 497328 543218
rect 497008 542898 497050 543134
rect 497286 542898 497328 543134
rect 497008 542866 497328 542898
rect 527728 543454 528048 543486
rect 527728 543218 527770 543454
rect 528006 543218 528048 543454
rect 527728 543134 528048 543218
rect 527728 542898 527770 543134
rect 528006 542898 528048 543134
rect 527728 542866 528048 542898
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 51568 525454 51888 525486
rect 51568 525218 51610 525454
rect 51846 525218 51888 525454
rect 51568 525134 51888 525218
rect 51568 524898 51610 525134
rect 51846 524898 51888 525134
rect 51568 524866 51888 524898
rect 82288 525454 82608 525486
rect 82288 525218 82330 525454
rect 82566 525218 82608 525454
rect 82288 525134 82608 525218
rect 82288 524898 82330 525134
rect 82566 524898 82608 525134
rect 82288 524866 82608 524898
rect 113008 525454 113328 525486
rect 113008 525218 113050 525454
rect 113286 525218 113328 525454
rect 113008 525134 113328 525218
rect 113008 524898 113050 525134
rect 113286 524898 113328 525134
rect 113008 524866 113328 524898
rect 143728 525454 144048 525486
rect 143728 525218 143770 525454
rect 144006 525218 144048 525454
rect 143728 525134 144048 525218
rect 143728 524898 143770 525134
rect 144006 524898 144048 525134
rect 143728 524866 144048 524898
rect 174448 525454 174768 525486
rect 174448 525218 174490 525454
rect 174726 525218 174768 525454
rect 174448 525134 174768 525218
rect 174448 524898 174490 525134
rect 174726 524898 174768 525134
rect 174448 524866 174768 524898
rect 205168 525454 205488 525486
rect 205168 525218 205210 525454
rect 205446 525218 205488 525454
rect 205168 525134 205488 525218
rect 205168 524898 205210 525134
rect 205446 524898 205488 525134
rect 205168 524866 205488 524898
rect 235888 525454 236208 525486
rect 235888 525218 235930 525454
rect 236166 525218 236208 525454
rect 235888 525134 236208 525218
rect 235888 524898 235930 525134
rect 236166 524898 236208 525134
rect 235888 524866 236208 524898
rect 266608 525454 266928 525486
rect 266608 525218 266650 525454
rect 266886 525218 266928 525454
rect 266608 525134 266928 525218
rect 266608 524898 266650 525134
rect 266886 524898 266928 525134
rect 266608 524866 266928 524898
rect 297328 525454 297648 525486
rect 297328 525218 297370 525454
rect 297606 525218 297648 525454
rect 297328 525134 297648 525218
rect 297328 524898 297370 525134
rect 297606 524898 297648 525134
rect 297328 524866 297648 524898
rect 328048 525454 328368 525486
rect 328048 525218 328090 525454
rect 328326 525218 328368 525454
rect 328048 525134 328368 525218
rect 328048 524898 328090 525134
rect 328326 524898 328368 525134
rect 328048 524866 328368 524898
rect 358768 525454 359088 525486
rect 358768 525218 358810 525454
rect 359046 525218 359088 525454
rect 358768 525134 359088 525218
rect 358768 524898 358810 525134
rect 359046 524898 359088 525134
rect 358768 524866 359088 524898
rect 389488 525454 389808 525486
rect 389488 525218 389530 525454
rect 389766 525218 389808 525454
rect 389488 525134 389808 525218
rect 389488 524898 389530 525134
rect 389766 524898 389808 525134
rect 389488 524866 389808 524898
rect 420208 525454 420528 525486
rect 420208 525218 420250 525454
rect 420486 525218 420528 525454
rect 420208 525134 420528 525218
rect 420208 524898 420250 525134
rect 420486 524898 420528 525134
rect 420208 524866 420528 524898
rect 450928 525454 451248 525486
rect 450928 525218 450970 525454
rect 451206 525218 451248 525454
rect 450928 525134 451248 525218
rect 450928 524898 450970 525134
rect 451206 524898 451248 525134
rect 450928 524866 451248 524898
rect 481648 525454 481968 525486
rect 481648 525218 481690 525454
rect 481926 525218 481968 525454
rect 481648 525134 481968 525218
rect 481648 524898 481690 525134
rect 481926 524898 481968 525134
rect 481648 524866 481968 524898
rect 512368 525454 512688 525486
rect 512368 525218 512410 525454
rect 512646 525218 512688 525454
rect 512368 525134 512688 525218
rect 512368 524898 512410 525134
rect 512646 524898 512688 525134
rect 512368 524866 512688 524898
rect 543088 525454 543408 525486
rect 543088 525218 543130 525454
rect 543366 525218 543408 525454
rect 543088 525134 543408 525218
rect 543088 524898 543130 525134
rect 543366 524898 543408 525134
rect 543088 524866 543408 524898
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 36208 507454 36528 507486
rect 36208 507218 36250 507454
rect 36486 507218 36528 507454
rect 36208 507134 36528 507218
rect 36208 506898 36250 507134
rect 36486 506898 36528 507134
rect 36208 506866 36528 506898
rect 66928 507454 67248 507486
rect 66928 507218 66970 507454
rect 67206 507218 67248 507454
rect 66928 507134 67248 507218
rect 66928 506898 66970 507134
rect 67206 506898 67248 507134
rect 66928 506866 67248 506898
rect 97648 507454 97968 507486
rect 97648 507218 97690 507454
rect 97926 507218 97968 507454
rect 97648 507134 97968 507218
rect 97648 506898 97690 507134
rect 97926 506898 97968 507134
rect 97648 506866 97968 506898
rect 128368 507454 128688 507486
rect 128368 507218 128410 507454
rect 128646 507218 128688 507454
rect 128368 507134 128688 507218
rect 128368 506898 128410 507134
rect 128646 506898 128688 507134
rect 128368 506866 128688 506898
rect 159088 507454 159408 507486
rect 159088 507218 159130 507454
rect 159366 507218 159408 507454
rect 159088 507134 159408 507218
rect 159088 506898 159130 507134
rect 159366 506898 159408 507134
rect 159088 506866 159408 506898
rect 189808 507454 190128 507486
rect 189808 507218 189850 507454
rect 190086 507218 190128 507454
rect 189808 507134 190128 507218
rect 189808 506898 189850 507134
rect 190086 506898 190128 507134
rect 189808 506866 190128 506898
rect 220528 507454 220848 507486
rect 220528 507218 220570 507454
rect 220806 507218 220848 507454
rect 220528 507134 220848 507218
rect 220528 506898 220570 507134
rect 220806 506898 220848 507134
rect 220528 506866 220848 506898
rect 251248 507454 251568 507486
rect 251248 507218 251290 507454
rect 251526 507218 251568 507454
rect 251248 507134 251568 507218
rect 251248 506898 251290 507134
rect 251526 506898 251568 507134
rect 251248 506866 251568 506898
rect 281968 507454 282288 507486
rect 281968 507218 282010 507454
rect 282246 507218 282288 507454
rect 281968 507134 282288 507218
rect 281968 506898 282010 507134
rect 282246 506898 282288 507134
rect 281968 506866 282288 506898
rect 312688 507454 313008 507486
rect 312688 507218 312730 507454
rect 312966 507218 313008 507454
rect 312688 507134 313008 507218
rect 312688 506898 312730 507134
rect 312966 506898 313008 507134
rect 312688 506866 313008 506898
rect 343408 507454 343728 507486
rect 343408 507218 343450 507454
rect 343686 507218 343728 507454
rect 343408 507134 343728 507218
rect 343408 506898 343450 507134
rect 343686 506898 343728 507134
rect 343408 506866 343728 506898
rect 374128 507454 374448 507486
rect 374128 507218 374170 507454
rect 374406 507218 374448 507454
rect 374128 507134 374448 507218
rect 374128 506898 374170 507134
rect 374406 506898 374448 507134
rect 374128 506866 374448 506898
rect 404848 507454 405168 507486
rect 404848 507218 404890 507454
rect 405126 507218 405168 507454
rect 404848 507134 405168 507218
rect 404848 506898 404890 507134
rect 405126 506898 405168 507134
rect 404848 506866 405168 506898
rect 435568 507454 435888 507486
rect 435568 507218 435610 507454
rect 435846 507218 435888 507454
rect 435568 507134 435888 507218
rect 435568 506898 435610 507134
rect 435846 506898 435888 507134
rect 435568 506866 435888 506898
rect 466288 507454 466608 507486
rect 466288 507218 466330 507454
rect 466566 507218 466608 507454
rect 466288 507134 466608 507218
rect 466288 506898 466330 507134
rect 466566 506898 466608 507134
rect 466288 506866 466608 506898
rect 497008 507454 497328 507486
rect 497008 507218 497050 507454
rect 497286 507218 497328 507454
rect 497008 507134 497328 507218
rect 497008 506898 497050 507134
rect 497286 506898 497328 507134
rect 497008 506866 497328 506898
rect 527728 507454 528048 507486
rect 527728 507218 527770 507454
rect 528006 507218 528048 507454
rect 527728 507134 528048 507218
rect 527728 506898 527770 507134
rect 528006 506898 528048 507134
rect 527728 506866 528048 506898
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 51568 489454 51888 489486
rect 51568 489218 51610 489454
rect 51846 489218 51888 489454
rect 51568 489134 51888 489218
rect 51568 488898 51610 489134
rect 51846 488898 51888 489134
rect 51568 488866 51888 488898
rect 82288 489454 82608 489486
rect 82288 489218 82330 489454
rect 82566 489218 82608 489454
rect 82288 489134 82608 489218
rect 82288 488898 82330 489134
rect 82566 488898 82608 489134
rect 82288 488866 82608 488898
rect 113008 489454 113328 489486
rect 113008 489218 113050 489454
rect 113286 489218 113328 489454
rect 113008 489134 113328 489218
rect 113008 488898 113050 489134
rect 113286 488898 113328 489134
rect 113008 488866 113328 488898
rect 143728 489454 144048 489486
rect 143728 489218 143770 489454
rect 144006 489218 144048 489454
rect 143728 489134 144048 489218
rect 143728 488898 143770 489134
rect 144006 488898 144048 489134
rect 143728 488866 144048 488898
rect 174448 489454 174768 489486
rect 174448 489218 174490 489454
rect 174726 489218 174768 489454
rect 174448 489134 174768 489218
rect 174448 488898 174490 489134
rect 174726 488898 174768 489134
rect 174448 488866 174768 488898
rect 205168 489454 205488 489486
rect 205168 489218 205210 489454
rect 205446 489218 205488 489454
rect 205168 489134 205488 489218
rect 205168 488898 205210 489134
rect 205446 488898 205488 489134
rect 205168 488866 205488 488898
rect 235888 489454 236208 489486
rect 235888 489218 235930 489454
rect 236166 489218 236208 489454
rect 235888 489134 236208 489218
rect 235888 488898 235930 489134
rect 236166 488898 236208 489134
rect 235888 488866 236208 488898
rect 266608 489454 266928 489486
rect 266608 489218 266650 489454
rect 266886 489218 266928 489454
rect 266608 489134 266928 489218
rect 266608 488898 266650 489134
rect 266886 488898 266928 489134
rect 266608 488866 266928 488898
rect 297328 489454 297648 489486
rect 297328 489218 297370 489454
rect 297606 489218 297648 489454
rect 297328 489134 297648 489218
rect 297328 488898 297370 489134
rect 297606 488898 297648 489134
rect 297328 488866 297648 488898
rect 328048 489454 328368 489486
rect 328048 489218 328090 489454
rect 328326 489218 328368 489454
rect 328048 489134 328368 489218
rect 328048 488898 328090 489134
rect 328326 488898 328368 489134
rect 328048 488866 328368 488898
rect 358768 489454 359088 489486
rect 358768 489218 358810 489454
rect 359046 489218 359088 489454
rect 358768 489134 359088 489218
rect 358768 488898 358810 489134
rect 359046 488898 359088 489134
rect 358768 488866 359088 488898
rect 389488 489454 389808 489486
rect 389488 489218 389530 489454
rect 389766 489218 389808 489454
rect 389488 489134 389808 489218
rect 389488 488898 389530 489134
rect 389766 488898 389808 489134
rect 389488 488866 389808 488898
rect 420208 489454 420528 489486
rect 420208 489218 420250 489454
rect 420486 489218 420528 489454
rect 420208 489134 420528 489218
rect 420208 488898 420250 489134
rect 420486 488898 420528 489134
rect 420208 488866 420528 488898
rect 450928 489454 451248 489486
rect 450928 489218 450970 489454
rect 451206 489218 451248 489454
rect 450928 489134 451248 489218
rect 450928 488898 450970 489134
rect 451206 488898 451248 489134
rect 450928 488866 451248 488898
rect 481648 489454 481968 489486
rect 481648 489218 481690 489454
rect 481926 489218 481968 489454
rect 481648 489134 481968 489218
rect 481648 488898 481690 489134
rect 481926 488898 481968 489134
rect 481648 488866 481968 488898
rect 512368 489454 512688 489486
rect 512368 489218 512410 489454
rect 512646 489218 512688 489454
rect 512368 489134 512688 489218
rect 512368 488898 512410 489134
rect 512646 488898 512688 489134
rect 512368 488866 512688 488898
rect 543088 489454 543408 489486
rect 543088 489218 543130 489454
rect 543366 489218 543408 489454
rect 543088 489134 543408 489218
rect 543088 488898 543130 489134
rect 543366 488898 543408 489134
rect 543088 488866 543408 488898
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 36208 471454 36528 471486
rect 36208 471218 36250 471454
rect 36486 471218 36528 471454
rect 36208 471134 36528 471218
rect 36208 470898 36250 471134
rect 36486 470898 36528 471134
rect 36208 470866 36528 470898
rect 66928 471454 67248 471486
rect 66928 471218 66970 471454
rect 67206 471218 67248 471454
rect 66928 471134 67248 471218
rect 66928 470898 66970 471134
rect 67206 470898 67248 471134
rect 66928 470866 67248 470898
rect 97648 471454 97968 471486
rect 97648 471218 97690 471454
rect 97926 471218 97968 471454
rect 97648 471134 97968 471218
rect 97648 470898 97690 471134
rect 97926 470898 97968 471134
rect 97648 470866 97968 470898
rect 128368 471454 128688 471486
rect 128368 471218 128410 471454
rect 128646 471218 128688 471454
rect 128368 471134 128688 471218
rect 128368 470898 128410 471134
rect 128646 470898 128688 471134
rect 128368 470866 128688 470898
rect 159088 471454 159408 471486
rect 159088 471218 159130 471454
rect 159366 471218 159408 471454
rect 159088 471134 159408 471218
rect 159088 470898 159130 471134
rect 159366 470898 159408 471134
rect 159088 470866 159408 470898
rect 189808 471454 190128 471486
rect 189808 471218 189850 471454
rect 190086 471218 190128 471454
rect 189808 471134 190128 471218
rect 189808 470898 189850 471134
rect 190086 470898 190128 471134
rect 189808 470866 190128 470898
rect 220528 471454 220848 471486
rect 220528 471218 220570 471454
rect 220806 471218 220848 471454
rect 220528 471134 220848 471218
rect 220528 470898 220570 471134
rect 220806 470898 220848 471134
rect 220528 470866 220848 470898
rect 251248 471454 251568 471486
rect 251248 471218 251290 471454
rect 251526 471218 251568 471454
rect 251248 471134 251568 471218
rect 251248 470898 251290 471134
rect 251526 470898 251568 471134
rect 251248 470866 251568 470898
rect 281968 471454 282288 471486
rect 281968 471218 282010 471454
rect 282246 471218 282288 471454
rect 281968 471134 282288 471218
rect 281968 470898 282010 471134
rect 282246 470898 282288 471134
rect 281968 470866 282288 470898
rect 312688 471454 313008 471486
rect 312688 471218 312730 471454
rect 312966 471218 313008 471454
rect 312688 471134 313008 471218
rect 312688 470898 312730 471134
rect 312966 470898 313008 471134
rect 312688 470866 313008 470898
rect 343408 471454 343728 471486
rect 343408 471218 343450 471454
rect 343686 471218 343728 471454
rect 343408 471134 343728 471218
rect 343408 470898 343450 471134
rect 343686 470898 343728 471134
rect 343408 470866 343728 470898
rect 374128 471454 374448 471486
rect 374128 471218 374170 471454
rect 374406 471218 374448 471454
rect 374128 471134 374448 471218
rect 374128 470898 374170 471134
rect 374406 470898 374448 471134
rect 374128 470866 374448 470898
rect 404848 471454 405168 471486
rect 404848 471218 404890 471454
rect 405126 471218 405168 471454
rect 404848 471134 405168 471218
rect 404848 470898 404890 471134
rect 405126 470898 405168 471134
rect 404848 470866 405168 470898
rect 435568 471454 435888 471486
rect 435568 471218 435610 471454
rect 435846 471218 435888 471454
rect 435568 471134 435888 471218
rect 435568 470898 435610 471134
rect 435846 470898 435888 471134
rect 435568 470866 435888 470898
rect 466288 471454 466608 471486
rect 466288 471218 466330 471454
rect 466566 471218 466608 471454
rect 466288 471134 466608 471218
rect 466288 470898 466330 471134
rect 466566 470898 466608 471134
rect 466288 470866 466608 470898
rect 497008 471454 497328 471486
rect 497008 471218 497050 471454
rect 497286 471218 497328 471454
rect 497008 471134 497328 471218
rect 497008 470898 497050 471134
rect 497286 470898 497328 471134
rect 497008 470866 497328 470898
rect 527728 471454 528048 471486
rect 527728 471218 527770 471454
rect 528006 471218 528048 471454
rect 527728 471134 528048 471218
rect 527728 470898 527770 471134
rect 528006 470898 528048 471134
rect 527728 470866 528048 470898
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 51568 453454 51888 453486
rect 51568 453218 51610 453454
rect 51846 453218 51888 453454
rect 51568 453134 51888 453218
rect 51568 452898 51610 453134
rect 51846 452898 51888 453134
rect 51568 452866 51888 452898
rect 82288 453454 82608 453486
rect 82288 453218 82330 453454
rect 82566 453218 82608 453454
rect 82288 453134 82608 453218
rect 82288 452898 82330 453134
rect 82566 452898 82608 453134
rect 82288 452866 82608 452898
rect 113008 453454 113328 453486
rect 113008 453218 113050 453454
rect 113286 453218 113328 453454
rect 113008 453134 113328 453218
rect 113008 452898 113050 453134
rect 113286 452898 113328 453134
rect 113008 452866 113328 452898
rect 143728 453454 144048 453486
rect 143728 453218 143770 453454
rect 144006 453218 144048 453454
rect 143728 453134 144048 453218
rect 143728 452898 143770 453134
rect 144006 452898 144048 453134
rect 143728 452866 144048 452898
rect 174448 453454 174768 453486
rect 174448 453218 174490 453454
rect 174726 453218 174768 453454
rect 174448 453134 174768 453218
rect 174448 452898 174490 453134
rect 174726 452898 174768 453134
rect 174448 452866 174768 452898
rect 205168 453454 205488 453486
rect 205168 453218 205210 453454
rect 205446 453218 205488 453454
rect 205168 453134 205488 453218
rect 205168 452898 205210 453134
rect 205446 452898 205488 453134
rect 205168 452866 205488 452898
rect 235888 453454 236208 453486
rect 235888 453218 235930 453454
rect 236166 453218 236208 453454
rect 235888 453134 236208 453218
rect 235888 452898 235930 453134
rect 236166 452898 236208 453134
rect 235888 452866 236208 452898
rect 266608 453454 266928 453486
rect 266608 453218 266650 453454
rect 266886 453218 266928 453454
rect 266608 453134 266928 453218
rect 266608 452898 266650 453134
rect 266886 452898 266928 453134
rect 266608 452866 266928 452898
rect 297328 453454 297648 453486
rect 297328 453218 297370 453454
rect 297606 453218 297648 453454
rect 297328 453134 297648 453218
rect 297328 452898 297370 453134
rect 297606 452898 297648 453134
rect 297328 452866 297648 452898
rect 328048 453454 328368 453486
rect 328048 453218 328090 453454
rect 328326 453218 328368 453454
rect 328048 453134 328368 453218
rect 328048 452898 328090 453134
rect 328326 452898 328368 453134
rect 328048 452866 328368 452898
rect 358768 453454 359088 453486
rect 358768 453218 358810 453454
rect 359046 453218 359088 453454
rect 358768 453134 359088 453218
rect 358768 452898 358810 453134
rect 359046 452898 359088 453134
rect 358768 452866 359088 452898
rect 389488 453454 389808 453486
rect 389488 453218 389530 453454
rect 389766 453218 389808 453454
rect 389488 453134 389808 453218
rect 389488 452898 389530 453134
rect 389766 452898 389808 453134
rect 389488 452866 389808 452898
rect 420208 453454 420528 453486
rect 420208 453218 420250 453454
rect 420486 453218 420528 453454
rect 420208 453134 420528 453218
rect 420208 452898 420250 453134
rect 420486 452898 420528 453134
rect 420208 452866 420528 452898
rect 450928 453454 451248 453486
rect 450928 453218 450970 453454
rect 451206 453218 451248 453454
rect 450928 453134 451248 453218
rect 450928 452898 450970 453134
rect 451206 452898 451248 453134
rect 450928 452866 451248 452898
rect 481648 453454 481968 453486
rect 481648 453218 481690 453454
rect 481926 453218 481968 453454
rect 481648 453134 481968 453218
rect 481648 452898 481690 453134
rect 481926 452898 481968 453134
rect 481648 452866 481968 452898
rect 512368 453454 512688 453486
rect 512368 453218 512410 453454
rect 512646 453218 512688 453454
rect 512368 453134 512688 453218
rect 512368 452898 512410 453134
rect 512646 452898 512688 453134
rect 512368 452866 512688 452898
rect 543088 453454 543408 453486
rect 543088 453218 543130 453454
rect 543366 453218 543408 453454
rect 543088 453134 543408 453218
rect 543088 452898 543130 453134
rect 543366 452898 543408 453134
rect 543088 452866 543408 452898
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 36208 435454 36528 435486
rect 36208 435218 36250 435454
rect 36486 435218 36528 435454
rect 36208 435134 36528 435218
rect 36208 434898 36250 435134
rect 36486 434898 36528 435134
rect 36208 434866 36528 434898
rect 66928 435454 67248 435486
rect 66928 435218 66970 435454
rect 67206 435218 67248 435454
rect 66928 435134 67248 435218
rect 66928 434898 66970 435134
rect 67206 434898 67248 435134
rect 66928 434866 67248 434898
rect 97648 435454 97968 435486
rect 97648 435218 97690 435454
rect 97926 435218 97968 435454
rect 97648 435134 97968 435218
rect 97648 434898 97690 435134
rect 97926 434898 97968 435134
rect 97648 434866 97968 434898
rect 128368 435454 128688 435486
rect 128368 435218 128410 435454
rect 128646 435218 128688 435454
rect 128368 435134 128688 435218
rect 128368 434898 128410 435134
rect 128646 434898 128688 435134
rect 128368 434866 128688 434898
rect 159088 435454 159408 435486
rect 159088 435218 159130 435454
rect 159366 435218 159408 435454
rect 159088 435134 159408 435218
rect 159088 434898 159130 435134
rect 159366 434898 159408 435134
rect 159088 434866 159408 434898
rect 189808 435454 190128 435486
rect 189808 435218 189850 435454
rect 190086 435218 190128 435454
rect 189808 435134 190128 435218
rect 189808 434898 189850 435134
rect 190086 434898 190128 435134
rect 189808 434866 190128 434898
rect 220528 435454 220848 435486
rect 220528 435218 220570 435454
rect 220806 435218 220848 435454
rect 220528 435134 220848 435218
rect 220528 434898 220570 435134
rect 220806 434898 220848 435134
rect 220528 434866 220848 434898
rect 251248 435454 251568 435486
rect 251248 435218 251290 435454
rect 251526 435218 251568 435454
rect 251248 435134 251568 435218
rect 251248 434898 251290 435134
rect 251526 434898 251568 435134
rect 251248 434866 251568 434898
rect 281968 435454 282288 435486
rect 281968 435218 282010 435454
rect 282246 435218 282288 435454
rect 281968 435134 282288 435218
rect 281968 434898 282010 435134
rect 282246 434898 282288 435134
rect 281968 434866 282288 434898
rect 312688 435454 313008 435486
rect 312688 435218 312730 435454
rect 312966 435218 313008 435454
rect 312688 435134 313008 435218
rect 312688 434898 312730 435134
rect 312966 434898 313008 435134
rect 312688 434866 313008 434898
rect 343408 435454 343728 435486
rect 343408 435218 343450 435454
rect 343686 435218 343728 435454
rect 343408 435134 343728 435218
rect 343408 434898 343450 435134
rect 343686 434898 343728 435134
rect 343408 434866 343728 434898
rect 374128 435454 374448 435486
rect 374128 435218 374170 435454
rect 374406 435218 374448 435454
rect 374128 435134 374448 435218
rect 374128 434898 374170 435134
rect 374406 434898 374448 435134
rect 374128 434866 374448 434898
rect 404848 435454 405168 435486
rect 404848 435218 404890 435454
rect 405126 435218 405168 435454
rect 404848 435134 405168 435218
rect 404848 434898 404890 435134
rect 405126 434898 405168 435134
rect 404848 434866 405168 434898
rect 435568 435454 435888 435486
rect 435568 435218 435610 435454
rect 435846 435218 435888 435454
rect 435568 435134 435888 435218
rect 435568 434898 435610 435134
rect 435846 434898 435888 435134
rect 435568 434866 435888 434898
rect 466288 435454 466608 435486
rect 466288 435218 466330 435454
rect 466566 435218 466608 435454
rect 466288 435134 466608 435218
rect 466288 434898 466330 435134
rect 466566 434898 466608 435134
rect 466288 434866 466608 434898
rect 497008 435454 497328 435486
rect 497008 435218 497050 435454
rect 497286 435218 497328 435454
rect 497008 435134 497328 435218
rect 497008 434898 497050 435134
rect 497286 434898 497328 435134
rect 497008 434866 497328 434898
rect 527728 435454 528048 435486
rect 527728 435218 527770 435454
rect 528006 435218 528048 435454
rect 527728 435134 528048 435218
rect 527728 434898 527770 435134
rect 528006 434898 528048 435134
rect 527728 434866 528048 434898
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 51568 417454 51888 417486
rect 51568 417218 51610 417454
rect 51846 417218 51888 417454
rect 51568 417134 51888 417218
rect 51568 416898 51610 417134
rect 51846 416898 51888 417134
rect 51568 416866 51888 416898
rect 82288 417454 82608 417486
rect 82288 417218 82330 417454
rect 82566 417218 82608 417454
rect 82288 417134 82608 417218
rect 82288 416898 82330 417134
rect 82566 416898 82608 417134
rect 82288 416866 82608 416898
rect 113008 417454 113328 417486
rect 113008 417218 113050 417454
rect 113286 417218 113328 417454
rect 113008 417134 113328 417218
rect 113008 416898 113050 417134
rect 113286 416898 113328 417134
rect 113008 416866 113328 416898
rect 143728 417454 144048 417486
rect 143728 417218 143770 417454
rect 144006 417218 144048 417454
rect 143728 417134 144048 417218
rect 143728 416898 143770 417134
rect 144006 416898 144048 417134
rect 143728 416866 144048 416898
rect 174448 417454 174768 417486
rect 174448 417218 174490 417454
rect 174726 417218 174768 417454
rect 174448 417134 174768 417218
rect 174448 416898 174490 417134
rect 174726 416898 174768 417134
rect 174448 416866 174768 416898
rect 205168 417454 205488 417486
rect 205168 417218 205210 417454
rect 205446 417218 205488 417454
rect 205168 417134 205488 417218
rect 205168 416898 205210 417134
rect 205446 416898 205488 417134
rect 205168 416866 205488 416898
rect 235888 417454 236208 417486
rect 235888 417218 235930 417454
rect 236166 417218 236208 417454
rect 235888 417134 236208 417218
rect 235888 416898 235930 417134
rect 236166 416898 236208 417134
rect 235888 416866 236208 416898
rect 266608 417454 266928 417486
rect 266608 417218 266650 417454
rect 266886 417218 266928 417454
rect 266608 417134 266928 417218
rect 266608 416898 266650 417134
rect 266886 416898 266928 417134
rect 266608 416866 266928 416898
rect 297328 417454 297648 417486
rect 297328 417218 297370 417454
rect 297606 417218 297648 417454
rect 297328 417134 297648 417218
rect 297328 416898 297370 417134
rect 297606 416898 297648 417134
rect 297328 416866 297648 416898
rect 328048 417454 328368 417486
rect 328048 417218 328090 417454
rect 328326 417218 328368 417454
rect 328048 417134 328368 417218
rect 328048 416898 328090 417134
rect 328326 416898 328368 417134
rect 328048 416866 328368 416898
rect 358768 417454 359088 417486
rect 358768 417218 358810 417454
rect 359046 417218 359088 417454
rect 358768 417134 359088 417218
rect 358768 416898 358810 417134
rect 359046 416898 359088 417134
rect 358768 416866 359088 416898
rect 389488 417454 389808 417486
rect 389488 417218 389530 417454
rect 389766 417218 389808 417454
rect 389488 417134 389808 417218
rect 389488 416898 389530 417134
rect 389766 416898 389808 417134
rect 389488 416866 389808 416898
rect 420208 417454 420528 417486
rect 420208 417218 420250 417454
rect 420486 417218 420528 417454
rect 420208 417134 420528 417218
rect 420208 416898 420250 417134
rect 420486 416898 420528 417134
rect 420208 416866 420528 416898
rect 450928 417454 451248 417486
rect 450928 417218 450970 417454
rect 451206 417218 451248 417454
rect 450928 417134 451248 417218
rect 450928 416898 450970 417134
rect 451206 416898 451248 417134
rect 450928 416866 451248 416898
rect 481648 417454 481968 417486
rect 481648 417218 481690 417454
rect 481926 417218 481968 417454
rect 481648 417134 481968 417218
rect 481648 416898 481690 417134
rect 481926 416898 481968 417134
rect 481648 416866 481968 416898
rect 512368 417454 512688 417486
rect 512368 417218 512410 417454
rect 512646 417218 512688 417454
rect 512368 417134 512688 417218
rect 512368 416898 512410 417134
rect 512646 416898 512688 417134
rect 512368 416866 512688 416898
rect 543088 417454 543408 417486
rect 543088 417218 543130 417454
rect 543366 417218 543408 417454
rect 543088 417134 543408 417218
rect 543088 416898 543130 417134
rect 543366 416898 543408 417134
rect 543088 416866 543408 416898
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 36208 399454 36528 399486
rect 36208 399218 36250 399454
rect 36486 399218 36528 399454
rect 36208 399134 36528 399218
rect 36208 398898 36250 399134
rect 36486 398898 36528 399134
rect 36208 398866 36528 398898
rect 66928 399454 67248 399486
rect 66928 399218 66970 399454
rect 67206 399218 67248 399454
rect 66928 399134 67248 399218
rect 66928 398898 66970 399134
rect 67206 398898 67248 399134
rect 66928 398866 67248 398898
rect 97648 399454 97968 399486
rect 97648 399218 97690 399454
rect 97926 399218 97968 399454
rect 97648 399134 97968 399218
rect 97648 398898 97690 399134
rect 97926 398898 97968 399134
rect 97648 398866 97968 398898
rect 128368 399454 128688 399486
rect 128368 399218 128410 399454
rect 128646 399218 128688 399454
rect 128368 399134 128688 399218
rect 128368 398898 128410 399134
rect 128646 398898 128688 399134
rect 128368 398866 128688 398898
rect 159088 399454 159408 399486
rect 159088 399218 159130 399454
rect 159366 399218 159408 399454
rect 159088 399134 159408 399218
rect 159088 398898 159130 399134
rect 159366 398898 159408 399134
rect 159088 398866 159408 398898
rect 189808 399454 190128 399486
rect 189808 399218 189850 399454
rect 190086 399218 190128 399454
rect 189808 399134 190128 399218
rect 189808 398898 189850 399134
rect 190086 398898 190128 399134
rect 189808 398866 190128 398898
rect 220528 399454 220848 399486
rect 220528 399218 220570 399454
rect 220806 399218 220848 399454
rect 220528 399134 220848 399218
rect 220528 398898 220570 399134
rect 220806 398898 220848 399134
rect 220528 398866 220848 398898
rect 251248 399454 251568 399486
rect 251248 399218 251290 399454
rect 251526 399218 251568 399454
rect 251248 399134 251568 399218
rect 251248 398898 251290 399134
rect 251526 398898 251568 399134
rect 251248 398866 251568 398898
rect 281968 399454 282288 399486
rect 281968 399218 282010 399454
rect 282246 399218 282288 399454
rect 281968 399134 282288 399218
rect 281968 398898 282010 399134
rect 282246 398898 282288 399134
rect 281968 398866 282288 398898
rect 312688 399454 313008 399486
rect 312688 399218 312730 399454
rect 312966 399218 313008 399454
rect 312688 399134 313008 399218
rect 312688 398898 312730 399134
rect 312966 398898 313008 399134
rect 312688 398866 313008 398898
rect 343408 399454 343728 399486
rect 343408 399218 343450 399454
rect 343686 399218 343728 399454
rect 343408 399134 343728 399218
rect 343408 398898 343450 399134
rect 343686 398898 343728 399134
rect 343408 398866 343728 398898
rect 374128 399454 374448 399486
rect 374128 399218 374170 399454
rect 374406 399218 374448 399454
rect 374128 399134 374448 399218
rect 374128 398898 374170 399134
rect 374406 398898 374448 399134
rect 374128 398866 374448 398898
rect 404848 399454 405168 399486
rect 404848 399218 404890 399454
rect 405126 399218 405168 399454
rect 404848 399134 405168 399218
rect 404848 398898 404890 399134
rect 405126 398898 405168 399134
rect 404848 398866 405168 398898
rect 435568 399454 435888 399486
rect 435568 399218 435610 399454
rect 435846 399218 435888 399454
rect 435568 399134 435888 399218
rect 435568 398898 435610 399134
rect 435846 398898 435888 399134
rect 435568 398866 435888 398898
rect 466288 399454 466608 399486
rect 466288 399218 466330 399454
rect 466566 399218 466608 399454
rect 466288 399134 466608 399218
rect 466288 398898 466330 399134
rect 466566 398898 466608 399134
rect 466288 398866 466608 398898
rect 497008 399454 497328 399486
rect 497008 399218 497050 399454
rect 497286 399218 497328 399454
rect 497008 399134 497328 399218
rect 497008 398898 497050 399134
rect 497286 398898 497328 399134
rect 497008 398866 497328 398898
rect 527728 399454 528048 399486
rect 527728 399218 527770 399454
rect 528006 399218 528048 399454
rect 527728 399134 528048 399218
rect 527728 398898 527770 399134
rect 528006 398898 528048 399134
rect 527728 398866 528048 398898
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 51568 381454 51888 381486
rect 51568 381218 51610 381454
rect 51846 381218 51888 381454
rect 51568 381134 51888 381218
rect 51568 380898 51610 381134
rect 51846 380898 51888 381134
rect 51568 380866 51888 380898
rect 82288 381454 82608 381486
rect 82288 381218 82330 381454
rect 82566 381218 82608 381454
rect 82288 381134 82608 381218
rect 82288 380898 82330 381134
rect 82566 380898 82608 381134
rect 82288 380866 82608 380898
rect 113008 381454 113328 381486
rect 113008 381218 113050 381454
rect 113286 381218 113328 381454
rect 113008 381134 113328 381218
rect 113008 380898 113050 381134
rect 113286 380898 113328 381134
rect 113008 380866 113328 380898
rect 143728 381454 144048 381486
rect 143728 381218 143770 381454
rect 144006 381218 144048 381454
rect 143728 381134 144048 381218
rect 143728 380898 143770 381134
rect 144006 380898 144048 381134
rect 143728 380866 144048 380898
rect 174448 381454 174768 381486
rect 174448 381218 174490 381454
rect 174726 381218 174768 381454
rect 174448 381134 174768 381218
rect 174448 380898 174490 381134
rect 174726 380898 174768 381134
rect 174448 380866 174768 380898
rect 205168 381454 205488 381486
rect 205168 381218 205210 381454
rect 205446 381218 205488 381454
rect 205168 381134 205488 381218
rect 205168 380898 205210 381134
rect 205446 380898 205488 381134
rect 205168 380866 205488 380898
rect 235888 381454 236208 381486
rect 235888 381218 235930 381454
rect 236166 381218 236208 381454
rect 235888 381134 236208 381218
rect 235888 380898 235930 381134
rect 236166 380898 236208 381134
rect 235888 380866 236208 380898
rect 266608 381454 266928 381486
rect 266608 381218 266650 381454
rect 266886 381218 266928 381454
rect 266608 381134 266928 381218
rect 266608 380898 266650 381134
rect 266886 380898 266928 381134
rect 266608 380866 266928 380898
rect 297328 381454 297648 381486
rect 297328 381218 297370 381454
rect 297606 381218 297648 381454
rect 297328 381134 297648 381218
rect 297328 380898 297370 381134
rect 297606 380898 297648 381134
rect 297328 380866 297648 380898
rect 328048 381454 328368 381486
rect 328048 381218 328090 381454
rect 328326 381218 328368 381454
rect 328048 381134 328368 381218
rect 328048 380898 328090 381134
rect 328326 380898 328368 381134
rect 328048 380866 328368 380898
rect 358768 381454 359088 381486
rect 358768 381218 358810 381454
rect 359046 381218 359088 381454
rect 358768 381134 359088 381218
rect 358768 380898 358810 381134
rect 359046 380898 359088 381134
rect 358768 380866 359088 380898
rect 389488 381454 389808 381486
rect 389488 381218 389530 381454
rect 389766 381218 389808 381454
rect 389488 381134 389808 381218
rect 389488 380898 389530 381134
rect 389766 380898 389808 381134
rect 389488 380866 389808 380898
rect 420208 381454 420528 381486
rect 420208 381218 420250 381454
rect 420486 381218 420528 381454
rect 420208 381134 420528 381218
rect 420208 380898 420250 381134
rect 420486 380898 420528 381134
rect 420208 380866 420528 380898
rect 450928 381454 451248 381486
rect 450928 381218 450970 381454
rect 451206 381218 451248 381454
rect 450928 381134 451248 381218
rect 450928 380898 450970 381134
rect 451206 380898 451248 381134
rect 450928 380866 451248 380898
rect 481648 381454 481968 381486
rect 481648 381218 481690 381454
rect 481926 381218 481968 381454
rect 481648 381134 481968 381218
rect 481648 380898 481690 381134
rect 481926 380898 481968 381134
rect 481648 380866 481968 380898
rect 512368 381454 512688 381486
rect 512368 381218 512410 381454
rect 512646 381218 512688 381454
rect 512368 381134 512688 381218
rect 512368 380898 512410 381134
rect 512646 380898 512688 381134
rect 512368 380866 512688 380898
rect 543088 381454 543408 381486
rect 543088 381218 543130 381454
rect 543366 381218 543408 381454
rect 543088 381134 543408 381218
rect 543088 380898 543130 381134
rect 543366 380898 543408 381134
rect 543088 380866 543408 380898
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 36208 363454 36528 363486
rect 36208 363218 36250 363454
rect 36486 363218 36528 363454
rect 36208 363134 36528 363218
rect 36208 362898 36250 363134
rect 36486 362898 36528 363134
rect 36208 362866 36528 362898
rect 66928 363454 67248 363486
rect 66928 363218 66970 363454
rect 67206 363218 67248 363454
rect 66928 363134 67248 363218
rect 66928 362898 66970 363134
rect 67206 362898 67248 363134
rect 66928 362866 67248 362898
rect 97648 363454 97968 363486
rect 97648 363218 97690 363454
rect 97926 363218 97968 363454
rect 97648 363134 97968 363218
rect 97648 362898 97690 363134
rect 97926 362898 97968 363134
rect 97648 362866 97968 362898
rect 128368 363454 128688 363486
rect 128368 363218 128410 363454
rect 128646 363218 128688 363454
rect 128368 363134 128688 363218
rect 128368 362898 128410 363134
rect 128646 362898 128688 363134
rect 128368 362866 128688 362898
rect 159088 363454 159408 363486
rect 159088 363218 159130 363454
rect 159366 363218 159408 363454
rect 159088 363134 159408 363218
rect 159088 362898 159130 363134
rect 159366 362898 159408 363134
rect 159088 362866 159408 362898
rect 189808 363454 190128 363486
rect 189808 363218 189850 363454
rect 190086 363218 190128 363454
rect 189808 363134 190128 363218
rect 189808 362898 189850 363134
rect 190086 362898 190128 363134
rect 189808 362866 190128 362898
rect 220528 363454 220848 363486
rect 220528 363218 220570 363454
rect 220806 363218 220848 363454
rect 220528 363134 220848 363218
rect 220528 362898 220570 363134
rect 220806 362898 220848 363134
rect 220528 362866 220848 362898
rect 251248 363454 251568 363486
rect 251248 363218 251290 363454
rect 251526 363218 251568 363454
rect 251248 363134 251568 363218
rect 251248 362898 251290 363134
rect 251526 362898 251568 363134
rect 251248 362866 251568 362898
rect 281968 363454 282288 363486
rect 281968 363218 282010 363454
rect 282246 363218 282288 363454
rect 281968 363134 282288 363218
rect 281968 362898 282010 363134
rect 282246 362898 282288 363134
rect 281968 362866 282288 362898
rect 312688 363454 313008 363486
rect 312688 363218 312730 363454
rect 312966 363218 313008 363454
rect 312688 363134 313008 363218
rect 312688 362898 312730 363134
rect 312966 362898 313008 363134
rect 312688 362866 313008 362898
rect 343408 363454 343728 363486
rect 343408 363218 343450 363454
rect 343686 363218 343728 363454
rect 343408 363134 343728 363218
rect 343408 362898 343450 363134
rect 343686 362898 343728 363134
rect 343408 362866 343728 362898
rect 374128 363454 374448 363486
rect 374128 363218 374170 363454
rect 374406 363218 374448 363454
rect 374128 363134 374448 363218
rect 374128 362898 374170 363134
rect 374406 362898 374448 363134
rect 374128 362866 374448 362898
rect 404848 363454 405168 363486
rect 404848 363218 404890 363454
rect 405126 363218 405168 363454
rect 404848 363134 405168 363218
rect 404848 362898 404890 363134
rect 405126 362898 405168 363134
rect 404848 362866 405168 362898
rect 435568 363454 435888 363486
rect 435568 363218 435610 363454
rect 435846 363218 435888 363454
rect 435568 363134 435888 363218
rect 435568 362898 435610 363134
rect 435846 362898 435888 363134
rect 435568 362866 435888 362898
rect 466288 363454 466608 363486
rect 466288 363218 466330 363454
rect 466566 363218 466608 363454
rect 466288 363134 466608 363218
rect 466288 362898 466330 363134
rect 466566 362898 466608 363134
rect 466288 362866 466608 362898
rect 497008 363454 497328 363486
rect 497008 363218 497050 363454
rect 497286 363218 497328 363454
rect 497008 363134 497328 363218
rect 497008 362898 497050 363134
rect 497286 362898 497328 363134
rect 497008 362866 497328 362898
rect 527728 363454 528048 363486
rect 527728 363218 527770 363454
rect 528006 363218 528048 363454
rect 527728 363134 528048 363218
rect 527728 362898 527770 363134
rect 528006 362898 528048 363134
rect 527728 362866 528048 362898
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 51568 345454 51888 345486
rect 51568 345218 51610 345454
rect 51846 345218 51888 345454
rect 51568 345134 51888 345218
rect 51568 344898 51610 345134
rect 51846 344898 51888 345134
rect 51568 344866 51888 344898
rect 82288 345454 82608 345486
rect 82288 345218 82330 345454
rect 82566 345218 82608 345454
rect 82288 345134 82608 345218
rect 82288 344898 82330 345134
rect 82566 344898 82608 345134
rect 82288 344866 82608 344898
rect 113008 345454 113328 345486
rect 113008 345218 113050 345454
rect 113286 345218 113328 345454
rect 113008 345134 113328 345218
rect 113008 344898 113050 345134
rect 113286 344898 113328 345134
rect 113008 344866 113328 344898
rect 143728 345454 144048 345486
rect 143728 345218 143770 345454
rect 144006 345218 144048 345454
rect 143728 345134 144048 345218
rect 143728 344898 143770 345134
rect 144006 344898 144048 345134
rect 143728 344866 144048 344898
rect 174448 345454 174768 345486
rect 174448 345218 174490 345454
rect 174726 345218 174768 345454
rect 174448 345134 174768 345218
rect 174448 344898 174490 345134
rect 174726 344898 174768 345134
rect 174448 344866 174768 344898
rect 205168 345454 205488 345486
rect 205168 345218 205210 345454
rect 205446 345218 205488 345454
rect 205168 345134 205488 345218
rect 205168 344898 205210 345134
rect 205446 344898 205488 345134
rect 205168 344866 205488 344898
rect 235888 345454 236208 345486
rect 235888 345218 235930 345454
rect 236166 345218 236208 345454
rect 235888 345134 236208 345218
rect 235888 344898 235930 345134
rect 236166 344898 236208 345134
rect 235888 344866 236208 344898
rect 266608 345454 266928 345486
rect 266608 345218 266650 345454
rect 266886 345218 266928 345454
rect 266608 345134 266928 345218
rect 266608 344898 266650 345134
rect 266886 344898 266928 345134
rect 266608 344866 266928 344898
rect 297328 345454 297648 345486
rect 297328 345218 297370 345454
rect 297606 345218 297648 345454
rect 297328 345134 297648 345218
rect 297328 344898 297370 345134
rect 297606 344898 297648 345134
rect 297328 344866 297648 344898
rect 328048 345454 328368 345486
rect 328048 345218 328090 345454
rect 328326 345218 328368 345454
rect 328048 345134 328368 345218
rect 328048 344898 328090 345134
rect 328326 344898 328368 345134
rect 328048 344866 328368 344898
rect 358768 345454 359088 345486
rect 358768 345218 358810 345454
rect 359046 345218 359088 345454
rect 358768 345134 359088 345218
rect 358768 344898 358810 345134
rect 359046 344898 359088 345134
rect 358768 344866 359088 344898
rect 389488 345454 389808 345486
rect 389488 345218 389530 345454
rect 389766 345218 389808 345454
rect 389488 345134 389808 345218
rect 389488 344898 389530 345134
rect 389766 344898 389808 345134
rect 389488 344866 389808 344898
rect 420208 345454 420528 345486
rect 420208 345218 420250 345454
rect 420486 345218 420528 345454
rect 420208 345134 420528 345218
rect 420208 344898 420250 345134
rect 420486 344898 420528 345134
rect 420208 344866 420528 344898
rect 450928 345454 451248 345486
rect 450928 345218 450970 345454
rect 451206 345218 451248 345454
rect 450928 345134 451248 345218
rect 450928 344898 450970 345134
rect 451206 344898 451248 345134
rect 450928 344866 451248 344898
rect 481648 345454 481968 345486
rect 481648 345218 481690 345454
rect 481926 345218 481968 345454
rect 481648 345134 481968 345218
rect 481648 344898 481690 345134
rect 481926 344898 481968 345134
rect 481648 344866 481968 344898
rect 512368 345454 512688 345486
rect 512368 345218 512410 345454
rect 512646 345218 512688 345454
rect 512368 345134 512688 345218
rect 512368 344898 512410 345134
rect 512646 344898 512688 345134
rect 512368 344866 512688 344898
rect 543088 345454 543408 345486
rect 543088 345218 543130 345454
rect 543366 345218 543408 345454
rect 543088 345134 543408 345218
rect 543088 344898 543130 345134
rect 543366 344898 543408 345134
rect 543088 344866 543408 344898
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 36208 327454 36528 327486
rect 36208 327218 36250 327454
rect 36486 327218 36528 327454
rect 36208 327134 36528 327218
rect 36208 326898 36250 327134
rect 36486 326898 36528 327134
rect 36208 326866 36528 326898
rect 66928 327454 67248 327486
rect 66928 327218 66970 327454
rect 67206 327218 67248 327454
rect 66928 327134 67248 327218
rect 66928 326898 66970 327134
rect 67206 326898 67248 327134
rect 66928 326866 67248 326898
rect 97648 327454 97968 327486
rect 97648 327218 97690 327454
rect 97926 327218 97968 327454
rect 97648 327134 97968 327218
rect 97648 326898 97690 327134
rect 97926 326898 97968 327134
rect 97648 326866 97968 326898
rect 128368 327454 128688 327486
rect 128368 327218 128410 327454
rect 128646 327218 128688 327454
rect 128368 327134 128688 327218
rect 128368 326898 128410 327134
rect 128646 326898 128688 327134
rect 128368 326866 128688 326898
rect 159088 327454 159408 327486
rect 159088 327218 159130 327454
rect 159366 327218 159408 327454
rect 159088 327134 159408 327218
rect 159088 326898 159130 327134
rect 159366 326898 159408 327134
rect 159088 326866 159408 326898
rect 189808 327454 190128 327486
rect 189808 327218 189850 327454
rect 190086 327218 190128 327454
rect 189808 327134 190128 327218
rect 189808 326898 189850 327134
rect 190086 326898 190128 327134
rect 189808 326866 190128 326898
rect 220528 327454 220848 327486
rect 220528 327218 220570 327454
rect 220806 327218 220848 327454
rect 220528 327134 220848 327218
rect 220528 326898 220570 327134
rect 220806 326898 220848 327134
rect 220528 326866 220848 326898
rect 251248 327454 251568 327486
rect 251248 327218 251290 327454
rect 251526 327218 251568 327454
rect 251248 327134 251568 327218
rect 251248 326898 251290 327134
rect 251526 326898 251568 327134
rect 251248 326866 251568 326898
rect 281968 327454 282288 327486
rect 281968 327218 282010 327454
rect 282246 327218 282288 327454
rect 281968 327134 282288 327218
rect 281968 326898 282010 327134
rect 282246 326898 282288 327134
rect 281968 326866 282288 326898
rect 312688 327454 313008 327486
rect 312688 327218 312730 327454
rect 312966 327218 313008 327454
rect 312688 327134 313008 327218
rect 312688 326898 312730 327134
rect 312966 326898 313008 327134
rect 312688 326866 313008 326898
rect 343408 327454 343728 327486
rect 343408 327218 343450 327454
rect 343686 327218 343728 327454
rect 343408 327134 343728 327218
rect 343408 326898 343450 327134
rect 343686 326898 343728 327134
rect 343408 326866 343728 326898
rect 374128 327454 374448 327486
rect 374128 327218 374170 327454
rect 374406 327218 374448 327454
rect 374128 327134 374448 327218
rect 374128 326898 374170 327134
rect 374406 326898 374448 327134
rect 374128 326866 374448 326898
rect 404848 327454 405168 327486
rect 404848 327218 404890 327454
rect 405126 327218 405168 327454
rect 404848 327134 405168 327218
rect 404848 326898 404890 327134
rect 405126 326898 405168 327134
rect 404848 326866 405168 326898
rect 435568 327454 435888 327486
rect 435568 327218 435610 327454
rect 435846 327218 435888 327454
rect 435568 327134 435888 327218
rect 435568 326898 435610 327134
rect 435846 326898 435888 327134
rect 435568 326866 435888 326898
rect 466288 327454 466608 327486
rect 466288 327218 466330 327454
rect 466566 327218 466608 327454
rect 466288 327134 466608 327218
rect 466288 326898 466330 327134
rect 466566 326898 466608 327134
rect 466288 326866 466608 326898
rect 497008 327454 497328 327486
rect 497008 327218 497050 327454
rect 497286 327218 497328 327454
rect 497008 327134 497328 327218
rect 497008 326898 497050 327134
rect 497286 326898 497328 327134
rect 497008 326866 497328 326898
rect 527728 327454 528048 327486
rect 527728 327218 527770 327454
rect 528006 327218 528048 327454
rect 527728 327134 528048 327218
rect 527728 326898 527770 327134
rect 528006 326898 528048 327134
rect 527728 326866 528048 326898
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 51568 309454 51888 309486
rect 51568 309218 51610 309454
rect 51846 309218 51888 309454
rect 51568 309134 51888 309218
rect 51568 308898 51610 309134
rect 51846 308898 51888 309134
rect 51568 308866 51888 308898
rect 82288 309454 82608 309486
rect 82288 309218 82330 309454
rect 82566 309218 82608 309454
rect 82288 309134 82608 309218
rect 82288 308898 82330 309134
rect 82566 308898 82608 309134
rect 82288 308866 82608 308898
rect 113008 309454 113328 309486
rect 113008 309218 113050 309454
rect 113286 309218 113328 309454
rect 113008 309134 113328 309218
rect 113008 308898 113050 309134
rect 113286 308898 113328 309134
rect 113008 308866 113328 308898
rect 143728 309454 144048 309486
rect 143728 309218 143770 309454
rect 144006 309218 144048 309454
rect 143728 309134 144048 309218
rect 143728 308898 143770 309134
rect 144006 308898 144048 309134
rect 143728 308866 144048 308898
rect 174448 309454 174768 309486
rect 174448 309218 174490 309454
rect 174726 309218 174768 309454
rect 174448 309134 174768 309218
rect 174448 308898 174490 309134
rect 174726 308898 174768 309134
rect 174448 308866 174768 308898
rect 205168 309454 205488 309486
rect 205168 309218 205210 309454
rect 205446 309218 205488 309454
rect 205168 309134 205488 309218
rect 205168 308898 205210 309134
rect 205446 308898 205488 309134
rect 205168 308866 205488 308898
rect 235888 309454 236208 309486
rect 235888 309218 235930 309454
rect 236166 309218 236208 309454
rect 235888 309134 236208 309218
rect 235888 308898 235930 309134
rect 236166 308898 236208 309134
rect 235888 308866 236208 308898
rect 266608 309454 266928 309486
rect 266608 309218 266650 309454
rect 266886 309218 266928 309454
rect 266608 309134 266928 309218
rect 266608 308898 266650 309134
rect 266886 308898 266928 309134
rect 266608 308866 266928 308898
rect 297328 309454 297648 309486
rect 297328 309218 297370 309454
rect 297606 309218 297648 309454
rect 297328 309134 297648 309218
rect 297328 308898 297370 309134
rect 297606 308898 297648 309134
rect 297328 308866 297648 308898
rect 328048 309454 328368 309486
rect 328048 309218 328090 309454
rect 328326 309218 328368 309454
rect 328048 309134 328368 309218
rect 328048 308898 328090 309134
rect 328326 308898 328368 309134
rect 328048 308866 328368 308898
rect 358768 309454 359088 309486
rect 358768 309218 358810 309454
rect 359046 309218 359088 309454
rect 358768 309134 359088 309218
rect 358768 308898 358810 309134
rect 359046 308898 359088 309134
rect 358768 308866 359088 308898
rect 389488 309454 389808 309486
rect 389488 309218 389530 309454
rect 389766 309218 389808 309454
rect 389488 309134 389808 309218
rect 389488 308898 389530 309134
rect 389766 308898 389808 309134
rect 389488 308866 389808 308898
rect 420208 309454 420528 309486
rect 420208 309218 420250 309454
rect 420486 309218 420528 309454
rect 420208 309134 420528 309218
rect 420208 308898 420250 309134
rect 420486 308898 420528 309134
rect 420208 308866 420528 308898
rect 450928 309454 451248 309486
rect 450928 309218 450970 309454
rect 451206 309218 451248 309454
rect 450928 309134 451248 309218
rect 450928 308898 450970 309134
rect 451206 308898 451248 309134
rect 450928 308866 451248 308898
rect 481648 309454 481968 309486
rect 481648 309218 481690 309454
rect 481926 309218 481968 309454
rect 481648 309134 481968 309218
rect 481648 308898 481690 309134
rect 481926 308898 481968 309134
rect 481648 308866 481968 308898
rect 512368 309454 512688 309486
rect 512368 309218 512410 309454
rect 512646 309218 512688 309454
rect 512368 309134 512688 309218
rect 512368 308898 512410 309134
rect 512646 308898 512688 309134
rect 512368 308866 512688 308898
rect 543088 309454 543408 309486
rect 543088 309218 543130 309454
rect 543366 309218 543408 309454
rect 543088 309134 543408 309218
rect 543088 308898 543130 309134
rect 543366 308898 543408 309134
rect 543088 308866 543408 308898
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 36208 291454 36528 291486
rect 36208 291218 36250 291454
rect 36486 291218 36528 291454
rect 36208 291134 36528 291218
rect 36208 290898 36250 291134
rect 36486 290898 36528 291134
rect 36208 290866 36528 290898
rect 66928 291454 67248 291486
rect 66928 291218 66970 291454
rect 67206 291218 67248 291454
rect 66928 291134 67248 291218
rect 66928 290898 66970 291134
rect 67206 290898 67248 291134
rect 66928 290866 67248 290898
rect 97648 291454 97968 291486
rect 97648 291218 97690 291454
rect 97926 291218 97968 291454
rect 97648 291134 97968 291218
rect 97648 290898 97690 291134
rect 97926 290898 97968 291134
rect 97648 290866 97968 290898
rect 128368 291454 128688 291486
rect 128368 291218 128410 291454
rect 128646 291218 128688 291454
rect 128368 291134 128688 291218
rect 128368 290898 128410 291134
rect 128646 290898 128688 291134
rect 128368 290866 128688 290898
rect 159088 291454 159408 291486
rect 159088 291218 159130 291454
rect 159366 291218 159408 291454
rect 159088 291134 159408 291218
rect 159088 290898 159130 291134
rect 159366 290898 159408 291134
rect 159088 290866 159408 290898
rect 189808 291454 190128 291486
rect 189808 291218 189850 291454
rect 190086 291218 190128 291454
rect 189808 291134 190128 291218
rect 189808 290898 189850 291134
rect 190086 290898 190128 291134
rect 189808 290866 190128 290898
rect 220528 291454 220848 291486
rect 220528 291218 220570 291454
rect 220806 291218 220848 291454
rect 220528 291134 220848 291218
rect 220528 290898 220570 291134
rect 220806 290898 220848 291134
rect 220528 290866 220848 290898
rect 251248 291454 251568 291486
rect 251248 291218 251290 291454
rect 251526 291218 251568 291454
rect 251248 291134 251568 291218
rect 251248 290898 251290 291134
rect 251526 290898 251568 291134
rect 251248 290866 251568 290898
rect 281968 291454 282288 291486
rect 281968 291218 282010 291454
rect 282246 291218 282288 291454
rect 281968 291134 282288 291218
rect 281968 290898 282010 291134
rect 282246 290898 282288 291134
rect 281968 290866 282288 290898
rect 312688 291454 313008 291486
rect 312688 291218 312730 291454
rect 312966 291218 313008 291454
rect 312688 291134 313008 291218
rect 312688 290898 312730 291134
rect 312966 290898 313008 291134
rect 312688 290866 313008 290898
rect 343408 291454 343728 291486
rect 343408 291218 343450 291454
rect 343686 291218 343728 291454
rect 343408 291134 343728 291218
rect 343408 290898 343450 291134
rect 343686 290898 343728 291134
rect 343408 290866 343728 290898
rect 374128 291454 374448 291486
rect 374128 291218 374170 291454
rect 374406 291218 374448 291454
rect 374128 291134 374448 291218
rect 374128 290898 374170 291134
rect 374406 290898 374448 291134
rect 374128 290866 374448 290898
rect 404848 291454 405168 291486
rect 404848 291218 404890 291454
rect 405126 291218 405168 291454
rect 404848 291134 405168 291218
rect 404848 290898 404890 291134
rect 405126 290898 405168 291134
rect 404848 290866 405168 290898
rect 435568 291454 435888 291486
rect 435568 291218 435610 291454
rect 435846 291218 435888 291454
rect 435568 291134 435888 291218
rect 435568 290898 435610 291134
rect 435846 290898 435888 291134
rect 435568 290866 435888 290898
rect 466288 291454 466608 291486
rect 466288 291218 466330 291454
rect 466566 291218 466608 291454
rect 466288 291134 466608 291218
rect 466288 290898 466330 291134
rect 466566 290898 466608 291134
rect 466288 290866 466608 290898
rect 497008 291454 497328 291486
rect 497008 291218 497050 291454
rect 497286 291218 497328 291454
rect 497008 291134 497328 291218
rect 497008 290898 497050 291134
rect 497286 290898 497328 291134
rect 497008 290866 497328 290898
rect 527728 291454 528048 291486
rect 527728 291218 527770 291454
rect 528006 291218 528048 291454
rect 527728 291134 528048 291218
rect 527728 290898 527770 291134
rect 528006 290898 528048 291134
rect 527728 290866 528048 290898
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 51568 273454 51888 273486
rect 51568 273218 51610 273454
rect 51846 273218 51888 273454
rect 51568 273134 51888 273218
rect 51568 272898 51610 273134
rect 51846 272898 51888 273134
rect 51568 272866 51888 272898
rect 82288 273454 82608 273486
rect 82288 273218 82330 273454
rect 82566 273218 82608 273454
rect 82288 273134 82608 273218
rect 82288 272898 82330 273134
rect 82566 272898 82608 273134
rect 82288 272866 82608 272898
rect 113008 273454 113328 273486
rect 113008 273218 113050 273454
rect 113286 273218 113328 273454
rect 113008 273134 113328 273218
rect 113008 272898 113050 273134
rect 113286 272898 113328 273134
rect 113008 272866 113328 272898
rect 143728 273454 144048 273486
rect 143728 273218 143770 273454
rect 144006 273218 144048 273454
rect 143728 273134 144048 273218
rect 143728 272898 143770 273134
rect 144006 272898 144048 273134
rect 143728 272866 144048 272898
rect 174448 273454 174768 273486
rect 174448 273218 174490 273454
rect 174726 273218 174768 273454
rect 174448 273134 174768 273218
rect 174448 272898 174490 273134
rect 174726 272898 174768 273134
rect 174448 272866 174768 272898
rect 205168 273454 205488 273486
rect 205168 273218 205210 273454
rect 205446 273218 205488 273454
rect 205168 273134 205488 273218
rect 205168 272898 205210 273134
rect 205446 272898 205488 273134
rect 205168 272866 205488 272898
rect 235888 273454 236208 273486
rect 235888 273218 235930 273454
rect 236166 273218 236208 273454
rect 235888 273134 236208 273218
rect 235888 272898 235930 273134
rect 236166 272898 236208 273134
rect 235888 272866 236208 272898
rect 266608 273454 266928 273486
rect 266608 273218 266650 273454
rect 266886 273218 266928 273454
rect 266608 273134 266928 273218
rect 266608 272898 266650 273134
rect 266886 272898 266928 273134
rect 266608 272866 266928 272898
rect 297328 273454 297648 273486
rect 297328 273218 297370 273454
rect 297606 273218 297648 273454
rect 297328 273134 297648 273218
rect 297328 272898 297370 273134
rect 297606 272898 297648 273134
rect 297328 272866 297648 272898
rect 328048 273454 328368 273486
rect 328048 273218 328090 273454
rect 328326 273218 328368 273454
rect 328048 273134 328368 273218
rect 328048 272898 328090 273134
rect 328326 272898 328368 273134
rect 328048 272866 328368 272898
rect 358768 273454 359088 273486
rect 358768 273218 358810 273454
rect 359046 273218 359088 273454
rect 358768 273134 359088 273218
rect 358768 272898 358810 273134
rect 359046 272898 359088 273134
rect 358768 272866 359088 272898
rect 389488 273454 389808 273486
rect 389488 273218 389530 273454
rect 389766 273218 389808 273454
rect 389488 273134 389808 273218
rect 389488 272898 389530 273134
rect 389766 272898 389808 273134
rect 389488 272866 389808 272898
rect 420208 273454 420528 273486
rect 420208 273218 420250 273454
rect 420486 273218 420528 273454
rect 420208 273134 420528 273218
rect 420208 272898 420250 273134
rect 420486 272898 420528 273134
rect 420208 272866 420528 272898
rect 450928 273454 451248 273486
rect 450928 273218 450970 273454
rect 451206 273218 451248 273454
rect 450928 273134 451248 273218
rect 450928 272898 450970 273134
rect 451206 272898 451248 273134
rect 450928 272866 451248 272898
rect 481648 273454 481968 273486
rect 481648 273218 481690 273454
rect 481926 273218 481968 273454
rect 481648 273134 481968 273218
rect 481648 272898 481690 273134
rect 481926 272898 481968 273134
rect 481648 272866 481968 272898
rect 512368 273454 512688 273486
rect 512368 273218 512410 273454
rect 512646 273218 512688 273454
rect 512368 273134 512688 273218
rect 512368 272898 512410 273134
rect 512646 272898 512688 273134
rect 512368 272866 512688 272898
rect 543088 273454 543408 273486
rect 543088 273218 543130 273454
rect 543366 273218 543408 273454
rect 543088 273134 543408 273218
rect 543088 272898 543130 273134
rect 543366 272898 543408 273134
rect 543088 272866 543408 272898
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 36208 255454 36528 255486
rect 36208 255218 36250 255454
rect 36486 255218 36528 255454
rect 36208 255134 36528 255218
rect 36208 254898 36250 255134
rect 36486 254898 36528 255134
rect 36208 254866 36528 254898
rect 66928 255454 67248 255486
rect 66928 255218 66970 255454
rect 67206 255218 67248 255454
rect 66928 255134 67248 255218
rect 66928 254898 66970 255134
rect 67206 254898 67248 255134
rect 66928 254866 67248 254898
rect 97648 255454 97968 255486
rect 97648 255218 97690 255454
rect 97926 255218 97968 255454
rect 97648 255134 97968 255218
rect 97648 254898 97690 255134
rect 97926 254898 97968 255134
rect 97648 254866 97968 254898
rect 128368 255454 128688 255486
rect 128368 255218 128410 255454
rect 128646 255218 128688 255454
rect 128368 255134 128688 255218
rect 128368 254898 128410 255134
rect 128646 254898 128688 255134
rect 128368 254866 128688 254898
rect 159088 255454 159408 255486
rect 159088 255218 159130 255454
rect 159366 255218 159408 255454
rect 159088 255134 159408 255218
rect 159088 254898 159130 255134
rect 159366 254898 159408 255134
rect 159088 254866 159408 254898
rect 189808 255454 190128 255486
rect 189808 255218 189850 255454
rect 190086 255218 190128 255454
rect 189808 255134 190128 255218
rect 189808 254898 189850 255134
rect 190086 254898 190128 255134
rect 189808 254866 190128 254898
rect 220528 255454 220848 255486
rect 220528 255218 220570 255454
rect 220806 255218 220848 255454
rect 220528 255134 220848 255218
rect 220528 254898 220570 255134
rect 220806 254898 220848 255134
rect 220528 254866 220848 254898
rect 251248 255454 251568 255486
rect 251248 255218 251290 255454
rect 251526 255218 251568 255454
rect 251248 255134 251568 255218
rect 251248 254898 251290 255134
rect 251526 254898 251568 255134
rect 251248 254866 251568 254898
rect 281968 255454 282288 255486
rect 281968 255218 282010 255454
rect 282246 255218 282288 255454
rect 281968 255134 282288 255218
rect 281968 254898 282010 255134
rect 282246 254898 282288 255134
rect 281968 254866 282288 254898
rect 312688 255454 313008 255486
rect 312688 255218 312730 255454
rect 312966 255218 313008 255454
rect 312688 255134 313008 255218
rect 312688 254898 312730 255134
rect 312966 254898 313008 255134
rect 312688 254866 313008 254898
rect 343408 255454 343728 255486
rect 343408 255218 343450 255454
rect 343686 255218 343728 255454
rect 343408 255134 343728 255218
rect 343408 254898 343450 255134
rect 343686 254898 343728 255134
rect 343408 254866 343728 254898
rect 374128 255454 374448 255486
rect 374128 255218 374170 255454
rect 374406 255218 374448 255454
rect 374128 255134 374448 255218
rect 374128 254898 374170 255134
rect 374406 254898 374448 255134
rect 374128 254866 374448 254898
rect 404848 255454 405168 255486
rect 404848 255218 404890 255454
rect 405126 255218 405168 255454
rect 404848 255134 405168 255218
rect 404848 254898 404890 255134
rect 405126 254898 405168 255134
rect 404848 254866 405168 254898
rect 435568 255454 435888 255486
rect 435568 255218 435610 255454
rect 435846 255218 435888 255454
rect 435568 255134 435888 255218
rect 435568 254898 435610 255134
rect 435846 254898 435888 255134
rect 435568 254866 435888 254898
rect 466288 255454 466608 255486
rect 466288 255218 466330 255454
rect 466566 255218 466608 255454
rect 466288 255134 466608 255218
rect 466288 254898 466330 255134
rect 466566 254898 466608 255134
rect 466288 254866 466608 254898
rect 497008 255454 497328 255486
rect 497008 255218 497050 255454
rect 497286 255218 497328 255454
rect 497008 255134 497328 255218
rect 497008 254898 497050 255134
rect 497286 254898 497328 255134
rect 497008 254866 497328 254898
rect 527728 255454 528048 255486
rect 527728 255218 527770 255454
rect 528006 255218 528048 255454
rect 527728 255134 528048 255218
rect 527728 254898 527770 255134
rect 528006 254898 528048 255134
rect 527728 254866 528048 254898
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 51568 237454 51888 237486
rect 51568 237218 51610 237454
rect 51846 237218 51888 237454
rect 51568 237134 51888 237218
rect 51568 236898 51610 237134
rect 51846 236898 51888 237134
rect 51568 236866 51888 236898
rect 82288 237454 82608 237486
rect 82288 237218 82330 237454
rect 82566 237218 82608 237454
rect 82288 237134 82608 237218
rect 82288 236898 82330 237134
rect 82566 236898 82608 237134
rect 82288 236866 82608 236898
rect 113008 237454 113328 237486
rect 113008 237218 113050 237454
rect 113286 237218 113328 237454
rect 113008 237134 113328 237218
rect 113008 236898 113050 237134
rect 113286 236898 113328 237134
rect 113008 236866 113328 236898
rect 143728 237454 144048 237486
rect 143728 237218 143770 237454
rect 144006 237218 144048 237454
rect 143728 237134 144048 237218
rect 143728 236898 143770 237134
rect 144006 236898 144048 237134
rect 143728 236866 144048 236898
rect 174448 237454 174768 237486
rect 174448 237218 174490 237454
rect 174726 237218 174768 237454
rect 174448 237134 174768 237218
rect 174448 236898 174490 237134
rect 174726 236898 174768 237134
rect 174448 236866 174768 236898
rect 205168 237454 205488 237486
rect 205168 237218 205210 237454
rect 205446 237218 205488 237454
rect 205168 237134 205488 237218
rect 205168 236898 205210 237134
rect 205446 236898 205488 237134
rect 205168 236866 205488 236898
rect 235888 237454 236208 237486
rect 235888 237218 235930 237454
rect 236166 237218 236208 237454
rect 235888 237134 236208 237218
rect 235888 236898 235930 237134
rect 236166 236898 236208 237134
rect 235888 236866 236208 236898
rect 266608 237454 266928 237486
rect 266608 237218 266650 237454
rect 266886 237218 266928 237454
rect 266608 237134 266928 237218
rect 266608 236898 266650 237134
rect 266886 236898 266928 237134
rect 266608 236866 266928 236898
rect 297328 237454 297648 237486
rect 297328 237218 297370 237454
rect 297606 237218 297648 237454
rect 297328 237134 297648 237218
rect 297328 236898 297370 237134
rect 297606 236898 297648 237134
rect 297328 236866 297648 236898
rect 328048 237454 328368 237486
rect 328048 237218 328090 237454
rect 328326 237218 328368 237454
rect 328048 237134 328368 237218
rect 328048 236898 328090 237134
rect 328326 236898 328368 237134
rect 328048 236866 328368 236898
rect 358768 237454 359088 237486
rect 358768 237218 358810 237454
rect 359046 237218 359088 237454
rect 358768 237134 359088 237218
rect 358768 236898 358810 237134
rect 359046 236898 359088 237134
rect 358768 236866 359088 236898
rect 389488 237454 389808 237486
rect 389488 237218 389530 237454
rect 389766 237218 389808 237454
rect 389488 237134 389808 237218
rect 389488 236898 389530 237134
rect 389766 236898 389808 237134
rect 389488 236866 389808 236898
rect 420208 237454 420528 237486
rect 420208 237218 420250 237454
rect 420486 237218 420528 237454
rect 420208 237134 420528 237218
rect 420208 236898 420250 237134
rect 420486 236898 420528 237134
rect 420208 236866 420528 236898
rect 450928 237454 451248 237486
rect 450928 237218 450970 237454
rect 451206 237218 451248 237454
rect 450928 237134 451248 237218
rect 450928 236898 450970 237134
rect 451206 236898 451248 237134
rect 450928 236866 451248 236898
rect 481648 237454 481968 237486
rect 481648 237218 481690 237454
rect 481926 237218 481968 237454
rect 481648 237134 481968 237218
rect 481648 236898 481690 237134
rect 481926 236898 481968 237134
rect 481648 236866 481968 236898
rect 512368 237454 512688 237486
rect 512368 237218 512410 237454
rect 512646 237218 512688 237454
rect 512368 237134 512688 237218
rect 512368 236898 512410 237134
rect 512646 236898 512688 237134
rect 512368 236866 512688 236898
rect 543088 237454 543408 237486
rect 543088 237218 543130 237454
rect 543366 237218 543408 237454
rect 543088 237134 543408 237218
rect 543088 236898 543130 237134
rect 543366 236898 543408 237134
rect 543088 236866 543408 236898
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 36208 219454 36528 219486
rect 36208 219218 36250 219454
rect 36486 219218 36528 219454
rect 36208 219134 36528 219218
rect 36208 218898 36250 219134
rect 36486 218898 36528 219134
rect 36208 218866 36528 218898
rect 66928 219454 67248 219486
rect 66928 219218 66970 219454
rect 67206 219218 67248 219454
rect 66928 219134 67248 219218
rect 66928 218898 66970 219134
rect 67206 218898 67248 219134
rect 66928 218866 67248 218898
rect 97648 219454 97968 219486
rect 97648 219218 97690 219454
rect 97926 219218 97968 219454
rect 97648 219134 97968 219218
rect 97648 218898 97690 219134
rect 97926 218898 97968 219134
rect 97648 218866 97968 218898
rect 128368 219454 128688 219486
rect 128368 219218 128410 219454
rect 128646 219218 128688 219454
rect 128368 219134 128688 219218
rect 128368 218898 128410 219134
rect 128646 218898 128688 219134
rect 128368 218866 128688 218898
rect 159088 219454 159408 219486
rect 159088 219218 159130 219454
rect 159366 219218 159408 219454
rect 159088 219134 159408 219218
rect 159088 218898 159130 219134
rect 159366 218898 159408 219134
rect 159088 218866 159408 218898
rect 189808 219454 190128 219486
rect 189808 219218 189850 219454
rect 190086 219218 190128 219454
rect 189808 219134 190128 219218
rect 189808 218898 189850 219134
rect 190086 218898 190128 219134
rect 189808 218866 190128 218898
rect 220528 219454 220848 219486
rect 220528 219218 220570 219454
rect 220806 219218 220848 219454
rect 220528 219134 220848 219218
rect 220528 218898 220570 219134
rect 220806 218898 220848 219134
rect 220528 218866 220848 218898
rect 251248 219454 251568 219486
rect 251248 219218 251290 219454
rect 251526 219218 251568 219454
rect 251248 219134 251568 219218
rect 251248 218898 251290 219134
rect 251526 218898 251568 219134
rect 251248 218866 251568 218898
rect 281968 219454 282288 219486
rect 281968 219218 282010 219454
rect 282246 219218 282288 219454
rect 281968 219134 282288 219218
rect 281968 218898 282010 219134
rect 282246 218898 282288 219134
rect 281968 218866 282288 218898
rect 312688 219454 313008 219486
rect 312688 219218 312730 219454
rect 312966 219218 313008 219454
rect 312688 219134 313008 219218
rect 312688 218898 312730 219134
rect 312966 218898 313008 219134
rect 312688 218866 313008 218898
rect 343408 219454 343728 219486
rect 343408 219218 343450 219454
rect 343686 219218 343728 219454
rect 343408 219134 343728 219218
rect 343408 218898 343450 219134
rect 343686 218898 343728 219134
rect 343408 218866 343728 218898
rect 374128 219454 374448 219486
rect 374128 219218 374170 219454
rect 374406 219218 374448 219454
rect 374128 219134 374448 219218
rect 374128 218898 374170 219134
rect 374406 218898 374448 219134
rect 374128 218866 374448 218898
rect 404848 219454 405168 219486
rect 404848 219218 404890 219454
rect 405126 219218 405168 219454
rect 404848 219134 405168 219218
rect 404848 218898 404890 219134
rect 405126 218898 405168 219134
rect 404848 218866 405168 218898
rect 435568 219454 435888 219486
rect 435568 219218 435610 219454
rect 435846 219218 435888 219454
rect 435568 219134 435888 219218
rect 435568 218898 435610 219134
rect 435846 218898 435888 219134
rect 435568 218866 435888 218898
rect 466288 219454 466608 219486
rect 466288 219218 466330 219454
rect 466566 219218 466608 219454
rect 466288 219134 466608 219218
rect 466288 218898 466330 219134
rect 466566 218898 466608 219134
rect 466288 218866 466608 218898
rect 497008 219454 497328 219486
rect 497008 219218 497050 219454
rect 497286 219218 497328 219454
rect 497008 219134 497328 219218
rect 497008 218898 497050 219134
rect 497286 218898 497328 219134
rect 497008 218866 497328 218898
rect 527728 219454 528048 219486
rect 527728 219218 527770 219454
rect 528006 219218 528048 219454
rect 527728 219134 528048 219218
rect 527728 218898 527770 219134
rect 528006 218898 528048 219134
rect 527728 218866 528048 218898
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 51568 201454 51888 201486
rect 51568 201218 51610 201454
rect 51846 201218 51888 201454
rect 51568 201134 51888 201218
rect 51568 200898 51610 201134
rect 51846 200898 51888 201134
rect 51568 200866 51888 200898
rect 82288 201454 82608 201486
rect 82288 201218 82330 201454
rect 82566 201218 82608 201454
rect 82288 201134 82608 201218
rect 82288 200898 82330 201134
rect 82566 200898 82608 201134
rect 82288 200866 82608 200898
rect 113008 201454 113328 201486
rect 113008 201218 113050 201454
rect 113286 201218 113328 201454
rect 113008 201134 113328 201218
rect 113008 200898 113050 201134
rect 113286 200898 113328 201134
rect 113008 200866 113328 200898
rect 143728 201454 144048 201486
rect 143728 201218 143770 201454
rect 144006 201218 144048 201454
rect 143728 201134 144048 201218
rect 143728 200898 143770 201134
rect 144006 200898 144048 201134
rect 143728 200866 144048 200898
rect 174448 201454 174768 201486
rect 174448 201218 174490 201454
rect 174726 201218 174768 201454
rect 174448 201134 174768 201218
rect 174448 200898 174490 201134
rect 174726 200898 174768 201134
rect 174448 200866 174768 200898
rect 205168 201454 205488 201486
rect 205168 201218 205210 201454
rect 205446 201218 205488 201454
rect 205168 201134 205488 201218
rect 205168 200898 205210 201134
rect 205446 200898 205488 201134
rect 205168 200866 205488 200898
rect 235888 201454 236208 201486
rect 235888 201218 235930 201454
rect 236166 201218 236208 201454
rect 235888 201134 236208 201218
rect 235888 200898 235930 201134
rect 236166 200898 236208 201134
rect 235888 200866 236208 200898
rect 266608 201454 266928 201486
rect 266608 201218 266650 201454
rect 266886 201218 266928 201454
rect 266608 201134 266928 201218
rect 266608 200898 266650 201134
rect 266886 200898 266928 201134
rect 266608 200866 266928 200898
rect 297328 201454 297648 201486
rect 297328 201218 297370 201454
rect 297606 201218 297648 201454
rect 297328 201134 297648 201218
rect 297328 200898 297370 201134
rect 297606 200898 297648 201134
rect 297328 200866 297648 200898
rect 328048 201454 328368 201486
rect 328048 201218 328090 201454
rect 328326 201218 328368 201454
rect 328048 201134 328368 201218
rect 328048 200898 328090 201134
rect 328326 200898 328368 201134
rect 328048 200866 328368 200898
rect 358768 201454 359088 201486
rect 358768 201218 358810 201454
rect 359046 201218 359088 201454
rect 358768 201134 359088 201218
rect 358768 200898 358810 201134
rect 359046 200898 359088 201134
rect 358768 200866 359088 200898
rect 389488 201454 389808 201486
rect 389488 201218 389530 201454
rect 389766 201218 389808 201454
rect 389488 201134 389808 201218
rect 389488 200898 389530 201134
rect 389766 200898 389808 201134
rect 389488 200866 389808 200898
rect 420208 201454 420528 201486
rect 420208 201218 420250 201454
rect 420486 201218 420528 201454
rect 420208 201134 420528 201218
rect 420208 200898 420250 201134
rect 420486 200898 420528 201134
rect 420208 200866 420528 200898
rect 450928 201454 451248 201486
rect 450928 201218 450970 201454
rect 451206 201218 451248 201454
rect 450928 201134 451248 201218
rect 450928 200898 450970 201134
rect 451206 200898 451248 201134
rect 450928 200866 451248 200898
rect 481648 201454 481968 201486
rect 481648 201218 481690 201454
rect 481926 201218 481968 201454
rect 481648 201134 481968 201218
rect 481648 200898 481690 201134
rect 481926 200898 481968 201134
rect 481648 200866 481968 200898
rect 512368 201454 512688 201486
rect 512368 201218 512410 201454
rect 512646 201218 512688 201454
rect 512368 201134 512688 201218
rect 512368 200898 512410 201134
rect 512646 200898 512688 201134
rect 512368 200866 512688 200898
rect 543088 201454 543408 201486
rect 543088 201218 543130 201454
rect 543366 201218 543408 201454
rect 543088 201134 543408 201218
rect 543088 200898 543130 201134
rect 543366 200898 543408 201134
rect 543088 200866 543408 200898
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 36208 183454 36528 183486
rect 36208 183218 36250 183454
rect 36486 183218 36528 183454
rect 36208 183134 36528 183218
rect 36208 182898 36250 183134
rect 36486 182898 36528 183134
rect 36208 182866 36528 182898
rect 66928 183454 67248 183486
rect 66928 183218 66970 183454
rect 67206 183218 67248 183454
rect 66928 183134 67248 183218
rect 66928 182898 66970 183134
rect 67206 182898 67248 183134
rect 66928 182866 67248 182898
rect 97648 183454 97968 183486
rect 97648 183218 97690 183454
rect 97926 183218 97968 183454
rect 97648 183134 97968 183218
rect 97648 182898 97690 183134
rect 97926 182898 97968 183134
rect 97648 182866 97968 182898
rect 128368 183454 128688 183486
rect 128368 183218 128410 183454
rect 128646 183218 128688 183454
rect 128368 183134 128688 183218
rect 128368 182898 128410 183134
rect 128646 182898 128688 183134
rect 128368 182866 128688 182898
rect 159088 183454 159408 183486
rect 159088 183218 159130 183454
rect 159366 183218 159408 183454
rect 159088 183134 159408 183218
rect 159088 182898 159130 183134
rect 159366 182898 159408 183134
rect 159088 182866 159408 182898
rect 189808 183454 190128 183486
rect 189808 183218 189850 183454
rect 190086 183218 190128 183454
rect 189808 183134 190128 183218
rect 189808 182898 189850 183134
rect 190086 182898 190128 183134
rect 189808 182866 190128 182898
rect 220528 183454 220848 183486
rect 220528 183218 220570 183454
rect 220806 183218 220848 183454
rect 220528 183134 220848 183218
rect 220528 182898 220570 183134
rect 220806 182898 220848 183134
rect 220528 182866 220848 182898
rect 251248 183454 251568 183486
rect 251248 183218 251290 183454
rect 251526 183218 251568 183454
rect 251248 183134 251568 183218
rect 251248 182898 251290 183134
rect 251526 182898 251568 183134
rect 251248 182866 251568 182898
rect 281968 183454 282288 183486
rect 281968 183218 282010 183454
rect 282246 183218 282288 183454
rect 281968 183134 282288 183218
rect 281968 182898 282010 183134
rect 282246 182898 282288 183134
rect 281968 182866 282288 182898
rect 312688 183454 313008 183486
rect 312688 183218 312730 183454
rect 312966 183218 313008 183454
rect 312688 183134 313008 183218
rect 312688 182898 312730 183134
rect 312966 182898 313008 183134
rect 312688 182866 313008 182898
rect 343408 183454 343728 183486
rect 343408 183218 343450 183454
rect 343686 183218 343728 183454
rect 343408 183134 343728 183218
rect 343408 182898 343450 183134
rect 343686 182898 343728 183134
rect 343408 182866 343728 182898
rect 374128 183454 374448 183486
rect 374128 183218 374170 183454
rect 374406 183218 374448 183454
rect 374128 183134 374448 183218
rect 374128 182898 374170 183134
rect 374406 182898 374448 183134
rect 374128 182866 374448 182898
rect 404848 183454 405168 183486
rect 404848 183218 404890 183454
rect 405126 183218 405168 183454
rect 404848 183134 405168 183218
rect 404848 182898 404890 183134
rect 405126 182898 405168 183134
rect 404848 182866 405168 182898
rect 435568 183454 435888 183486
rect 435568 183218 435610 183454
rect 435846 183218 435888 183454
rect 435568 183134 435888 183218
rect 435568 182898 435610 183134
rect 435846 182898 435888 183134
rect 435568 182866 435888 182898
rect 466288 183454 466608 183486
rect 466288 183218 466330 183454
rect 466566 183218 466608 183454
rect 466288 183134 466608 183218
rect 466288 182898 466330 183134
rect 466566 182898 466608 183134
rect 466288 182866 466608 182898
rect 497008 183454 497328 183486
rect 497008 183218 497050 183454
rect 497286 183218 497328 183454
rect 497008 183134 497328 183218
rect 497008 182898 497050 183134
rect 497286 182898 497328 183134
rect 497008 182866 497328 182898
rect 527728 183454 528048 183486
rect 527728 183218 527770 183454
rect 528006 183218 528048 183454
rect 527728 183134 528048 183218
rect 527728 182898 527770 183134
rect 528006 182898 528048 183134
rect 527728 182866 528048 182898
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 51568 165454 51888 165486
rect 51568 165218 51610 165454
rect 51846 165218 51888 165454
rect 51568 165134 51888 165218
rect 51568 164898 51610 165134
rect 51846 164898 51888 165134
rect 51568 164866 51888 164898
rect 82288 165454 82608 165486
rect 82288 165218 82330 165454
rect 82566 165218 82608 165454
rect 82288 165134 82608 165218
rect 82288 164898 82330 165134
rect 82566 164898 82608 165134
rect 82288 164866 82608 164898
rect 113008 165454 113328 165486
rect 113008 165218 113050 165454
rect 113286 165218 113328 165454
rect 113008 165134 113328 165218
rect 113008 164898 113050 165134
rect 113286 164898 113328 165134
rect 113008 164866 113328 164898
rect 143728 165454 144048 165486
rect 143728 165218 143770 165454
rect 144006 165218 144048 165454
rect 143728 165134 144048 165218
rect 143728 164898 143770 165134
rect 144006 164898 144048 165134
rect 143728 164866 144048 164898
rect 174448 165454 174768 165486
rect 174448 165218 174490 165454
rect 174726 165218 174768 165454
rect 174448 165134 174768 165218
rect 174448 164898 174490 165134
rect 174726 164898 174768 165134
rect 174448 164866 174768 164898
rect 205168 165454 205488 165486
rect 205168 165218 205210 165454
rect 205446 165218 205488 165454
rect 205168 165134 205488 165218
rect 205168 164898 205210 165134
rect 205446 164898 205488 165134
rect 205168 164866 205488 164898
rect 235888 165454 236208 165486
rect 235888 165218 235930 165454
rect 236166 165218 236208 165454
rect 235888 165134 236208 165218
rect 235888 164898 235930 165134
rect 236166 164898 236208 165134
rect 235888 164866 236208 164898
rect 266608 165454 266928 165486
rect 266608 165218 266650 165454
rect 266886 165218 266928 165454
rect 266608 165134 266928 165218
rect 266608 164898 266650 165134
rect 266886 164898 266928 165134
rect 266608 164866 266928 164898
rect 297328 165454 297648 165486
rect 297328 165218 297370 165454
rect 297606 165218 297648 165454
rect 297328 165134 297648 165218
rect 297328 164898 297370 165134
rect 297606 164898 297648 165134
rect 297328 164866 297648 164898
rect 328048 165454 328368 165486
rect 328048 165218 328090 165454
rect 328326 165218 328368 165454
rect 328048 165134 328368 165218
rect 328048 164898 328090 165134
rect 328326 164898 328368 165134
rect 328048 164866 328368 164898
rect 358768 165454 359088 165486
rect 358768 165218 358810 165454
rect 359046 165218 359088 165454
rect 358768 165134 359088 165218
rect 358768 164898 358810 165134
rect 359046 164898 359088 165134
rect 358768 164866 359088 164898
rect 389488 165454 389808 165486
rect 389488 165218 389530 165454
rect 389766 165218 389808 165454
rect 389488 165134 389808 165218
rect 389488 164898 389530 165134
rect 389766 164898 389808 165134
rect 389488 164866 389808 164898
rect 420208 165454 420528 165486
rect 420208 165218 420250 165454
rect 420486 165218 420528 165454
rect 420208 165134 420528 165218
rect 420208 164898 420250 165134
rect 420486 164898 420528 165134
rect 420208 164866 420528 164898
rect 450928 165454 451248 165486
rect 450928 165218 450970 165454
rect 451206 165218 451248 165454
rect 450928 165134 451248 165218
rect 450928 164898 450970 165134
rect 451206 164898 451248 165134
rect 450928 164866 451248 164898
rect 481648 165454 481968 165486
rect 481648 165218 481690 165454
rect 481926 165218 481968 165454
rect 481648 165134 481968 165218
rect 481648 164898 481690 165134
rect 481926 164898 481968 165134
rect 481648 164866 481968 164898
rect 512368 165454 512688 165486
rect 512368 165218 512410 165454
rect 512646 165218 512688 165454
rect 512368 165134 512688 165218
rect 512368 164898 512410 165134
rect 512646 164898 512688 165134
rect 512368 164866 512688 164898
rect 543088 165454 543408 165486
rect 543088 165218 543130 165454
rect 543366 165218 543408 165454
rect 543088 165134 543408 165218
rect 543088 164898 543130 165134
rect 543366 164898 543408 165134
rect 543088 164866 543408 164898
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 36208 147454 36528 147486
rect 36208 147218 36250 147454
rect 36486 147218 36528 147454
rect 36208 147134 36528 147218
rect 36208 146898 36250 147134
rect 36486 146898 36528 147134
rect 36208 146866 36528 146898
rect 66928 147454 67248 147486
rect 66928 147218 66970 147454
rect 67206 147218 67248 147454
rect 66928 147134 67248 147218
rect 66928 146898 66970 147134
rect 67206 146898 67248 147134
rect 66928 146866 67248 146898
rect 97648 147454 97968 147486
rect 97648 147218 97690 147454
rect 97926 147218 97968 147454
rect 97648 147134 97968 147218
rect 97648 146898 97690 147134
rect 97926 146898 97968 147134
rect 97648 146866 97968 146898
rect 128368 147454 128688 147486
rect 128368 147218 128410 147454
rect 128646 147218 128688 147454
rect 128368 147134 128688 147218
rect 128368 146898 128410 147134
rect 128646 146898 128688 147134
rect 128368 146866 128688 146898
rect 159088 147454 159408 147486
rect 159088 147218 159130 147454
rect 159366 147218 159408 147454
rect 159088 147134 159408 147218
rect 159088 146898 159130 147134
rect 159366 146898 159408 147134
rect 159088 146866 159408 146898
rect 189808 147454 190128 147486
rect 189808 147218 189850 147454
rect 190086 147218 190128 147454
rect 189808 147134 190128 147218
rect 189808 146898 189850 147134
rect 190086 146898 190128 147134
rect 189808 146866 190128 146898
rect 220528 147454 220848 147486
rect 220528 147218 220570 147454
rect 220806 147218 220848 147454
rect 220528 147134 220848 147218
rect 220528 146898 220570 147134
rect 220806 146898 220848 147134
rect 220528 146866 220848 146898
rect 251248 147454 251568 147486
rect 251248 147218 251290 147454
rect 251526 147218 251568 147454
rect 251248 147134 251568 147218
rect 251248 146898 251290 147134
rect 251526 146898 251568 147134
rect 251248 146866 251568 146898
rect 281968 147454 282288 147486
rect 281968 147218 282010 147454
rect 282246 147218 282288 147454
rect 281968 147134 282288 147218
rect 281968 146898 282010 147134
rect 282246 146898 282288 147134
rect 281968 146866 282288 146898
rect 312688 147454 313008 147486
rect 312688 147218 312730 147454
rect 312966 147218 313008 147454
rect 312688 147134 313008 147218
rect 312688 146898 312730 147134
rect 312966 146898 313008 147134
rect 312688 146866 313008 146898
rect 343408 147454 343728 147486
rect 343408 147218 343450 147454
rect 343686 147218 343728 147454
rect 343408 147134 343728 147218
rect 343408 146898 343450 147134
rect 343686 146898 343728 147134
rect 343408 146866 343728 146898
rect 374128 147454 374448 147486
rect 374128 147218 374170 147454
rect 374406 147218 374448 147454
rect 374128 147134 374448 147218
rect 374128 146898 374170 147134
rect 374406 146898 374448 147134
rect 374128 146866 374448 146898
rect 404848 147454 405168 147486
rect 404848 147218 404890 147454
rect 405126 147218 405168 147454
rect 404848 147134 405168 147218
rect 404848 146898 404890 147134
rect 405126 146898 405168 147134
rect 404848 146866 405168 146898
rect 435568 147454 435888 147486
rect 435568 147218 435610 147454
rect 435846 147218 435888 147454
rect 435568 147134 435888 147218
rect 435568 146898 435610 147134
rect 435846 146898 435888 147134
rect 435568 146866 435888 146898
rect 466288 147454 466608 147486
rect 466288 147218 466330 147454
rect 466566 147218 466608 147454
rect 466288 147134 466608 147218
rect 466288 146898 466330 147134
rect 466566 146898 466608 147134
rect 466288 146866 466608 146898
rect 497008 147454 497328 147486
rect 497008 147218 497050 147454
rect 497286 147218 497328 147454
rect 497008 147134 497328 147218
rect 497008 146898 497050 147134
rect 497286 146898 497328 147134
rect 497008 146866 497328 146898
rect 527728 147454 528048 147486
rect 527728 147218 527770 147454
rect 528006 147218 528048 147454
rect 527728 147134 528048 147218
rect 527728 146898 527770 147134
rect 528006 146898 528048 147134
rect 527728 146866 528048 146898
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 51568 129454 51888 129486
rect 51568 129218 51610 129454
rect 51846 129218 51888 129454
rect 51568 129134 51888 129218
rect 51568 128898 51610 129134
rect 51846 128898 51888 129134
rect 51568 128866 51888 128898
rect 82288 129454 82608 129486
rect 82288 129218 82330 129454
rect 82566 129218 82608 129454
rect 82288 129134 82608 129218
rect 82288 128898 82330 129134
rect 82566 128898 82608 129134
rect 82288 128866 82608 128898
rect 113008 129454 113328 129486
rect 113008 129218 113050 129454
rect 113286 129218 113328 129454
rect 113008 129134 113328 129218
rect 113008 128898 113050 129134
rect 113286 128898 113328 129134
rect 113008 128866 113328 128898
rect 143728 129454 144048 129486
rect 143728 129218 143770 129454
rect 144006 129218 144048 129454
rect 143728 129134 144048 129218
rect 143728 128898 143770 129134
rect 144006 128898 144048 129134
rect 143728 128866 144048 128898
rect 174448 129454 174768 129486
rect 174448 129218 174490 129454
rect 174726 129218 174768 129454
rect 174448 129134 174768 129218
rect 174448 128898 174490 129134
rect 174726 128898 174768 129134
rect 174448 128866 174768 128898
rect 205168 129454 205488 129486
rect 205168 129218 205210 129454
rect 205446 129218 205488 129454
rect 205168 129134 205488 129218
rect 205168 128898 205210 129134
rect 205446 128898 205488 129134
rect 205168 128866 205488 128898
rect 235888 129454 236208 129486
rect 235888 129218 235930 129454
rect 236166 129218 236208 129454
rect 235888 129134 236208 129218
rect 235888 128898 235930 129134
rect 236166 128898 236208 129134
rect 235888 128866 236208 128898
rect 266608 129454 266928 129486
rect 266608 129218 266650 129454
rect 266886 129218 266928 129454
rect 266608 129134 266928 129218
rect 266608 128898 266650 129134
rect 266886 128898 266928 129134
rect 266608 128866 266928 128898
rect 297328 129454 297648 129486
rect 297328 129218 297370 129454
rect 297606 129218 297648 129454
rect 297328 129134 297648 129218
rect 297328 128898 297370 129134
rect 297606 128898 297648 129134
rect 297328 128866 297648 128898
rect 328048 129454 328368 129486
rect 328048 129218 328090 129454
rect 328326 129218 328368 129454
rect 328048 129134 328368 129218
rect 328048 128898 328090 129134
rect 328326 128898 328368 129134
rect 328048 128866 328368 128898
rect 358768 129454 359088 129486
rect 358768 129218 358810 129454
rect 359046 129218 359088 129454
rect 358768 129134 359088 129218
rect 358768 128898 358810 129134
rect 359046 128898 359088 129134
rect 358768 128866 359088 128898
rect 389488 129454 389808 129486
rect 389488 129218 389530 129454
rect 389766 129218 389808 129454
rect 389488 129134 389808 129218
rect 389488 128898 389530 129134
rect 389766 128898 389808 129134
rect 389488 128866 389808 128898
rect 420208 129454 420528 129486
rect 420208 129218 420250 129454
rect 420486 129218 420528 129454
rect 420208 129134 420528 129218
rect 420208 128898 420250 129134
rect 420486 128898 420528 129134
rect 420208 128866 420528 128898
rect 450928 129454 451248 129486
rect 450928 129218 450970 129454
rect 451206 129218 451248 129454
rect 450928 129134 451248 129218
rect 450928 128898 450970 129134
rect 451206 128898 451248 129134
rect 450928 128866 451248 128898
rect 481648 129454 481968 129486
rect 481648 129218 481690 129454
rect 481926 129218 481968 129454
rect 481648 129134 481968 129218
rect 481648 128898 481690 129134
rect 481926 128898 481968 129134
rect 481648 128866 481968 128898
rect 512368 129454 512688 129486
rect 512368 129218 512410 129454
rect 512646 129218 512688 129454
rect 512368 129134 512688 129218
rect 512368 128898 512410 129134
rect 512646 128898 512688 129134
rect 512368 128866 512688 128898
rect 543088 129454 543408 129486
rect 543088 129218 543130 129454
rect 543366 129218 543408 129454
rect 543088 129134 543408 129218
rect 543088 128898 543130 129134
rect 543366 128898 543408 129134
rect 543088 128866 543408 128898
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 36208 111454 36528 111486
rect 36208 111218 36250 111454
rect 36486 111218 36528 111454
rect 36208 111134 36528 111218
rect 36208 110898 36250 111134
rect 36486 110898 36528 111134
rect 36208 110866 36528 110898
rect 66928 111454 67248 111486
rect 66928 111218 66970 111454
rect 67206 111218 67248 111454
rect 66928 111134 67248 111218
rect 66928 110898 66970 111134
rect 67206 110898 67248 111134
rect 66928 110866 67248 110898
rect 97648 111454 97968 111486
rect 97648 111218 97690 111454
rect 97926 111218 97968 111454
rect 97648 111134 97968 111218
rect 97648 110898 97690 111134
rect 97926 110898 97968 111134
rect 97648 110866 97968 110898
rect 128368 111454 128688 111486
rect 128368 111218 128410 111454
rect 128646 111218 128688 111454
rect 128368 111134 128688 111218
rect 128368 110898 128410 111134
rect 128646 110898 128688 111134
rect 128368 110866 128688 110898
rect 159088 111454 159408 111486
rect 159088 111218 159130 111454
rect 159366 111218 159408 111454
rect 159088 111134 159408 111218
rect 159088 110898 159130 111134
rect 159366 110898 159408 111134
rect 159088 110866 159408 110898
rect 189808 111454 190128 111486
rect 189808 111218 189850 111454
rect 190086 111218 190128 111454
rect 189808 111134 190128 111218
rect 189808 110898 189850 111134
rect 190086 110898 190128 111134
rect 189808 110866 190128 110898
rect 220528 111454 220848 111486
rect 220528 111218 220570 111454
rect 220806 111218 220848 111454
rect 220528 111134 220848 111218
rect 220528 110898 220570 111134
rect 220806 110898 220848 111134
rect 220528 110866 220848 110898
rect 251248 111454 251568 111486
rect 251248 111218 251290 111454
rect 251526 111218 251568 111454
rect 251248 111134 251568 111218
rect 251248 110898 251290 111134
rect 251526 110898 251568 111134
rect 251248 110866 251568 110898
rect 281968 111454 282288 111486
rect 281968 111218 282010 111454
rect 282246 111218 282288 111454
rect 281968 111134 282288 111218
rect 281968 110898 282010 111134
rect 282246 110898 282288 111134
rect 281968 110866 282288 110898
rect 312688 111454 313008 111486
rect 312688 111218 312730 111454
rect 312966 111218 313008 111454
rect 312688 111134 313008 111218
rect 312688 110898 312730 111134
rect 312966 110898 313008 111134
rect 312688 110866 313008 110898
rect 343408 111454 343728 111486
rect 343408 111218 343450 111454
rect 343686 111218 343728 111454
rect 343408 111134 343728 111218
rect 343408 110898 343450 111134
rect 343686 110898 343728 111134
rect 343408 110866 343728 110898
rect 374128 111454 374448 111486
rect 374128 111218 374170 111454
rect 374406 111218 374448 111454
rect 374128 111134 374448 111218
rect 374128 110898 374170 111134
rect 374406 110898 374448 111134
rect 374128 110866 374448 110898
rect 404848 111454 405168 111486
rect 404848 111218 404890 111454
rect 405126 111218 405168 111454
rect 404848 111134 405168 111218
rect 404848 110898 404890 111134
rect 405126 110898 405168 111134
rect 404848 110866 405168 110898
rect 435568 111454 435888 111486
rect 435568 111218 435610 111454
rect 435846 111218 435888 111454
rect 435568 111134 435888 111218
rect 435568 110898 435610 111134
rect 435846 110898 435888 111134
rect 435568 110866 435888 110898
rect 466288 111454 466608 111486
rect 466288 111218 466330 111454
rect 466566 111218 466608 111454
rect 466288 111134 466608 111218
rect 466288 110898 466330 111134
rect 466566 110898 466608 111134
rect 466288 110866 466608 110898
rect 497008 111454 497328 111486
rect 497008 111218 497050 111454
rect 497286 111218 497328 111454
rect 497008 111134 497328 111218
rect 497008 110898 497050 111134
rect 497286 110898 497328 111134
rect 497008 110866 497328 110898
rect 527728 111454 528048 111486
rect 527728 111218 527770 111454
rect 528006 111218 528048 111454
rect 527728 111134 528048 111218
rect 527728 110898 527770 111134
rect 528006 110898 528048 111134
rect 527728 110866 528048 110898
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 51568 93454 51888 93486
rect 51568 93218 51610 93454
rect 51846 93218 51888 93454
rect 51568 93134 51888 93218
rect 51568 92898 51610 93134
rect 51846 92898 51888 93134
rect 51568 92866 51888 92898
rect 82288 93454 82608 93486
rect 82288 93218 82330 93454
rect 82566 93218 82608 93454
rect 82288 93134 82608 93218
rect 82288 92898 82330 93134
rect 82566 92898 82608 93134
rect 82288 92866 82608 92898
rect 113008 93454 113328 93486
rect 113008 93218 113050 93454
rect 113286 93218 113328 93454
rect 113008 93134 113328 93218
rect 113008 92898 113050 93134
rect 113286 92898 113328 93134
rect 113008 92866 113328 92898
rect 143728 93454 144048 93486
rect 143728 93218 143770 93454
rect 144006 93218 144048 93454
rect 143728 93134 144048 93218
rect 143728 92898 143770 93134
rect 144006 92898 144048 93134
rect 143728 92866 144048 92898
rect 174448 93454 174768 93486
rect 174448 93218 174490 93454
rect 174726 93218 174768 93454
rect 174448 93134 174768 93218
rect 174448 92898 174490 93134
rect 174726 92898 174768 93134
rect 174448 92866 174768 92898
rect 205168 93454 205488 93486
rect 205168 93218 205210 93454
rect 205446 93218 205488 93454
rect 205168 93134 205488 93218
rect 205168 92898 205210 93134
rect 205446 92898 205488 93134
rect 205168 92866 205488 92898
rect 235888 93454 236208 93486
rect 235888 93218 235930 93454
rect 236166 93218 236208 93454
rect 235888 93134 236208 93218
rect 235888 92898 235930 93134
rect 236166 92898 236208 93134
rect 235888 92866 236208 92898
rect 266608 93454 266928 93486
rect 266608 93218 266650 93454
rect 266886 93218 266928 93454
rect 266608 93134 266928 93218
rect 266608 92898 266650 93134
rect 266886 92898 266928 93134
rect 266608 92866 266928 92898
rect 297328 93454 297648 93486
rect 297328 93218 297370 93454
rect 297606 93218 297648 93454
rect 297328 93134 297648 93218
rect 297328 92898 297370 93134
rect 297606 92898 297648 93134
rect 297328 92866 297648 92898
rect 328048 93454 328368 93486
rect 328048 93218 328090 93454
rect 328326 93218 328368 93454
rect 328048 93134 328368 93218
rect 328048 92898 328090 93134
rect 328326 92898 328368 93134
rect 328048 92866 328368 92898
rect 358768 93454 359088 93486
rect 358768 93218 358810 93454
rect 359046 93218 359088 93454
rect 358768 93134 359088 93218
rect 358768 92898 358810 93134
rect 359046 92898 359088 93134
rect 358768 92866 359088 92898
rect 389488 93454 389808 93486
rect 389488 93218 389530 93454
rect 389766 93218 389808 93454
rect 389488 93134 389808 93218
rect 389488 92898 389530 93134
rect 389766 92898 389808 93134
rect 389488 92866 389808 92898
rect 420208 93454 420528 93486
rect 420208 93218 420250 93454
rect 420486 93218 420528 93454
rect 420208 93134 420528 93218
rect 420208 92898 420250 93134
rect 420486 92898 420528 93134
rect 420208 92866 420528 92898
rect 450928 93454 451248 93486
rect 450928 93218 450970 93454
rect 451206 93218 451248 93454
rect 450928 93134 451248 93218
rect 450928 92898 450970 93134
rect 451206 92898 451248 93134
rect 450928 92866 451248 92898
rect 481648 93454 481968 93486
rect 481648 93218 481690 93454
rect 481926 93218 481968 93454
rect 481648 93134 481968 93218
rect 481648 92898 481690 93134
rect 481926 92898 481968 93134
rect 481648 92866 481968 92898
rect 512368 93454 512688 93486
rect 512368 93218 512410 93454
rect 512646 93218 512688 93454
rect 512368 93134 512688 93218
rect 512368 92898 512410 93134
rect 512646 92898 512688 93134
rect 512368 92866 512688 92898
rect 543088 93454 543408 93486
rect 543088 93218 543130 93454
rect 543366 93218 543408 93454
rect 543088 93134 543408 93218
rect 543088 92898 543130 93134
rect 543366 92898 543408 93134
rect 543088 92866 543408 92898
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 36208 75454 36528 75486
rect 36208 75218 36250 75454
rect 36486 75218 36528 75454
rect 36208 75134 36528 75218
rect 36208 74898 36250 75134
rect 36486 74898 36528 75134
rect 36208 74866 36528 74898
rect 66928 75454 67248 75486
rect 66928 75218 66970 75454
rect 67206 75218 67248 75454
rect 66928 75134 67248 75218
rect 66928 74898 66970 75134
rect 67206 74898 67248 75134
rect 66928 74866 67248 74898
rect 97648 75454 97968 75486
rect 97648 75218 97690 75454
rect 97926 75218 97968 75454
rect 97648 75134 97968 75218
rect 97648 74898 97690 75134
rect 97926 74898 97968 75134
rect 97648 74866 97968 74898
rect 128368 75454 128688 75486
rect 128368 75218 128410 75454
rect 128646 75218 128688 75454
rect 128368 75134 128688 75218
rect 128368 74898 128410 75134
rect 128646 74898 128688 75134
rect 128368 74866 128688 74898
rect 159088 75454 159408 75486
rect 159088 75218 159130 75454
rect 159366 75218 159408 75454
rect 159088 75134 159408 75218
rect 159088 74898 159130 75134
rect 159366 74898 159408 75134
rect 159088 74866 159408 74898
rect 189808 75454 190128 75486
rect 189808 75218 189850 75454
rect 190086 75218 190128 75454
rect 189808 75134 190128 75218
rect 189808 74898 189850 75134
rect 190086 74898 190128 75134
rect 189808 74866 190128 74898
rect 220528 75454 220848 75486
rect 220528 75218 220570 75454
rect 220806 75218 220848 75454
rect 220528 75134 220848 75218
rect 220528 74898 220570 75134
rect 220806 74898 220848 75134
rect 220528 74866 220848 74898
rect 251248 75454 251568 75486
rect 251248 75218 251290 75454
rect 251526 75218 251568 75454
rect 251248 75134 251568 75218
rect 251248 74898 251290 75134
rect 251526 74898 251568 75134
rect 251248 74866 251568 74898
rect 281968 75454 282288 75486
rect 281968 75218 282010 75454
rect 282246 75218 282288 75454
rect 281968 75134 282288 75218
rect 281968 74898 282010 75134
rect 282246 74898 282288 75134
rect 281968 74866 282288 74898
rect 312688 75454 313008 75486
rect 312688 75218 312730 75454
rect 312966 75218 313008 75454
rect 312688 75134 313008 75218
rect 312688 74898 312730 75134
rect 312966 74898 313008 75134
rect 312688 74866 313008 74898
rect 343408 75454 343728 75486
rect 343408 75218 343450 75454
rect 343686 75218 343728 75454
rect 343408 75134 343728 75218
rect 343408 74898 343450 75134
rect 343686 74898 343728 75134
rect 343408 74866 343728 74898
rect 374128 75454 374448 75486
rect 374128 75218 374170 75454
rect 374406 75218 374448 75454
rect 374128 75134 374448 75218
rect 374128 74898 374170 75134
rect 374406 74898 374448 75134
rect 374128 74866 374448 74898
rect 404848 75454 405168 75486
rect 404848 75218 404890 75454
rect 405126 75218 405168 75454
rect 404848 75134 405168 75218
rect 404848 74898 404890 75134
rect 405126 74898 405168 75134
rect 404848 74866 405168 74898
rect 435568 75454 435888 75486
rect 435568 75218 435610 75454
rect 435846 75218 435888 75454
rect 435568 75134 435888 75218
rect 435568 74898 435610 75134
rect 435846 74898 435888 75134
rect 435568 74866 435888 74898
rect 466288 75454 466608 75486
rect 466288 75218 466330 75454
rect 466566 75218 466608 75454
rect 466288 75134 466608 75218
rect 466288 74898 466330 75134
rect 466566 74898 466608 75134
rect 466288 74866 466608 74898
rect 497008 75454 497328 75486
rect 497008 75218 497050 75454
rect 497286 75218 497328 75454
rect 497008 75134 497328 75218
rect 497008 74898 497050 75134
rect 497286 74898 497328 75134
rect 497008 74866 497328 74898
rect 527728 75454 528048 75486
rect 527728 75218 527770 75454
rect 528006 75218 528048 75454
rect 527728 75134 528048 75218
rect 527728 74898 527770 75134
rect 528006 74898 528048 75134
rect 527728 74866 528048 74898
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 51568 57454 51888 57486
rect 51568 57218 51610 57454
rect 51846 57218 51888 57454
rect 51568 57134 51888 57218
rect 51568 56898 51610 57134
rect 51846 56898 51888 57134
rect 51568 56866 51888 56898
rect 82288 57454 82608 57486
rect 82288 57218 82330 57454
rect 82566 57218 82608 57454
rect 82288 57134 82608 57218
rect 82288 56898 82330 57134
rect 82566 56898 82608 57134
rect 82288 56866 82608 56898
rect 113008 57454 113328 57486
rect 113008 57218 113050 57454
rect 113286 57218 113328 57454
rect 113008 57134 113328 57218
rect 113008 56898 113050 57134
rect 113286 56898 113328 57134
rect 113008 56866 113328 56898
rect 143728 57454 144048 57486
rect 143728 57218 143770 57454
rect 144006 57218 144048 57454
rect 143728 57134 144048 57218
rect 143728 56898 143770 57134
rect 144006 56898 144048 57134
rect 143728 56866 144048 56898
rect 174448 57454 174768 57486
rect 174448 57218 174490 57454
rect 174726 57218 174768 57454
rect 174448 57134 174768 57218
rect 174448 56898 174490 57134
rect 174726 56898 174768 57134
rect 174448 56866 174768 56898
rect 205168 57454 205488 57486
rect 205168 57218 205210 57454
rect 205446 57218 205488 57454
rect 205168 57134 205488 57218
rect 205168 56898 205210 57134
rect 205446 56898 205488 57134
rect 205168 56866 205488 56898
rect 235888 57454 236208 57486
rect 235888 57218 235930 57454
rect 236166 57218 236208 57454
rect 235888 57134 236208 57218
rect 235888 56898 235930 57134
rect 236166 56898 236208 57134
rect 235888 56866 236208 56898
rect 266608 57454 266928 57486
rect 266608 57218 266650 57454
rect 266886 57218 266928 57454
rect 266608 57134 266928 57218
rect 266608 56898 266650 57134
rect 266886 56898 266928 57134
rect 266608 56866 266928 56898
rect 297328 57454 297648 57486
rect 297328 57218 297370 57454
rect 297606 57218 297648 57454
rect 297328 57134 297648 57218
rect 297328 56898 297370 57134
rect 297606 56898 297648 57134
rect 297328 56866 297648 56898
rect 328048 57454 328368 57486
rect 328048 57218 328090 57454
rect 328326 57218 328368 57454
rect 328048 57134 328368 57218
rect 328048 56898 328090 57134
rect 328326 56898 328368 57134
rect 328048 56866 328368 56898
rect 358768 57454 359088 57486
rect 358768 57218 358810 57454
rect 359046 57218 359088 57454
rect 358768 57134 359088 57218
rect 358768 56898 358810 57134
rect 359046 56898 359088 57134
rect 358768 56866 359088 56898
rect 389488 57454 389808 57486
rect 389488 57218 389530 57454
rect 389766 57218 389808 57454
rect 389488 57134 389808 57218
rect 389488 56898 389530 57134
rect 389766 56898 389808 57134
rect 389488 56866 389808 56898
rect 420208 57454 420528 57486
rect 420208 57218 420250 57454
rect 420486 57218 420528 57454
rect 420208 57134 420528 57218
rect 420208 56898 420250 57134
rect 420486 56898 420528 57134
rect 420208 56866 420528 56898
rect 450928 57454 451248 57486
rect 450928 57218 450970 57454
rect 451206 57218 451248 57454
rect 450928 57134 451248 57218
rect 450928 56898 450970 57134
rect 451206 56898 451248 57134
rect 450928 56866 451248 56898
rect 481648 57454 481968 57486
rect 481648 57218 481690 57454
rect 481926 57218 481968 57454
rect 481648 57134 481968 57218
rect 481648 56898 481690 57134
rect 481926 56898 481968 57134
rect 481648 56866 481968 56898
rect 512368 57454 512688 57486
rect 512368 57218 512410 57454
rect 512646 57218 512688 57454
rect 512368 57134 512688 57218
rect 512368 56898 512410 57134
rect 512646 56898 512688 57134
rect 512368 56866 512688 56898
rect 543088 57454 543408 57486
rect 543088 57218 543130 57454
rect 543366 57218 543408 57454
rect 543088 57134 543408 57218
rect 543088 56898 543130 57134
rect 543366 56898 543408 57134
rect 543088 56866 543408 56898
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 36208 39454 36528 39486
rect 36208 39218 36250 39454
rect 36486 39218 36528 39454
rect 36208 39134 36528 39218
rect 36208 38898 36250 39134
rect 36486 38898 36528 39134
rect 36208 38866 36528 38898
rect 66928 39454 67248 39486
rect 66928 39218 66970 39454
rect 67206 39218 67248 39454
rect 66928 39134 67248 39218
rect 66928 38898 66970 39134
rect 67206 38898 67248 39134
rect 66928 38866 67248 38898
rect 97648 39454 97968 39486
rect 97648 39218 97690 39454
rect 97926 39218 97968 39454
rect 97648 39134 97968 39218
rect 97648 38898 97690 39134
rect 97926 38898 97968 39134
rect 97648 38866 97968 38898
rect 128368 39454 128688 39486
rect 128368 39218 128410 39454
rect 128646 39218 128688 39454
rect 128368 39134 128688 39218
rect 128368 38898 128410 39134
rect 128646 38898 128688 39134
rect 128368 38866 128688 38898
rect 159088 39454 159408 39486
rect 159088 39218 159130 39454
rect 159366 39218 159408 39454
rect 159088 39134 159408 39218
rect 159088 38898 159130 39134
rect 159366 38898 159408 39134
rect 159088 38866 159408 38898
rect 189808 39454 190128 39486
rect 189808 39218 189850 39454
rect 190086 39218 190128 39454
rect 189808 39134 190128 39218
rect 189808 38898 189850 39134
rect 190086 38898 190128 39134
rect 189808 38866 190128 38898
rect 220528 39454 220848 39486
rect 220528 39218 220570 39454
rect 220806 39218 220848 39454
rect 220528 39134 220848 39218
rect 220528 38898 220570 39134
rect 220806 38898 220848 39134
rect 220528 38866 220848 38898
rect 251248 39454 251568 39486
rect 251248 39218 251290 39454
rect 251526 39218 251568 39454
rect 251248 39134 251568 39218
rect 251248 38898 251290 39134
rect 251526 38898 251568 39134
rect 251248 38866 251568 38898
rect 281968 39454 282288 39486
rect 281968 39218 282010 39454
rect 282246 39218 282288 39454
rect 281968 39134 282288 39218
rect 281968 38898 282010 39134
rect 282246 38898 282288 39134
rect 281968 38866 282288 38898
rect 312688 39454 313008 39486
rect 312688 39218 312730 39454
rect 312966 39218 313008 39454
rect 312688 39134 313008 39218
rect 312688 38898 312730 39134
rect 312966 38898 313008 39134
rect 312688 38866 313008 38898
rect 343408 39454 343728 39486
rect 343408 39218 343450 39454
rect 343686 39218 343728 39454
rect 343408 39134 343728 39218
rect 343408 38898 343450 39134
rect 343686 38898 343728 39134
rect 343408 38866 343728 38898
rect 374128 39454 374448 39486
rect 374128 39218 374170 39454
rect 374406 39218 374448 39454
rect 374128 39134 374448 39218
rect 374128 38898 374170 39134
rect 374406 38898 374448 39134
rect 374128 38866 374448 38898
rect 404848 39454 405168 39486
rect 404848 39218 404890 39454
rect 405126 39218 405168 39454
rect 404848 39134 405168 39218
rect 404848 38898 404890 39134
rect 405126 38898 405168 39134
rect 404848 38866 405168 38898
rect 435568 39454 435888 39486
rect 435568 39218 435610 39454
rect 435846 39218 435888 39454
rect 435568 39134 435888 39218
rect 435568 38898 435610 39134
rect 435846 38898 435888 39134
rect 435568 38866 435888 38898
rect 466288 39454 466608 39486
rect 466288 39218 466330 39454
rect 466566 39218 466608 39454
rect 466288 39134 466608 39218
rect 466288 38898 466330 39134
rect 466566 38898 466608 39134
rect 466288 38866 466608 38898
rect 497008 39454 497328 39486
rect 497008 39218 497050 39454
rect 497286 39218 497328 39454
rect 497008 39134 497328 39218
rect 497008 38898 497050 39134
rect 497286 38898 497328 39134
rect 497008 38866 497328 38898
rect 527728 39454 528048 39486
rect 527728 39218 527770 39454
rect 528006 39218 528048 39454
rect 527728 39134 528048 39218
rect 527728 38898 527770 39134
rect 528006 38898 528048 39134
rect 527728 38866 528048 38898
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 30000
rect 37794 3454 38414 30000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 7174 42134 30000
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 10894 45854 30000
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 30000
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 30000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 30000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 30000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 30000
rect 73794 3454 74414 30000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 30000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 30000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 30000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 30000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 30000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 30000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 30000
rect 109794 3454 110414 30000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 30000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 30000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 30000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 30000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 30000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 30000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 30000
rect 145794 3454 146414 30000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 7174 150134 30000
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 30000
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 30000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 30000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 30000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 30000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 30000
rect 181794 3454 182414 30000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 30000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 30000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 30000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 30000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 30000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 30000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 30000
rect 217794 3454 218414 30000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 30000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 30000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 30000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 30000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 30000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 30000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 30000
rect 253794 3454 254414 30000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 30000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 30000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 30000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 30000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 30000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 30000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 30000
rect 289794 3454 290414 30000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 30000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 30000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 30000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 30000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 30000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 30000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 30000
rect 325794 3454 326414 30000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 30000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 30000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 30000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 30000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 30000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 30000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 30000
rect 361794 3454 362414 30000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 30000
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 30000
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 30000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 30000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 30000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 30000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 30000
rect 397794 3454 398414 30000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 30000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 30000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 30000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 30000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 30000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 30000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 30000
rect 433794 3454 434414 30000
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 30000
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 30000
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 30000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 30000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 30000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 30000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 30000
rect 469794 3454 470414 30000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 7174 474134 30000
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 10894 477854 30000
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 30000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 30000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 30000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 30000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 30000
rect 505794 3454 506414 30000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 7174 510134 30000
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 10894 513854 30000
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 30000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 30000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 30000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 28894 531854 30000
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 30000
rect 541794 3454 542414 30000
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 7174 546134 30000
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 10894 549854 30000
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 14614 553574 30000
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 51610 669218 51846 669454
rect 51610 668898 51846 669134
rect 82330 669218 82566 669454
rect 82330 668898 82566 669134
rect 113050 669218 113286 669454
rect 113050 668898 113286 669134
rect 143770 669218 144006 669454
rect 143770 668898 144006 669134
rect 174490 669218 174726 669454
rect 174490 668898 174726 669134
rect 205210 669218 205446 669454
rect 205210 668898 205446 669134
rect 235930 669218 236166 669454
rect 235930 668898 236166 669134
rect 266650 669218 266886 669454
rect 266650 668898 266886 669134
rect 297370 669218 297606 669454
rect 297370 668898 297606 669134
rect 328090 669218 328326 669454
rect 328090 668898 328326 669134
rect 358810 669218 359046 669454
rect 358810 668898 359046 669134
rect 389530 669218 389766 669454
rect 389530 668898 389766 669134
rect 420250 669218 420486 669454
rect 420250 668898 420486 669134
rect 450970 669218 451206 669454
rect 450970 668898 451206 669134
rect 481690 669218 481926 669454
rect 481690 668898 481926 669134
rect 512410 669218 512646 669454
rect 512410 668898 512646 669134
rect 543130 669218 543366 669454
rect 543130 668898 543366 669134
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 36250 651218 36486 651454
rect 36250 650898 36486 651134
rect 66970 651218 67206 651454
rect 66970 650898 67206 651134
rect 97690 651218 97926 651454
rect 97690 650898 97926 651134
rect 128410 651218 128646 651454
rect 128410 650898 128646 651134
rect 159130 651218 159366 651454
rect 159130 650898 159366 651134
rect 189850 651218 190086 651454
rect 189850 650898 190086 651134
rect 220570 651218 220806 651454
rect 220570 650898 220806 651134
rect 251290 651218 251526 651454
rect 251290 650898 251526 651134
rect 282010 651218 282246 651454
rect 282010 650898 282246 651134
rect 312730 651218 312966 651454
rect 312730 650898 312966 651134
rect 343450 651218 343686 651454
rect 343450 650898 343686 651134
rect 374170 651218 374406 651454
rect 374170 650898 374406 651134
rect 404890 651218 405126 651454
rect 404890 650898 405126 651134
rect 435610 651218 435846 651454
rect 435610 650898 435846 651134
rect 466330 651218 466566 651454
rect 466330 650898 466566 651134
rect 497050 651218 497286 651454
rect 497050 650898 497286 651134
rect 527770 651218 528006 651454
rect 527770 650898 528006 651134
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 51610 633218 51846 633454
rect 51610 632898 51846 633134
rect 82330 633218 82566 633454
rect 82330 632898 82566 633134
rect 113050 633218 113286 633454
rect 113050 632898 113286 633134
rect 143770 633218 144006 633454
rect 143770 632898 144006 633134
rect 174490 633218 174726 633454
rect 174490 632898 174726 633134
rect 205210 633218 205446 633454
rect 205210 632898 205446 633134
rect 235930 633218 236166 633454
rect 235930 632898 236166 633134
rect 266650 633218 266886 633454
rect 266650 632898 266886 633134
rect 297370 633218 297606 633454
rect 297370 632898 297606 633134
rect 328090 633218 328326 633454
rect 328090 632898 328326 633134
rect 358810 633218 359046 633454
rect 358810 632898 359046 633134
rect 389530 633218 389766 633454
rect 389530 632898 389766 633134
rect 420250 633218 420486 633454
rect 420250 632898 420486 633134
rect 450970 633218 451206 633454
rect 450970 632898 451206 633134
rect 481690 633218 481926 633454
rect 481690 632898 481926 633134
rect 512410 633218 512646 633454
rect 512410 632898 512646 633134
rect 543130 633218 543366 633454
rect 543130 632898 543366 633134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 36250 615218 36486 615454
rect 36250 614898 36486 615134
rect 66970 615218 67206 615454
rect 66970 614898 67206 615134
rect 97690 615218 97926 615454
rect 97690 614898 97926 615134
rect 128410 615218 128646 615454
rect 128410 614898 128646 615134
rect 159130 615218 159366 615454
rect 159130 614898 159366 615134
rect 189850 615218 190086 615454
rect 189850 614898 190086 615134
rect 220570 615218 220806 615454
rect 220570 614898 220806 615134
rect 251290 615218 251526 615454
rect 251290 614898 251526 615134
rect 282010 615218 282246 615454
rect 282010 614898 282246 615134
rect 312730 615218 312966 615454
rect 312730 614898 312966 615134
rect 343450 615218 343686 615454
rect 343450 614898 343686 615134
rect 374170 615218 374406 615454
rect 374170 614898 374406 615134
rect 404890 615218 405126 615454
rect 404890 614898 405126 615134
rect 435610 615218 435846 615454
rect 435610 614898 435846 615134
rect 466330 615218 466566 615454
rect 466330 614898 466566 615134
rect 497050 615218 497286 615454
rect 497050 614898 497286 615134
rect 527770 615218 528006 615454
rect 527770 614898 528006 615134
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 51610 597218 51846 597454
rect 51610 596898 51846 597134
rect 82330 597218 82566 597454
rect 82330 596898 82566 597134
rect 113050 597218 113286 597454
rect 113050 596898 113286 597134
rect 143770 597218 144006 597454
rect 143770 596898 144006 597134
rect 174490 597218 174726 597454
rect 174490 596898 174726 597134
rect 205210 597218 205446 597454
rect 205210 596898 205446 597134
rect 235930 597218 236166 597454
rect 235930 596898 236166 597134
rect 266650 597218 266886 597454
rect 266650 596898 266886 597134
rect 297370 597218 297606 597454
rect 297370 596898 297606 597134
rect 328090 597218 328326 597454
rect 328090 596898 328326 597134
rect 358810 597218 359046 597454
rect 358810 596898 359046 597134
rect 389530 597218 389766 597454
rect 389530 596898 389766 597134
rect 420250 597218 420486 597454
rect 420250 596898 420486 597134
rect 450970 597218 451206 597454
rect 450970 596898 451206 597134
rect 481690 597218 481926 597454
rect 481690 596898 481926 597134
rect 512410 597218 512646 597454
rect 512410 596898 512646 597134
rect 543130 597218 543366 597454
rect 543130 596898 543366 597134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 36250 579218 36486 579454
rect 36250 578898 36486 579134
rect 66970 579218 67206 579454
rect 66970 578898 67206 579134
rect 97690 579218 97926 579454
rect 97690 578898 97926 579134
rect 128410 579218 128646 579454
rect 128410 578898 128646 579134
rect 159130 579218 159366 579454
rect 159130 578898 159366 579134
rect 189850 579218 190086 579454
rect 189850 578898 190086 579134
rect 220570 579218 220806 579454
rect 220570 578898 220806 579134
rect 251290 579218 251526 579454
rect 251290 578898 251526 579134
rect 282010 579218 282246 579454
rect 282010 578898 282246 579134
rect 312730 579218 312966 579454
rect 312730 578898 312966 579134
rect 343450 579218 343686 579454
rect 343450 578898 343686 579134
rect 374170 579218 374406 579454
rect 374170 578898 374406 579134
rect 404890 579218 405126 579454
rect 404890 578898 405126 579134
rect 435610 579218 435846 579454
rect 435610 578898 435846 579134
rect 466330 579218 466566 579454
rect 466330 578898 466566 579134
rect 497050 579218 497286 579454
rect 497050 578898 497286 579134
rect 527770 579218 528006 579454
rect 527770 578898 528006 579134
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 51610 561218 51846 561454
rect 51610 560898 51846 561134
rect 82330 561218 82566 561454
rect 82330 560898 82566 561134
rect 113050 561218 113286 561454
rect 113050 560898 113286 561134
rect 143770 561218 144006 561454
rect 143770 560898 144006 561134
rect 174490 561218 174726 561454
rect 174490 560898 174726 561134
rect 205210 561218 205446 561454
rect 205210 560898 205446 561134
rect 235930 561218 236166 561454
rect 235930 560898 236166 561134
rect 266650 561218 266886 561454
rect 266650 560898 266886 561134
rect 297370 561218 297606 561454
rect 297370 560898 297606 561134
rect 328090 561218 328326 561454
rect 328090 560898 328326 561134
rect 358810 561218 359046 561454
rect 358810 560898 359046 561134
rect 389530 561218 389766 561454
rect 389530 560898 389766 561134
rect 420250 561218 420486 561454
rect 420250 560898 420486 561134
rect 450970 561218 451206 561454
rect 450970 560898 451206 561134
rect 481690 561218 481926 561454
rect 481690 560898 481926 561134
rect 512410 561218 512646 561454
rect 512410 560898 512646 561134
rect 543130 561218 543366 561454
rect 543130 560898 543366 561134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 36250 543218 36486 543454
rect 36250 542898 36486 543134
rect 66970 543218 67206 543454
rect 66970 542898 67206 543134
rect 97690 543218 97926 543454
rect 97690 542898 97926 543134
rect 128410 543218 128646 543454
rect 128410 542898 128646 543134
rect 159130 543218 159366 543454
rect 159130 542898 159366 543134
rect 189850 543218 190086 543454
rect 189850 542898 190086 543134
rect 220570 543218 220806 543454
rect 220570 542898 220806 543134
rect 251290 543218 251526 543454
rect 251290 542898 251526 543134
rect 282010 543218 282246 543454
rect 282010 542898 282246 543134
rect 312730 543218 312966 543454
rect 312730 542898 312966 543134
rect 343450 543218 343686 543454
rect 343450 542898 343686 543134
rect 374170 543218 374406 543454
rect 374170 542898 374406 543134
rect 404890 543218 405126 543454
rect 404890 542898 405126 543134
rect 435610 543218 435846 543454
rect 435610 542898 435846 543134
rect 466330 543218 466566 543454
rect 466330 542898 466566 543134
rect 497050 543218 497286 543454
rect 497050 542898 497286 543134
rect 527770 543218 528006 543454
rect 527770 542898 528006 543134
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 51610 525218 51846 525454
rect 51610 524898 51846 525134
rect 82330 525218 82566 525454
rect 82330 524898 82566 525134
rect 113050 525218 113286 525454
rect 113050 524898 113286 525134
rect 143770 525218 144006 525454
rect 143770 524898 144006 525134
rect 174490 525218 174726 525454
rect 174490 524898 174726 525134
rect 205210 525218 205446 525454
rect 205210 524898 205446 525134
rect 235930 525218 236166 525454
rect 235930 524898 236166 525134
rect 266650 525218 266886 525454
rect 266650 524898 266886 525134
rect 297370 525218 297606 525454
rect 297370 524898 297606 525134
rect 328090 525218 328326 525454
rect 328090 524898 328326 525134
rect 358810 525218 359046 525454
rect 358810 524898 359046 525134
rect 389530 525218 389766 525454
rect 389530 524898 389766 525134
rect 420250 525218 420486 525454
rect 420250 524898 420486 525134
rect 450970 525218 451206 525454
rect 450970 524898 451206 525134
rect 481690 525218 481926 525454
rect 481690 524898 481926 525134
rect 512410 525218 512646 525454
rect 512410 524898 512646 525134
rect 543130 525218 543366 525454
rect 543130 524898 543366 525134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 36250 507218 36486 507454
rect 36250 506898 36486 507134
rect 66970 507218 67206 507454
rect 66970 506898 67206 507134
rect 97690 507218 97926 507454
rect 97690 506898 97926 507134
rect 128410 507218 128646 507454
rect 128410 506898 128646 507134
rect 159130 507218 159366 507454
rect 159130 506898 159366 507134
rect 189850 507218 190086 507454
rect 189850 506898 190086 507134
rect 220570 507218 220806 507454
rect 220570 506898 220806 507134
rect 251290 507218 251526 507454
rect 251290 506898 251526 507134
rect 282010 507218 282246 507454
rect 282010 506898 282246 507134
rect 312730 507218 312966 507454
rect 312730 506898 312966 507134
rect 343450 507218 343686 507454
rect 343450 506898 343686 507134
rect 374170 507218 374406 507454
rect 374170 506898 374406 507134
rect 404890 507218 405126 507454
rect 404890 506898 405126 507134
rect 435610 507218 435846 507454
rect 435610 506898 435846 507134
rect 466330 507218 466566 507454
rect 466330 506898 466566 507134
rect 497050 507218 497286 507454
rect 497050 506898 497286 507134
rect 527770 507218 528006 507454
rect 527770 506898 528006 507134
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 51610 489218 51846 489454
rect 51610 488898 51846 489134
rect 82330 489218 82566 489454
rect 82330 488898 82566 489134
rect 113050 489218 113286 489454
rect 113050 488898 113286 489134
rect 143770 489218 144006 489454
rect 143770 488898 144006 489134
rect 174490 489218 174726 489454
rect 174490 488898 174726 489134
rect 205210 489218 205446 489454
rect 205210 488898 205446 489134
rect 235930 489218 236166 489454
rect 235930 488898 236166 489134
rect 266650 489218 266886 489454
rect 266650 488898 266886 489134
rect 297370 489218 297606 489454
rect 297370 488898 297606 489134
rect 328090 489218 328326 489454
rect 328090 488898 328326 489134
rect 358810 489218 359046 489454
rect 358810 488898 359046 489134
rect 389530 489218 389766 489454
rect 389530 488898 389766 489134
rect 420250 489218 420486 489454
rect 420250 488898 420486 489134
rect 450970 489218 451206 489454
rect 450970 488898 451206 489134
rect 481690 489218 481926 489454
rect 481690 488898 481926 489134
rect 512410 489218 512646 489454
rect 512410 488898 512646 489134
rect 543130 489218 543366 489454
rect 543130 488898 543366 489134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 36250 471218 36486 471454
rect 36250 470898 36486 471134
rect 66970 471218 67206 471454
rect 66970 470898 67206 471134
rect 97690 471218 97926 471454
rect 97690 470898 97926 471134
rect 128410 471218 128646 471454
rect 128410 470898 128646 471134
rect 159130 471218 159366 471454
rect 159130 470898 159366 471134
rect 189850 471218 190086 471454
rect 189850 470898 190086 471134
rect 220570 471218 220806 471454
rect 220570 470898 220806 471134
rect 251290 471218 251526 471454
rect 251290 470898 251526 471134
rect 282010 471218 282246 471454
rect 282010 470898 282246 471134
rect 312730 471218 312966 471454
rect 312730 470898 312966 471134
rect 343450 471218 343686 471454
rect 343450 470898 343686 471134
rect 374170 471218 374406 471454
rect 374170 470898 374406 471134
rect 404890 471218 405126 471454
rect 404890 470898 405126 471134
rect 435610 471218 435846 471454
rect 435610 470898 435846 471134
rect 466330 471218 466566 471454
rect 466330 470898 466566 471134
rect 497050 471218 497286 471454
rect 497050 470898 497286 471134
rect 527770 471218 528006 471454
rect 527770 470898 528006 471134
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 51610 453218 51846 453454
rect 51610 452898 51846 453134
rect 82330 453218 82566 453454
rect 82330 452898 82566 453134
rect 113050 453218 113286 453454
rect 113050 452898 113286 453134
rect 143770 453218 144006 453454
rect 143770 452898 144006 453134
rect 174490 453218 174726 453454
rect 174490 452898 174726 453134
rect 205210 453218 205446 453454
rect 205210 452898 205446 453134
rect 235930 453218 236166 453454
rect 235930 452898 236166 453134
rect 266650 453218 266886 453454
rect 266650 452898 266886 453134
rect 297370 453218 297606 453454
rect 297370 452898 297606 453134
rect 328090 453218 328326 453454
rect 328090 452898 328326 453134
rect 358810 453218 359046 453454
rect 358810 452898 359046 453134
rect 389530 453218 389766 453454
rect 389530 452898 389766 453134
rect 420250 453218 420486 453454
rect 420250 452898 420486 453134
rect 450970 453218 451206 453454
rect 450970 452898 451206 453134
rect 481690 453218 481926 453454
rect 481690 452898 481926 453134
rect 512410 453218 512646 453454
rect 512410 452898 512646 453134
rect 543130 453218 543366 453454
rect 543130 452898 543366 453134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 36250 435218 36486 435454
rect 36250 434898 36486 435134
rect 66970 435218 67206 435454
rect 66970 434898 67206 435134
rect 97690 435218 97926 435454
rect 97690 434898 97926 435134
rect 128410 435218 128646 435454
rect 128410 434898 128646 435134
rect 159130 435218 159366 435454
rect 159130 434898 159366 435134
rect 189850 435218 190086 435454
rect 189850 434898 190086 435134
rect 220570 435218 220806 435454
rect 220570 434898 220806 435134
rect 251290 435218 251526 435454
rect 251290 434898 251526 435134
rect 282010 435218 282246 435454
rect 282010 434898 282246 435134
rect 312730 435218 312966 435454
rect 312730 434898 312966 435134
rect 343450 435218 343686 435454
rect 343450 434898 343686 435134
rect 374170 435218 374406 435454
rect 374170 434898 374406 435134
rect 404890 435218 405126 435454
rect 404890 434898 405126 435134
rect 435610 435218 435846 435454
rect 435610 434898 435846 435134
rect 466330 435218 466566 435454
rect 466330 434898 466566 435134
rect 497050 435218 497286 435454
rect 497050 434898 497286 435134
rect 527770 435218 528006 435454
rect 527770 434898 528006 435134
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 51610 417218 51846 417454
rect 51610 416898 51846 417134
rect 82330 417218 82566 417454
rect 82330 416898 82566 417134
rect 113050 417218 113286 417454
rect 113050 416898 113286 417134
rect 143770 417218 144006 417454
rect 143770 416898 144006 417134
rect 174490 417218 174726 417454
rect 174490 416898 174726 417134
rect 205210 417218 205446 417454
rect 205210 416898 205446 417134
rect 235930 417218 236166 417454
rect 235930 416898 236166 417134
rect 266650 417218 266886 417454
rect 266650 416898 266886 417134
rect 297370 417218 297606 417454
rect 297370 416898 297606 417134
rect 328090 417218 328326 417454
rect 328090 416898 328326 417134
rect 358810 417218 359046 417454
rect 358810 416898 359046 417134
rect 389530 417218 389766 417454
rect 389530 416898 389766 417134
rect 420250 417218 420486 417454
rect 420250 416898 420486 417134
rect 450970 417218 451206 417454
rect 450970 416898 451206 417134
rect 481690 417218 481926 417454
rect 481690 416898 481926 417134
rect 512410 417218 512646 417454
rect 512410 416898 512646 417134
rect 543130 417218 543366 417454
rect 543130 416898 543366 417134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 36250 399218 36486 399454
rect 36250 398898 36486 399134
rect 66970 399218 67206 399454
rect 66970 398898 67206 399134
rect 97690 399218 97926 399454
rect 97690 398898 97926 399134
rect 128410 399218 128646 399454
rect 128410 398898 128646 399134
rect 159130 399218 159366 399454
rect 159130 398898 159366 399134
rect 189850 399218 190086 399454
rect 189850 398898 190086 399134
rect 220570 399218 220806 399454
rect 220570 398898 220806 399134
rect 251290 399218 251526 399454
rect 251290 398898 251526 399134
rect 282010 399218 282246 399454
rect 282010 398898 282246 399134
rect 312730 399218 312966 399454
rect 312730 398898 312966 399134
rect 343450 399218 343686 399454
rect 343450 398898 343686 399134
rect 374170 399218 374406 399454
rect 374170 398898 374406 399134
rect 404890 399218 405126 399454
rect 404890 398898 405126 399134
rect 435610 399218 435846 399454
rect 435610 398898 435846 399134
rect 466330 399218 466566 399454
rect 466330 398898 466566 399134
rect 497050 399218 497286 399454
rect 497050 398898 497286 399134
rect 527770 399218 528006 399454
rect 527770 398898 528006 399134
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 51610 381218 51846 381454
rect 51610 380898 51846 381134
rect 82330 381218 82566 381454
rect 82330 380898 82566 381134
rect 113050 381218 113286 381454
rect 113050 380898 113286 381134
rect 143770 381218 144006 381454
rect 143770 380898 144006 381134
rect 174490 381218 174726 381454
rect 174490 380898 174726 381134
rect 205210 381218 205446 381454
rect 205210 380898 205446 381134
rect 235930 381218 236166 381454
rect 235930 380898 236166 381134
rect 266650 381218 266886 381454
rect 266650 380898 266886 381134
rect 297370 381218 297606 381454
rect 297370 380898 297606 381134
rect 328090 381218 328326 381454
rect 328090 380898 328326 381134
rect 358810 381218 359046 381454
rect 358810 380898 359046 381134
rect 389530 381218 389766 381454
rect 389530 380898 389766 381134
rect 420250 381218 420486 381454
rect 420250 380898 420486 381134
rect 450970 381218 451206 381454
rect 450970 380898 451206 381134
rect 481690 381218 481926 381454
rect 481690 380898 481926 381134
rect 512410 381218 512646 381454
rect 512410 380898 512646 381134
rect 543130 381218 543366 381454
rect 543130 380898 543366 381134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 36250 363218 36486 363454
rect 36250 362898 36486 363134
rect 66970 363218 67206 363454
rect 66970 362898 67206 363134
rect 97690 363218 97926 363454
rect 97690 362898 97926 363134
rect 128410 363218 128646 363454
rect 128410 362898 128646 363134
rect 159130 363218 159366 363454
rect 159130 362898 159366 363134
rect 189850 363218 190086 363454
rect 189850 362898 190086 363134
rect 220570 363218 220806 363454
rect 220570 362898 220806 363134
rect 251290 363218 251526 363454
rect 251290 362898 251526 363134
rect 282010 363218 282246 363454
rect 282010 362898 282246 363134
rect 312730 363218 312966 363454
rect 312730 362898 312966 363134
rect 343450 363218 343686 363454
rect 343450 362898 343686 363134
rect 374170 363218 374406 363454
rect 374170 362898 374406 363134
rect 404890 363218 405126 363454
rect 404890 362898 405126 363134
rect 435610 363218 435846 363454
rect 435610 362898 435846 363134
rect 466330 363218 466566 363454
rect 466330 362898 466566 363134
rect 497050 363218 497286 363454
rect 497050 362898 497286 363134
rect 527770 363218 528006 363454
rect 527770 362898 528006 363134
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 51610 345218 51846 345454
rect 51610 344898 51846 345134
rect 82330 345218 82566 345454
rect 82330 344898 82566 345134
rect 113050 345218 113286 345454
rect 113050 344898 113286 345134
rect 143770 345218 144006 345454
rect 143770 344898 144006 345134
rect 174490 345218 174726 345454
rect 174490 344898 174726 345134
rect 205210 345218 205446 345454
rect 205210 344898 205446 345134
rect 235930 345218 236166 345454
rect 235930 344898 236166 345134
rect 266650 345218 266886 345454
rect 266650 344898 266886 345134
rect 297370 345218 297606 345454
rect 297370 344898 297606 345134
rect 328090 345218 328326 345454
rect 328090 344898 328326 345134
rect 358810 345218 359046 345454
rect 358810 344898 359046 345134
rect 389530 345218 389766 345454
rect 389530 344898 389766 345134
rect 420250 345218 420486 345454
rect 420250 344898 420486 345134
rect 450970 345218 451206 345454
rect 450970 344898 451206 345134
rect 481690 345218 481926 345454
rect 481690 344898 481926 345134
rect 512410 345218 512646 345454
rect 512410 344898 512646 345134
rect 543130 345218 543366 345454
rect 543130 344898 543366 345134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 36250 327218 36486 327454
rect 36250 326898 36486 327134
rect 66970 327218 67206 327454
rect 66970 326898 67206 327134
rect 97690 327218 97926 327454
rect 97690 326898 97926 327134
rect 128410 327218 128646 327454
rect 128410 326898 128646 327134
rect 159130 327218 159366 327454
rect 159130 326898 159366 327134
rect 189850 327218 190086 327454
rect 189850 326898 190086 327134
rect 220570 327218 220806 327454
rect 220570 326898 220806 327134
rect 251290 327218 251526 327454
rect 251290 326898 251526 327134
rect 282010 327218 282246 327454
rect 282010 326898 282246 327134
rect 312730 327218 312966 327454
rect 312730 326898 312966 327134
rect 343450 327218 343686 327454
rect 343450 326898 343686 327134
rect 374170 327218 374406 327454
rect 374170 326898 374406 327134
rect 404890 327218 405126 327454
rect 404890 326898 405126 327134
rect 435610 327218 435846 327454
rect 435610 326898 435846 327134
rect 466330 327218 466566 327454
rect 466330 326898 466566 327134
rect 497050 327218 497286 327454
rect 497050 326898 497286 327134
rect 527770 327218 528006 327454
rect 527770 326898 528006 327134
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 51610 309218 51846 309454
rect 51610 308898 51846 309134
rect 82330 309218 82566 309454
rect 82330 308898 82566 309134
rect 113050 309218 113286 309454
rect 113050 308898 113286 309134
rect 143770 309218 144006 309454
rect 143770 308898 144006 309134
rect 174490 309218 174726 309454
rect 174490 308898 174726 309134
rect 205210 309218 205446 309454
rect 205210 308898 205446 309134
rect 235930 309218 236166 309454
rect 235930 308898 236166 309134
rect 266650 309218 266886 309454
rect 266650 308898 266886 309134
rect 297370 309218 297606 309454
rect 297370 308898 297606 309134
rect 328090 309218 328326 309454
rect 328090 308898 328326 309134
rect 358810 309218 359046 309454
rect 358810 308898 359046 309134
rect 389530 309218 389766 309454
rect 389530 308898 389766 309134
rect 420250 309218 420486 309454
rect 420250 308898 420486 309134
rect 450970 309218 451206 309454
rect 450970 308898 451206 309134
rect 481690 309218 481926 309454
rect 481690 308898 481926 309134
rect 512410 309218 512646 309454
rect 512410 308898 512646 309134
rect 543130 309218 543366 309454
rect 543130 308898 543366 309134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 36250 291218 36486 291454
rect 36250 290898 36486 291134
rect 66970 291218 67206 291454
rect 66970 290898 67206 291134
rect 97690 291218 97926 291454
rect 97690 290898 97926 291134
rect 128410 291218 128646 291454
rect 128410 290898 128646 291134
rect 159130 291218 159366 291454
rect 159130 290898 159366 291134
rect 189850 291218 190086 291454
rect 189850 290898 190086 291134
rect 220570 291218 220806 291454
rect 220570 290898 220806 291134
rect 251290 291218 251526 291454
rect 251290 290898 251526 291134
rect 282010 291218 282246 291454
rect 282010 290898 282246 291134
rect 312730 291218 312966 291454
rect 312730 290898 312966 291134
rect 343450 291218 343686 291454
rect 343450 290898 343686 291134
rect 374170 291218 374406 291454
rect 374170 290898 374406 291134
rect 404890 291218 405126 291454
rect 404890 290898 405126 291134
rect 435610 291218 435846 291454
rect 435610 290898 435846 291134
rect 466330 291218 466566 291454
rect 466330 290898 466566 291134
rect 497050 291218 497286 291454
rect 497050 290898 497286 291134
rect 527770 291218 528006 291454
rect 527770 290898 528006 291134
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 51610 273218 51846 273454
rect 51610 272898 51846 273134
rect 82330 273218 82566 273454
rect 82330 272898 82566 273134
rect 113050 273218 113286 273454
rect 113050 272898 113286 273134
rect 143770 273218 144006 273454
rect 143770 272898 144006 273134
rect 174490 273218 174726 273454
rect 174490 272898 174726 273134
rect 205210 273218 205446 273454
rect 205210 272898 205446 273134
rect 235930 273218 236166 273454
rect 235930 272898 236166 273134
rect 266650 273218 266886 273454
rect 266650 272898 266886 273134
rect 297370 273218 297606 273454
rect 297370 272898 297606 273134
rect 328090 273218 328326 273454
rect 328090 272898 328326 273134
rect 358810 273218 359046 273454
rect 358810 272898 359046 273134
rect 389530 273218 389766 273454
rect 389530 272898 389766 273134
rect 420250 273218 420486 273454
rect 420250 272898 420486 273134
rect 450970 273218 451206 273454
rect 450970 272898 451206 273134
rect 481690 273218 481926 273454
rect 481690 272898 481926 273134
rect 512410 273218 512646 273454
rect 512410 272898 512646 273134
rect 543130 273218 543366 273454
rect 543130 272898 543366 273134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 36250 255218 36486 255454
rect 36250 254898 36486 255134
rect 66970 255218 67206 255454
rect 66970 254898 67206 255134
rect 97690 255218 97926 255454
rect 97690 254898 97926 255134
rect 128410 255218 128646 255454
rect 128410 254898 128646 255134
rect 159130 255218 159366 255454
rect 159130 254898 159366 255134
rect 189850 255218 190086 255454
rect 189850 254898 190086 255134
rect 220570 255218 220806 255454
rect 220570 254898 220806 255134
rect 251290 255218 251526 255454
rect 251290 254898 251526 255134
rect 282010 255218 282246 255454
rect 282010 254898 282246 255134
rect 312730 255218 312966 255454
rect 312730 254898 312966 255134
rect 343450 255218 343686 255454
rect 343450 254898 343686 255134
rect 374170 255218 374406 255454
rect 374170 254898 374406 255134
rect 404890 255218 405126 255454
rect 404890 254898 405126 255134
rect 435610 255218 435846 255454
rect 435610 254898 435846 255134
rect 466330 255218 466566 255454
rect 466330 254898 466566 255134
rect 497050 255218 497286 255454
rect 497050 254898 497286 255134
rect 527770 255218 528006 255454
rect 527770 254898 528006 255134
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 51610 237218 51846 237454
rect 51610 236898 51846 237134
rect 82330 237218 82566 237454
rect 82330 236898 82566 237134
rect 113050 237218 113286 237454
rect 113050 236898 113286 237134
rect 143770 237218 144006 237454
rect 143770 236898 144006 237134
rect 174490 237218 174726 237454
rect 174490 236898 174726 237134
rect 205210 237218 205446 237454
rect 205210 236898 205446 237134
rect 235930 237218 236166 237454
rect 235930 236898 236166 237134
rect 266650 237218 266886 237454
rect 266650 236898 266886 237134
rect 297370 237218 297606 237454
rect 297370 236898 297606 237134
rect 328090 237218 328326 237454
rect 328090 236898 328326 237134
rect 358810 237218 359046 237454
rect 358810 236898 359046 237134
rect 389530 237218 389766 237454
rect 389530 236898 389766 237134
rect 420250 237218 420486 237454
rect 420250 236898 420486 237134
rect 450970 237218 451206 237454
rect 450970 236898 451206 237134
rect 481690 237218 481926 237454
rect 481690 236898 481926 237134
rect 512410 237218 512646 237454
rect 512410 236898 512646 237134
rect 543130 237218 543366 237454
rect 543130 236898 543366 237134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 36250 219218 36486 219454
rect 36250 218898 36486 219134
rect 66970 219218 67206 219454
rect 66970 218898 67206 219134
rect 97690 219218 97926 219454
rect 97690 218898 97926 219134
rect 128410 219218 128646 219454
rect 128410 218898 128646 219134
rect 159130 219218 159366 219454
rect 159130 218898 159366 219134
rect 189850 219218 190086 219454
rect 189850 218898 190086 219134
rect 220570 219218 220806 219454
rect 220570 218898 220806 219134
rect 251290 219218 251526 219454
rect 251290 218898 251526 219134
rect 282010 219218 282246 219454
rect 282010 218898 282246 219134
rect 312730 219218 312966 219454
rect 312730 218898 312966 219134
rect 343450 219218 343686 219454
rect 343450 218898 343686 219134
rect 374170 219218 374406 219454
rect 374170 218898 374406 219134
rect 404890 219218 405126 219454
rect 404890 218898 405126 219134
rect 435610 219218 435846 219454
rect 435610 218898 435846 219134
rect 466330 219218 466566 219454
rect 466330 218898 466566 219134
rect 497050 219218 497286 219454
rect 497050 218898 497286 219134
rect 527770 219218 528006 219454
rect 527770 218898 528006 219134
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 51610 201218 51846 201454
rect 51610 200898 51846 201134
rect 82330 201218 82566 201454
rect 82330 200898 82566 201134
rect 113050 201218 113286 201454
rect 113050 200898 113286 201134
rect 143770 201218 144006 201454
rect 143770 200898 144006 201134
rect 174490 201218 174726 201454
rect 174490 200898 174726 201134
rect 205210 201218 205446 201454
rect 205210 200898 205446 201134
rect 235930 201218 236166 201454
rect 235930 200898 236166 201134
rect 266650 201218 266886 201454
rect 266650 200898 266886 201134
rect 297370 201218 297606 201454
rect 297370 200898 297606 201134
rect 328090 201218 328326 201454
rect 328090 200898 328326 201134
rect 358810 201218 359046 201454
rect 358810 200898 359046 201134
rect 389530 201218 389766 201454
rect 389530 200898 389766 201134
rect 420250 201218 420486 201454
rect 420250 200898 420486 201134
rect 450970 201218 451206 201454
rect 450970 200898 451206 201134
rect 481690 201218 481926 201454
rect 481690 200898 481926 201134
rect 512410 201218 512646 201454
rect 512410 200898 512646 201134
rect 543130 201218 543366 201454
rect 543130 200898 543366 201134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 36250 183218 36486 183454
rect 36250 182898 36486 183134
rect 66970 183218 67206 183454
rect 66970 182898 67206 183134
rect 97690 183218 97926 183454
rect 97690 182898 97926 183134
rect 128410 183218 128646 183454
rect 128410 182898 128646 183134
rect 159130 183218 159366 183454
rect 159130 182898 159366 183134
rect 189850 183218 190086 183454
rect 189850 182898 190086 183134
rect 220570 183218 220806 183454
rect 220570 182898 220806 183134
rect 251290 183218 251526 183454
rect 251290 182898 251526 183134
rect 282010 183218 282246 183454
rect 282010 182898 282246 183134
rect 312730 183218 312966 183454
rect 312730 182898 312966 183134
rect 343450 183218 343686 183454
rect 343450 182898 343686 183134
rect 374170 183218 374406 183454
rect 374170 182898 374406 183134
rect 404890 183218 405126 183454
rect 404890 182898 405126 183134
rect 435610 183218 435846 183454
rect 435610 182898 435846 183134
rect 466330 183218 466566 183454
rect 466330 182898 466566 183134
rect 497050 183218 497286 183454
rect 497050 182898 497286 183134
rect 527770 183218 528006 183454
rect 527770 182898 528006 183134
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 51610 165218 51846 165454
rect 51610 164898 51846 165134
rect 82330 165218 82566 165454
rect 82330 164898 82566 165134
rect 113050 165218 113286 165454
rect 113050 164898 113286 165134
rect 143770 165218 144006 165454
rect 143770 164898 144006 165134
rect 174490 165218 174726 165454
rect 174490 164898 174726 165134
rect 205210 165218 205446 165454
rect 205210 164898 205446 165134
rect 235930 165218 236166 165454
rect 235930 164898 236166 165134
rect 266650 165218 266886 165454
rect 266650 164898 266886 165134
rect 297370 165218 297606 165454
rect 297370 164898 297606 165134
rect 328090 165218 328326 165454
rect 328090 164898 328326 165134
rect 358810 165218 359046 165454
rect 358810 164898 359046 165134
rect 389530 165218 389766 165454
rect 389530 164898 389766 165134
rect 420250 165218 420486 165454
rect 420250 164898 420486 165134
rect 450970 165218 451206 165454
rect 450970 164898 451206 165134
rect 481690 165218 481926 165454
rect 481690 164898 481926 165134
rect 512410 165218 512646 165454
rect 512410 164898 512646 165134
rect 543130 165218 543366 165454
rect 543130 164898 543366 165134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 36250 147218 36486 147454
rect 36250 146898 36486 147134
rect 66970 147218 67206 147454
rect 66970 146898 67206 147134
rect 97690 147218 97926 147454
rect 97690 146898 97926 147134
rect 128410 147218 128646 147454
rect 128410 146898 128646 147134
rect 159130 147218 159366 147454
rect 159130 146898 159366 147134
rect 189850 147218 190086 147454
rect 189850 146898 190086 147134
rect 220570 147218 220806 147454
rect 220570 146898 220806 147134
rect 251290 147218 251526 147454
rect 251290 146898 251526 147134
rect 282010 147218 282246 147454
rect 282010 146898 282246 147134
rect 312730 147218 312966 147454
rect 312730 146898 312966 147134
rect 343450 147218 343686 147454
rect 343450 146898 343686 147134
rect 374170 147218 374406 147454
rect 374170 146898 374406 147134
rect 404890 147218 405126 147454
rect 404890 146898 405126 147134
rect 435610 147218 435846 147454
rect 435610 146898 435846 147134
rect 466330 147218 466566 147454
rect 466330 146898 466566 147134
rect 497050 147218 497286 147454
rect 497050 146898 497286 147134
rect 527770 147218 528006 147454
rect 527770 146898 528006 147134
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 51610 129218 51846 129454
rect 51610 128898 51846 129134
rect 82330 129218 82566 129454
rect 82330 128898 82566 129134
rect 113050 129218 113286 129454
rect 113050 128898 113286 129134
rect 143770 129218 144006 129454
rect 143770 128898 144006 129134
rect 174490 129218 174726 129454
rect 174490 128898 174726 129134
rect 205210 129218 205446 129454
rect 205210 128898 205446 129134
rect 235930 129218 236166 129454
rect 235930 128898 236166 129134
rect 266650 129218 266886 129454
rect 266650 128898 266886 129134
rect 297370 129218 297606 129454
rect 297370 128898 297606 129134
rect 328090 129218 328326 129454
rect 328090 128898 328326 129134
rect 358810 129218 359046 129454
rect 358810 128898 359046 129134
rect 389530 129218 389766 129454
rect 389530 128898 389766 129134
rect 420250 129218 420486 129454
rect 420250 128898 420486 129134
rect 450970 129218 451206 129454
rect 450970 128898 451206 129134
rect 481690 129218 481926 129454
rect 481690 128898 481926 129134
rect 512410 129218 512646 129454
rect 512410 128898 512646 129134
rect 543130 129218 543366 129454
rect 543130 128898 543366 129134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 36250 111218 36486 111454
rect 36250 110898 36486 111134
rect 66970 111218 67206 111454
rect 66970 110898 67206 111134
rect 97690 111218 97926 111454
rect 97690 110898 97926 111134
rect 128410 111218 128646 111454
rect 128410 110898 128646 111134
rect 159130 111218 159366 111454
rect 159130 110898 159366 111134
rect 189850 111218 190086 111454
rect 189850 110898 190086 111134
rect 220570 111218 220806 111454
rect 220570 110898 220806 111134
rect 251290 111218 251526 111454
rect 251290 110898 251526 111134
rect 282010 111218 282246 111454
rect 282010 110898 282246 111134
rect 312730 111218 312966 111454
rect 312730 110898 312966 111134
rect 343450 111218 343686 111454
rect 343450 110898 343686 111134
rect 374170 111218 374406 111454
rect 374170 110898 374406 111134
rect 404890 111218 405126 111454
rect 404890 110898 405126 111134
rect 435610 111218 435846 111454
rect 435610 110898 435846 111134
rect 466330 111218 466566 111454
rect 466330 110898 466566 111134
rect 497050 111218 497286 111454
rect 497050 110898 497286 111134
rect 527770 111218 528006 111454
rect 527770 110898 528006 111134
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 51610 93218 51846 93454
rect 51610 92898 51846 93134
rect 82330 93218 82566 93454
rect 82330 92898 82566 93134
rect 113050 93218 113286 93454
rect 113050 92898 113286 93134
rect 143770 93218 144006 93454
rect 143770 92898 144006 93134
rect 174490 93218 174726 93454
rect 174490 92898 174726 93134
rect 205210 93218 205446 93454
rect 205210 92898 205446 93134
rect 235930 93218 236166 93454
rect 235930 92898 236166 93134
rect 266650 93218 266886 93454
rect 266650 92898 266886 93134
rect 297370 93218 297606 93454
rect 297370 92898 297606 93134
rect 328090 93218 328326 93454
rect 328090 92898 328326 93134
rect 358810 93218 359046 93454
rect 358810 92898 359046 93134
rect 389530 93218 389766 93454
rect 389530 92898 389766 93134
rect 420250 93218 420486 93454
rect 420250 92898 420486 93134
rect 450970 93218 451206 93454
rect 450970 92898 451206 93134
rect 481690 93218 481926 93454
rect 481690 92898 481926 93134
rect 512410 93218 512646 93454
rect 512410 92898 512646 93134
rect 543130 93218 543366 93454
rect 543130 92898 543366 93134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 36250 75218 36486 75454
rect 36250 74898 36486 75134
rect 66970 75218 67206 75454
rect 66970 74898 67206 75134
rect 97690 75218 97926 75454
rect 97690 74898 97926 75134
rect 128410 75218 128646 75454
rect 128410 74898 128646 75134
rect 159130 75218 159366 75454
rect 159130 74898 159366 75134
rect 189850 75218 190086 75454
rect 189850 74898 190086 75134
rect 220570 75218 220806 75454
rect 220570 74898 220806 75134
rect 251290 75218 251526 75454
rect 251290 74898 251526 75134
rect 282010 75218 282246 75454
rect 282010 74898 282246 75134
rect 312730 75218 312966 75454
rect 312730 74898 312966 75134
rect 343450 75218 343686 75454
rect 343450 74898 343686 75134
rect 374170 75218 374406 75454
rect 374170 74898 374406 75134
rect 404890 75218 405126 75454
rect 404890 74898 405126 75134
rect 435610 75218 435846 75454
rect 435610 74898 435846 75134
rect 466330 75218 466566 75454
rect 466330 74898 466566 75134
rect 497050 75218 497286 75454
rect 497050 74898 497286 75134
rect 527770 75218 528006 75454
rect 527770 74898 528006 75134
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 51610 57218 51846 57454
rect 51610 56898 51846 57134
rect 82330 57218 82566 57454
rect 82330 56898 82566 57134
rect 113050 57218 113286 57454
rect 113050 56898 113286 57134
rect 143770 57218 144006 57454
rect 143770 56898 144006 57134
rect 174490 57218 174726 57454
rect 174490 56898 174726 57134
rect 205210 57218 205446 57454
rect 205210 56898 205446 57134
rect 235930 57218 236166 57454
rect 235930 56898 236166 57134
rect 266650 57218 266886 57454
rect 266650 56898 266886 57134
rect 297370 57218 297606 57454
rect 297370 56898 297606 57134
rect 328090 57218 328326 57454
rect 328090 56898 328326 57134
rect 358810 57218 359046 57454
rect 358810 56898 359046 57134
rect 389530 57218 389766 57454
rect 389530 56898 389766 57134
rect 420250 57218 420486 57454
rect 420250 56898 420486 57134
rect 450970 57218 451206 57454
rect 450970 56898 451206 57134
rect 481690 57218 481926 57454
rect 481690 56898 481926 57134
rect 512410 57218 512646 57454
rect 512410 56898 512646 57134
rect 543130 57218 543366 57454
rect 543130 56898 543366 57134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 36250 39218 36486 39454
rect 36250 38898 36486 39134
rect 66970 39218 67206 39454
rect 66970 38898 67206 39134
rect 97690 39218 97926 39454
rect 97690 38898 97926 39134
rect 128410 39218 128646 39454
rect 128410 38898 128646 39134
rect 159130 39218 159366 39454
rect 159130 38898 159366 39134
rect 189850 39218 190086 39454
rect 189850 38898 190086 39134
rect 220570 39218 220806 39454
rect 220570 38898 220806 39134
rect 251290 39218 251526 39454
rect 251290 38898 251526 39134
rect 282010 39218 282246 39454
rect 282010 38898 282246 39134
rect 312730 39218 312966 39454
rect 312730 38898 312966 39134
rect 343450 39218 343686 39454
rect 343450 38898 343686 39134
rect 374170 39218 374406 39454
rect 374170 38898 374406 39134
rect 404890 39218 405126 39454
rect 404890 38898 405126 39134
rect 435610 39218 435846 39454
rect 435610 38898 435846 39134
rect 466330 39218 466566 39454
rect 466330 38898 466566 39134
rect 497050 39218 497286 39454
rect 497050 38898 497286 39134
rect 527770 39218 528006 39454
rect 527770 38898 528006 39134
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 51610 669454
rect 51846 669218 82330 669454
rect 82566 669218 113050 669454
rect 113286 669218 143770 669454
rect 144006 669218 174490 669454
rect 174726 669218 205210 669454
rect 205446 669218 235930 669454
rect 236166 669218 266650 669454
rect 266886 669218 297370 669454
rect 297606 669218 328090 669454
rect 328326 669218 358810 669454
rect 359046 669218 389530 669454
rect 389766 669218 420250 669454
rect 420486 669218 450970 669454
rect 451206 669218 481690 669454
rect 481926 669218 512410 669454
rect 512646 669218 543130 669454
rect 543366 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 51610 669134
rect 51846 668898 82330 669134
rect 82566 668898 113050 669134
rect 113286 668898 143770 669134
rect 144006 668898 174490 669134
rect 174726 668898 205210 669134
rect 205446 668898 235930 669134
rect 236166 668898 266650 669134
rect 266886 668898 297370 669134
rect 297606 668898 328090 669134
rect 328326 668898 358810 669134
rect 359046 668898 389530 669134
rect 389766 668898 420250 669134
rect 420486 668898 450970 669134
rect 451206 668898 481690 669134
rect 481926 668898 512410 669134
rect 512646 668898 543130 669134
rect 543366 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 36250 651454
rect 36486 651218 66970 651454
rect 67206 651218 97690 651454
rect 97926 651218 128410 651454
rect 128646 651218 159130 651454
rect 159366 651218 189850 651454
rect 190086 651218 220570 651454
rect 220806 651218 251290 651454
rect 251526 651218 282010 651454
rect 282246 651218 312730 651454
rect 312966 651218 343450 651454
rect 343686 651218 374170 651454
rect 374406 651218 404890 651454
rect 405126 651218 435610 651454
rect 435846 651218 466330 651454
rect 466566 651218 497050 651454
rect 497286 651218 527770 651454
rect 528006 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 36250 651134
rect 36486 650898 66970 651134
rect 67206 650898 97690 651134
rect 97926 650898 128410 651134
rect 128646 650898 159130 651134
rect 159366 650898 189850 651134
rect 190086 650898 220570 651134
rect 220806 650898 251290 651134
rect 251526 650898 282010 651134
rect 282246 650898 312730 651134
rect 312966 650898 343450 651134
rect 343686 650898 374170 651134
rect 374406 650898 404890 651134
rect 405126 650898 435610 651134
rect 435846 650898 466330 651134
rect 466566 650898 497050 651134
rect 497286 650898 527770 651134
rect 528006 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 51610 633454
rect 51846 633218 82330 633454
rect 82566 633218 113050 633454
rect 113286 633218 143770 633454
rect 144006 633218 174490 633454
rect 174726 633218 205210 633454
rect 205446 633218 235930 633454
rect 236166 633218 266650 633454
rect 266886 633218 297370 633454
rect 297606 633218 328090 633454
rect 328326 633218 358810 633454
rect 359046 633218 389530 633454
rect 389766 633218 420250 633454
rect 420486 633218 450970 633454
rect 451206 633218 481690 633454
rect 481926 633218 512410 633454
rect 512646 633218 543130 633454
rect 543366 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 51610 633134
rect 51846 632898 82330 633134
rect 82566 632898 113050 633134
rect 113286 632898 143770 633134
rect 144006 632898 174490 633134
rect 174726 632898 205210 633134
rect 205446 632898 235930 633134
rect 236166 632898 266650 633134
rect 266886 632898 297370 633134
rect 297606 632898 328090 633134
rect 328326 632898 358810 633134
rect 359046 632898 389530 633134
rect 389766 632898 420250 633134
rect 420486 632898 450970 633134
rect 451206 632898 481690 633134
rect 481926 632898 512410 633134
rect 512646 632898 543130 633134
rect 543366 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 36250 615454
rect 36486 615218 66970 615454
rect 67206 615218 97690 615454
rect 97926 615218 128410 615454
rect 128646 615218 159130 615454
rect 159366 615218 189850 615454
rect 190086 615218 220570 615454
rect 220806 615218 251290 615454
rect 251526 615218 282010 615454
rect 282246 615218 312730 615454
rect 312966 615218 343450 615454
rect 343686 615218 374170 615454
rect 374406 615218 404890 615454
rect 405126 615218 435610 615454
rect 435846 615218 466330 615454
rect 466566 615218 497050 615454
rect 497286 615218 527770 615454
rect 528006 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 36250 615134
rect 36486 614898 66970 615134
rect 67206 614898 97690 615134
rect 97926 614898 128410 615134
rect 128646 614898 159130 615134
rect 159366 614898 189850 615134
rect 190086 614898 220570 615134
rect 220806 614898 251290 615134
rect 251526 614898 282010 615134
rect 282246 614898 312730 615134
rect 312966 614898 343450 615134
rect 343686 614898 374170 615134
rect 374406 614898 404890 615134
rect 405126 614898 435610 615134
rect 435846 614898 466330 615134
rect 466566 614898 497050 615134
rect 497286 614898 527770 615134
rect 528006 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 51610 597454
rect 51846 597218 82330 597454
rect 82566 597218 113050 597454
rect 113286 597218 143770 597454
rect 144006 597218 174490 597454
rect 174726 597218 205210 597454
rect 205446 597218 235930 597454
rect 236166 597218 266650 597454
rect 266886 597218 297370 597454
rect 297606 597218 328090 597454
rect 328326 597218 358810 597454
rect 359046 597218 389530 597454
rect 389766 597218 420250 597454
rect 420486 597218 450970 597454
rect 451206 597218 481690 597454
rect 481926 597218 512410 597454
rect 512646 597218 543130 597454
rect 543366 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 51610 597134
rect 51846 596898 82330 597134
rect 82566 596898 113050 597134
rect 113286 596898 143770 597134
rect 144006 596898 174490 597134
rect 174726 596898 205210 597134
rect 205446 596898 235930 597134
rect 236166 596898 266650 597134
rect 266886 596898 297370 597134
rect 297606 596898 328090 597134
rect 328326 596898 358810 597134
rect 359046 596898 389530 597134
rect 389766 596898 420250 597134
rect 420486 596898 450970 597134
rect 451206 596898 481690 597134
rect 481926 596898 512410 597134
rect 512646 596898 543130 597134
rect 543366 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 36250 579454
rect 36486 579218 66970 579454
rect 67206 579218 97690 579454
rect 97926 579218 128410 579454
rect 128646 579218 159130 579454
rect 159366 579218 189850 579454
rect 190086 579218 220570 579454
rect 220806 579218 251290 579454
rect 251526 579218 282010 579454
rect 282246 579218 312730 579454
rect 312966 579218 343450 579454
rect 343686 579218 374170 579454
rect 374406 579218 404890 579454
rect 405126 579218 435610 579454
rect 435846 579218 466330 579454
rect 466566 579218 497050 579454
rect 497286 579218 527770 579454
rect 528006 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 36250 579134
rect 36486 578898 66970 579134
rect 67206 578898 97690 579134
rect 97926 578898 128410 579134
rect 128646 578898 159130 579134
rect 159366 578898 189850 579134
rect 190086 578898 220570 579134
rect 220806 578898 251290 579134
rect 251526 578898 282010 579134
rect 282246 578898 312730 579134
rect 312966 578898 343450 579134
rect 343686 578898 374170 579134
rect 374406 578898 404890 579134
rect 405126 578898 435610 579134
rect 435846 578898 466330 579134
rect 466566 578898 497050 579134
rect 497286 578898 527770 579134
rect 528006 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 51610 561454
rect 51846 561218 82330 561454
rect 82566 561218 113050 561454
rect 113286 561218 143770 561454
rect 144006 561218 174490 561454
rect 174726 561218 205210 561454
rect 205446 561218 235930 561454
rect 236166 561218 266650 561454
rect 266886 561218 297370 561454
rect 297606 561218 328090 561454
rect 328326 561218 358810 561454
rect 359046 561218 389530 561454
rect 389766 561218 420250 561454
rect 420486 561218 450970 561454
rect 451206 561218 481690 561454
rect 481926 561218 512410 561454
rect 512646 561218 543130 561454
rect 543366 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 51610 561134
rect 51846 560898 82330 561134
rect 82566 560898 113050 561134
rect 113286 560898 143770 561134
rect 144006 560898 174490 561134
rect 174726 560898 205210 561134
rect 205446 560898 235930 561134
rect 236166 560898 266650 561134
rect 266886 560898 297370 561134
rect 297606 560898 328090 561134
rect 328326 560898 358810 561134
rect 359046 560898 389530 561134
rect 389766 560898 420250 561134
rect 420486 560898 450970 561134
rect 451206 560898 481690 561134
rect 481926 560898 512410 561134
rect 512646 560898 543130 561134
rect 543366 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 36250 543454
rect 36486 543218 66970 543454
rect 67206 543218 97690 543454
rect 97926 543218 128410 543454
rect 128646 543218 159130 543454
rect 159366 543218 189850 543454
rect 190086 543218 220570 543454
rect 220806 543218 251290 543454
rect 251526 543218 282010 543454
rect 282246 543218 312730 543454
rect 312966 543218 343450 543454
rect 343686 543218 374170 543454
rect 374406 543218 404890 543454
rect 405126 543218 435610 543454
rect 435846 543218 466330 543454
rect 466566 543218 497050 543454
rect 497286 543218 527770 543454
rect 528006 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 36250 543134
rect 36486 542898 66970 543134
rect 67206 542898 97690 543134
rect 97926 542898 128410 543134
rect 128646 542898 159130 543134
rect 159366 542898 189850 543134
rect 190086 542898 220570 543134
rect 220806 542898 251290 543134
rect 251526 542898 282010 543134
rect 282246 542898 312730 543134
rect 312966 542898 343450 543134
rect 343686 542898 374170 543134
rect 374406 542898 404890 543134
rect 405126 542898 435610 543134
rect 435846 542898 466330 543134
rect 466566 542898 497050 543134
rect 497286 542898 527770 543134
rect 528006 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 51610 525454
rect 51846 525218 82330 525454
rect 82566 525218 113050 525454
rect 113286 525218 143770 525454
rect 144006 525218 174490 525454
rect 174726 525218 205210 525454
rect 205446 525218 235930 525454
rect 236166 525218 266650 525454
rect 266886 525218 297370 525454
rect 297606 525218 328090 525454
rect 328326 525218 358810 525454
rect 359046 525218 389530 525454
rect 389766 525218 420250 525454
rect 420486 525218 450970 525454
rect 451206 525218 481690 525454
rect 481926 525218 512410 525454
rect 512646 525218 543130 525454
rect 543366 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 51610 525134
rect 51846 524898 82330 525134
rect 82566 524898 113050 525134
rect 113286 524898 143770 525134
rect 144006 524898 174490 525134
rect 174726 524898 205210 525134
rect 205446 524898 235930 525134
rect 236166 524898 266650 525134
rect 266886 524898 297370 525134
rect 297606 524898 328090 525134
rect 328326 524898 358810 525134
rect 359046 524898 389530 525134
rect 389766 524898 420250 525134
rect 420486 524898 450970 525134
rect 451206 524898 481690 525134
rect 481926 524898 512410 525134
rect 512646 524898 543130 525134
rect 543366 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 36250 507454
rect 36486 507218 66970 507454
rect 67206 507218 97690 507454
rect 97926 507218 128410 507454
rect 128646 507218 159130 507454
rect 159366 507218 189850 507454
rect 190086 507218 220570 507454
rect 220806 507218 251290 507454
rect 251526 507218 282010 507454
rect 282246 507218 312730 507454
rect 312966 507218 343450 507454
rect 343686 507218 374170 507454
rect 374406 507218 404890 507454
rect 405126 507218 435610 507454
rect 435846 507218 466330 507454
rect 466566 507218 497050 507454
rect 497286 507218 527770 507454
rect 528006 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 36250 507134
rect 36486 506898 66970 507134
rect 67206 506898 97690 507134
rect 97926 506898 128410 507134
rect 128646 506898 159130 507134
rect 159366 506898 189850 507134
rect 190086 506898 220570 507134
rect 220806 506898 251290 507134
rect 251526 506898 282010 507134
rect 282246 506898 312730 507134
rect 312966 506898 343450 507134
rect 343686 506898 374170 507134
rect 374406 506898 404890 507134
rect 405126 506898 435610 507134
rect 435846 506898 466330 507134
rect 466566 506898 497050 507134
rect 497286 506898 527770 507134
rect 528006 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 51610 489454
rect 51846 489218 82330 489454
rect 82566 489218 113050 489454
rect 113286 489218 143770 489454
rect 144006 489218 174490 489454
rect 174726 489218 205210 489454
rect 205446 489218 235930 489454
rect 236166 489218 266650 489454
rect 266886 489218 297370 489454
rect 297606 489218 328090 489454
rect 328326 489218 358810 489454
rect 359046 489218 389530 489454
rect 389766 489218 420250 489454
rect 420486 489218 450970 489454
rect 451206 489218 481690 489454
rect 481926 489218 512410 489454
rect 512646 489218 543130 489454
rect 543366 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 51610 489134
rect 51846 488898 82330 489134
rect 82566 488898 113050 489134
rect 113286 488898 143770 489134
rect 144006 488898 174490 489134
rect 174726 488898 205210 489134
rect 205446 488898 235930 489134
rect 236166 488898 266650 489134
rect 266886 488898 297370 489134
rect 297606 488898 328090 489134
rect 328326 488898 358810 489134
rect 359046 488898 389530 489134
rect 389766 488898 420250 489134
rect 420486 488898 450970 489134
rect 451206 488898 481690 489134
rect 481926 488898 512410 489134
rect 512646 488898 543130 489134
rect 543366 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 36250 471454
rect 36486 471218 66970 471454
rect 67206 471218 97690 471454
rect 97926 471218 128410 471454
rect 128646 471218 159130 471454
rect 159366 471218 189850 471454
rect 190086 471218 220570 471454
rect 220806 471218 251290 471454
rect 251526 471218 282010 471454
rect 282246 471218 312730 471454
rect 312966 471218 343450 471454
rect 343686 471218 374170 471454
rect 374406 471218 404890 471454
rect 405126 471218 435610 471454
rect 435846 471218 466330 471454
rect 466566 471218 497050 471454
rect 497286 471218 527770 471454
rect 528006 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 36250 471134
rect 36486 470898 66970 471134
rect 67206 470898 97690 471134
rect 97926 470898 128410 471134
rect 128646 470898 159130 471134
rect 159366 470898 189850 471134
rect 190086 470898 220570 471134
rect 220806 470898 251290 471134
rect 251526 470898 282010 471134
rect 282246 470898 312730 471134
rect 312966 470898 343450 471134
rect 343686 470898 374170 471134
rect 374406 470898 404890 471134
rect 405126 470898 435610 471134
rect 435846 470898 466330 471134
rect 466566 470898 497050 471134
rect 497286 470898 527770 471134
rect 528006 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 51610 453454
rect 51846 453218 82330 453454
rect 82566 453218 113050 453454
rect 113286 453218 143770 453454
rect 144006 453218 174490 453454
rect 174726 453218 205210 453454
rect 205446 453218 235930 453454
rect 236166 453218 266650 453454
rect 266886 453218 297370 453454
rect 297606 453218 328090 453454
rect 328326 453218 358810 453454
rect 359046 453218 389530 453454
rect 389766 453218 420250 453454
rect 420486 453218 450970 453454
rect 451206 453218 481690 453454
rect 481926 453218 512410 453454
rect 512646 453218 543130 453454
rect 543366 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 51610 453134
rect 51846 452898 82330 453134
rect 82566 452898 113050 453134
rect 113286 452898 143770 453134
rect 144006 452898 174490 453134
rect 174726 452898 205210 453134
rect 205446 452898 235930 453134
rect 236166 452898 266650 453134
rect 266886 452898 297370 453134
rect 297606 452898 328090 453134
rect 328326 452898 358810 453134
rect 359046 452898 389530 453134
rect 389766 452898 420250 453134
rect 420486 452898 450970 453134
rect 451206 452898 481690 453134
rect 481926 452898 512410 453134
rect 512646 452898 543130 453134
rect 543366 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 36250 435454
rect 36486 435218 66970 435454
rect 67206 435218 97690 435454
rect 97926 435218 128410 435454
rect 128646 435218 159130 435454
rect 159366 435218 189850 435454
rect 190086 435218 220570 435454
rect 220806 435218 251290 435454
rect 251526 435218 282010 435454
rect 282246 435218 312730 435454
rect 312966 435218 343450 435454
rect 343686 435218 374170 435454
rect 374406 435218 404890 435454
rect 405126 435218 435610 435454
rect 435846 435218 466330 435454
rect 466566 435218 497050 435454
rect 497286 435218 527770 435454
rect 528006 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 36250 435134
rect 36486 434898 66970 435134
rect 67206 434898 97690 435134
rect 97926 434898 128410 435134
rect 128646 434898 159130 435134
rect 159366 434898 189850 435134
rect 190086 434898 220570 435134
rect 220806 434898 251290 435134
rect 251526 434898 282010 435134
rect 282246 434898 312730 435134
rect 312966 434898 343450 435134
rect 343686 434898 374170 435134
rect 374406 434898 404890 435134
rect 405126 434898 435610 435134
rect 435846 434898 466330 435134
rect 466566 434898 497050 435134
rect 497286 434898 527770 435134
rect 528006 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 51610 417454
rect 51846 417218 82330 417454
rect 82566 417218 113050 417454
rect 113286 417218 143770 417454
rect 144006 417218 174490 417454
rect 174726 417218 205210 417454
rect 205446 417218 235930 417454
rect 236166 417218 266650 417454
rect 266886 417218 297370 417454
rect 297606 417218 328090 417454
rect 328326 417218 358810 417454
rect 359046 417218 389530 417454
rect 389766 417218 420250 417454
rect 420486 417218 450970 417454
rect 451206 417218 481690 417454
rect 481926 417218 512410 417454
rect 512646 417218 543130 417454
rect 543366 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 51610 417134
rect 51846 416898 82330 417134
rect 82566 416898 113050 417134
rect 113286 416898 143770 417134
rect 144006 416898 174490 417134
rect 174726 416898 205210 417134
rect 205446 416898 235930 417134
rect 236166 416898 266650 417134
rect 266886 416898 297370 417134
rect 297606 416898 328090 417134
rect 328326 416898 358810 417134
rect 359046 416898 389530 417134
rect 389766 416898 420250 417134
rect 420486 416898 450970 417134
rect 451206 416898 481690 417134
rect 481926 416898 512410 417134
rect 512646 416898 543130 417134
rect 543366 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 36250 399454
rect 36486 399218 66970 399454
rect 67206 399218 97690 399454
rect 97926 399218 128410 399454
rect 128646 399218 159130 399454
rect 159366 399218 189850 399454
rect 190086 399218 220570 399454
rect 220806 399218 251290 399454
rect 251526 399218 282010 399454
rect 282246 399218 312730 399454
rect 312966 399218 343450 399454
rect 343686 399218 374170 399454
rect 374406 399218 404890 399454
rect 405126 399218 435610 399454
rect 435846 399218 466330 399454
rect 466566 399218 497050 399454
rect 497286 399218 527770 399454
rect 528006 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 36250 399134
rect 36486 398898 66970 399134
rect 67206 398898 97690 399134
rect 97926 398898 128410 399134
rect 128646 398898 159130 399134
rect 159366 398898 189850 399134
rect 190086 398898 220570 399134
rect 220806 398898 251290 399134
rect 251526 398898 282010 399134
rect 282246 398898 312730 399134
rect 312966 398898 343450 399134
rect 343686 398898 374170 399134
rect 374406 398898 404890 399134
rect 405126 398898 435610 399134
rect 435846 398898 466330 399134
rect 466566 398898 497050 399134
rect 497286 398898 527770 399134
rect 528006 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 51610 381454
rect 51846 381218 82330 381454
rect 82566 381218 113050 381454
rect 113286 381218 143770 381454
rect 144006 381218 174490 381454
rect 174726 381218 205210 381454
rect 205446 381218 235930 381454
rect 236166 381218 266650 381454
rect 266886 381218 297370 381454
rect 297606 381218 328090 381454
rect 328326 381218 358810 381454
rect 359046 381218 389530 381454
rect 389766 381218 420250 381454
rect 420486 381218 450970 381454
rect 451206 381218 481690 381454
rect 481926 381218 512410 381454
rect 512646 381218 543130 381454
rect 543366 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 51610 381134
rect 51846 380898 82330 381134
rect 82566 380898 113050 381134
rect 113286 380898 143770 381134
rect 144006 380898 174490 381134
rect 174726 380898 205210 381134
rect 205446 380898 235930 381134
rect 236166 380898 266650 381134
rect 266886 380898 297370 381134
rect 297606 380898 328090 381134
rect 328326 380898 358810 381134
rect 359046 380898 389530 381134
rect 389766 380898 420250 381134
rect 420486 380898 450970 381134
rect 451206 380898 481690 381134
rect 481926 380898 512410 381134
rect 512646 380898 543130 381134
rect 543366 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 36250 363454
rect 36486 363218 66970 363454
rect 67206 363218 97690 363454
rect 97926 363218 128410 363454
rect 128646 363218 159130 363454
rect 159366 363218 189850 363454
rect 190086 363218 220570 363454
rect 220806 363218 251290 363454
rect 251526 363218 282010 363454
rect 282246 363218 312730 363454
rect 312966 363218 343450 363454
rect 343686 363218 374170 363454
rect 374406 363218 404890 363454
rect 405126 363218 435610 363454
rect 435846 363218 466330 363454
rect 466566 363218 497050 363454
rect 497286 363218 527770 363454
rect 528006 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 36250 363134
rect 36486 362898 66970 363134
rect 67206 362898 97690 363134
rect 97926 362898 128410 363134
rect 128646 362898 159130 363134
rect 159366 362898 189850 363134
rect 190086 362898 220570 363134
rect 220806 362898 251290 363134
rect 251526 362898 282010 363134
rect 282246 362898 312730 363134
rect 312966 362898 343450 363134
rect 343686 362898 374170 363134
rect 374406 362898 404890 363134
rect 405126 362898 435610 363134
rect 435846 362898 466330 363134
rect 466566 362898 497050 363134
rect 497286 362898 527770 363134
rect 528006 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 51610 345454
rect 51846 345218 82330 345454
rect 82566 345218 113050 345454
rect 113286 345218 143770 345454
rect 144006 345218 174490 345454
rect 174726 345218 205210 345454
rect 205446 345218 235930 345454
rect 236166 345218 266650 345454
rect 266886 345218 297370 345454
rect 297606 345218 328090 345454
rect 328326 345218 358810 345454
rect 359046 345218 389530 345454
rect 389766 345218 420250 345454
rect 420486 345218 450970 345454
rect 451206 345218 481690 345454
rect 481926 345218 512410 345454
rect 512646 345218 543130 345454
rect 543366 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 51610 345134
rect 51846 344898 82330 345134
rect 82566 344898 113050 345134
rect 113286 344898 143770 345134
rect 144006 344898 174490 345134
rect 174726 344898 205210 345134
rect 205446 344898 235930 345134
rect 236166 344898 266650 345134
rect 266886 344898 297370 345134
rect 297606 344898 328090 345134
rect 328326 344898 358810 345134
rect 359046 344898 389530 345134
rect 389766 344898 420250 345134
rect 420486 344898 450970 345134
rect 451206 344898 481690 345134
rect 481926 344898 512410 345134
rect 512646 344898 543130 345134
rect 543366 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 36250 327454
rect 36486 327218 66970 327454
rect 67206 327218 97690 327454
rect 97926 327218 128410 327454
rect 128646 327218 159130 327454
rect 159366 327218 189850 327454
rect 190086 327218 220570 327454
rect 220806 327218 251290 327454
rect 251526 327218 282010 327454
rect 282246 327218 312730 327454
rect 312966 327218 343450 327454
rect 343686 327218 374170 327454
rect 374406 327218 404890 327454
rect 405126 327218 435610 327454
rect 435846 327218 466330 327454
rect 466566 327218 497050 327454
rect 497286 327218 527770 327454
rect 528006 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 36250 327134
rect 36486 326898 66970 327134
rect 67206 326898 97690 327134
rect 97926 326898 128410 327134
rect 128646 326898 159130 327134
rect 159366 326898 189850 327134
rect 190086 326898 220570 327134
rect 220806 326898 251290 327134
rect 251526 326898 282010 327134
rect 282246 326898 312730 327134
rect 312966 326898 343450 327134
rect 343686 326898 374170 327134
rect 374406 326898 404890 327134
rect 405126 326898 435610 327134
rect 435846 326898 466330 327134
rect 466566 326898 497050 327134
rect 497286 326898 527770 327134
rect 528006 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 51610 309454
rect 51846 309218 82330 309454
rect 82566 309218 113050 309454
rect 113286 309218 143770 309454
rect 144006 309218 174490 309454
rect 174726 309218 205210 309454
rect 205446 309218 235930 309454
rect 236166 309218 266650 309454
rect 266886 309218 297370 309454
rect 297606 309218 328090 309454
rect 328326 309218 358810 309454
rect 359046 309218 389530 309454
rect 389766 309218 420250 309454
rect 420486 309218 450970 309454
rect 451206 309218 481690 309454
rect 481926 309218 512410 309454
rect 512646 309218 543130 309454
rect 543366 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 51610 309134
rect 51846 308898 82330 309134
rect 82566 308898 113050 309134
rect 113286 308898 143770 309134
rect 144006 308898 174490 309134
rect 174726 308898 205210 309134
rect 205446 308898 235930 309134
rect 236166 308898 266650 309134
rect 266886 308898 297370 309134
rect 297606 308898 328090 309134
rect 328326 308898 358810 309134
rect 359046 308898 389530 309134
rect 389766 308898 420250 309134
rect 420486 308898 450970 309134
rect 451206 308898 481690 309134
rect 481926 308898 512410 309134
rect 512646 308898 543130 309134
rect 543366 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 36250 291454
rect 36486 291218 66970 291454
rect 67206 291218 97690 291454
rect 97926 291218 128410 291454
rect 128646 291218 159130 291454
rect 159366 291218 189850 291454
rect 190086 291218 220570 291454
rect 220806 291218 251290 291454
rect 251526 291218 282010 291454
rect 282246 291218 312730 291454
rect 312966 291218 343450 291454
rect 343686 291218 374170 291454
rect 374406 291218 404890 291454
rect 405126 291218 435610 291454
rect 435846 291218 466330 291454
rect 466566 291218 497050 291454
rect 497286 291218 527770 291454
rect 528006 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 36250 291134
rect 36486 290898 66970 291134
rect 67206 290898 97690 291134
rect 97926 290898 128410 291134
rect 128646 290898 159130 291134
rect 159366 290898 189850 291134
rect 190086 290898 220570 291134
rect 220806 290898 251290 291134
rect 251526 290898 282010 291134
rect 282246 290898 312730 291134
rect 312966 290898 343450 291134
rect 343686 290898 374170 291134
rect 374406 290898 404890 291134
rect 405126 290898 435610 291134
rect 435846 290898 466330 291134
rect 466566 290898 497050 291134
rect 497286 290898 527770 291134
rect 528006 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 51610 273454
rect 51846 273218 82330 273454
rect 82566 273218 113050 273454
rect 113286 273218 143770 273454
rect 144006 273218 174490 273454
rect 174726 273218 205210 273454
rect 205446 273218 235930 273454
rect 236166 273218 266650 273454
rect 266886 273218 297370 273454
rect 297606 273218 328090 273454
rect 328326 273218 358810 273454
rect 359046 273218 389530 273454
rect 389766 273218 420250 273454
rect 420486 273218 450970 273454
rect 451206 273218 481690 273454
rect 481926 273218 512410 273454
rect 512646 273218 543130 273454
rect 543366 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 51610 273134
rect 51846 272898 82330 273134
rect 82566 272898 113050 273134
rect 113286 272898 143770 273134
rect 144006 272898 174490 273134
rect 174726 272898 205210 273134
rect 205446 272898 235930 273134
rect 236166 272898 266650 273134
rect 266886 272898 297370 273134
rect 297606 272898 328090 273134
rect 328326 272898 358810 273134
rect 359046 272898 389530 273134
rect 389766 272898 420250 273134
rect 420486 272898 450970 273134
rect 451206 272898 481690 273134
rect 481926 272898 512410 273134
rect 512646 272898 543130 273134
rect 543366 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 36250 255454
rect 36486 255218 66970 255454
rect 67206 255218 97690 255454
rect 97926 255218 128410 255454
rect 128646 255218 159130 255454
rect 159366 255218 189850 255454
rect 190086 255218 220570 255454
rect 220806 255218 251290 255454
rect 251526 255218 282010 255454
rect 282246 255218 312730 255454
rect 312966 255218 343450 255454
rect 343686 255218 374170 255454
rect 374406 255218 404890 255454
rect 405126 255218 435610 255454
rect 435846 255218 466330 255454
rect 466566 255218 497050 255454
rect 497286 255218 527770 255454
rect 528006 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 36250 255134
rect 36486 254898 66970 255134
rect 67206 254898 97690 255134
rect 97926 254898 128410 255134
rect 128646 254898 159130 255134
rect 159366 254898 189850 255134
rect 190086 254898 220570 255134
rect 220806 254898 251290 255134
rect 251526 254898 282010 255134
rect 282246 254898 312730 255134
rect 312966 254898 343450 255134
rect 343686 254898 374170 255134
rect 374406 254898 404890 255134
rect 405126 254898 435610 255134
rect 435846 254898 466330 255134
rect 466566 254898 497050 255134
rect 497286 254898 527770 255134
rect 528006 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 51610 237454
rect 51846 237218 82330 237454
rect 82566 237218 113050 237454
rect 113286 237218 143770 237454
rect 144006 237218 174490 237454
rect 174726 237218 205210 237454
rect 205446 237218 235930 237454
rect 236166 237218 266650 237454
rect 266886 237218 297370 237454
rect 297606 237218 328090 237454
rect 328326 237218 358810 237454
rect 359046 237218 389530 237454
rect 389766 237218 420250 237454
rect 420486 237218 450970 237454
rect 451206 237218 481690 237454
rect 481926 237218 512410 237454
rect 512646 237218 543130 237454
rect 543366 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 51610 237134
rect 51846 236898 82330 237134
rect 82566 236898 113050 237134
rect 113286 236898 143770 237134
rect 144006 236898 174490 237134
rect 174726 236898 205210 237134
rect 205446 236898 235930 237134
rect 236166 236898 266650 237134
rect 266886 236898 297370 237134
rect 297606 236898 328090 237134
rect 328326 236898 358810 237134
rect 359046 236898 389530 237134
rect 389766 236898 420250 237134
rect 420486 236898 450970 237134
rect 451206 236898 481690 237134
rect 481926 236898 512410 237134
rect 512646 236898 543130 237134
rect 543366 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 36250 219454
rect 36486 219218 66970 219454
rect 67206 219218 97690 219454
rect 97926 219218 128410 219454
rect 128646 219218 159130 219454
rect 159366 219218 189850 219454
rect 190086 219218 220570 219454
rect 220806 219218 251290 219454
rect 251526 219218 282010 219454
rect 282246 219218 312730 219454
rect 312966 219218 343450 219454
rect 343686 219218 374170 219454
rect 374406 219218 404890 219454
rect 405126 219218 435610 219454
rect 435846 219218 466330 219454
rect 466566 219218 497050 219454
rect 497286 219218 527770 219454
rect 528006 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 36250 219134
rect 36486 218898 66970 219134
rect 67206 218898 97690 219134
rect 97926 218898 128410 219134
rect 128646 218898 159130 219134
rect 159366 218898 189850 219134
rect 190086 218898 220570 219134
rect 220806 218898 251290 219134
rect 251526 218898 282010 219134
rect 282246 218898 312730 219134
rect 312966 218898 343450 219134
rect 343686 218898 374170 219134
rect 374406 218898 404890 219134
rect 405126 218898 435610 219134
rect 435846 218898 466330 219134
rect 466566 218898 497050 219134
rect 497286 218898 527770 219134
rect 528006 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 51610 201454
rect 51846 201218 82330 201454
rect 82566 201218 113050 201454
rect 113286 201218 143770 201454
rect 144006 201218 174490 201454
rect 174726 201218 205210 201454
rect 205446 201218 235930 201454
rect 236166 201218 266650 201454
rect 266886 201218 297370 201454
rect 297606 201218 328090 201454
rect 328326 201218 358810 201454
rect 359046 201218 389530 201454
rect 389766 201218 420250 201454
rect 420486 201218 450970 201454
rect 451206 201218 481690 201454
rect 481926 201218 512410 201454
rect 512646 201218 543130 201454
rect 543366 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 51610 201134
rect 51846 200898 82330 201134
rect 82566 200898 113050 201134
rect 113286 200898 143770 201134
rect 144006 200898 174490 201134
rect 174726 200898 205210 201134
rect 205446 200898 235930 201134
rect 236166 200898 266650 201134
rect 266886 200898 297370 201134
rect 297606 200898 328090 201134
rect 328326 200898 358810 201134
rect 359046 200898 389530 201134
rect 389766 200898 420250 201134
rect 420486 200898 450970 201134
rect 451206 200898 481690 201134
rect 481926 200898 512410 201134
rect 512646 200898 543130 201134
rect 543366 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 36250 183454
rect 36486 183218 66970 183454
rect 67206 183218 97690 183454
rect 97926 183218 128410 183454
rect 128646 183218 159130 183454
rect 159366 183218 189850 183454
rect 190086 183218 220570 183454
rect 220806 183218 251290 183454
rect 251526 183218 282010 183454
rect 282246 183218 312730 183454
rect 312966 183218 343450 183454
rect 343686 183218 374170 183454
rect 374406 183218 404890 183454
rect 405126 183218 435610 183454
rect 435846 183218 466330 183454
rect 466566 183218 497050 183454
rect 497286 183218 527770 183454
rect 528006 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 36250 183134
rect 36486 182898 66970 183134
rect 67206 182898 97690 183134
rect 97926 182898 128410 183134
rect 128646 182898 159130 183134
rect 159366 182898 189850 183134
rect 190086 182898 220570 183134
rect 220806 182898 251290 183134
rect 251526 182898 282010 183134
rect 282246 182898 312730 183134
rect 312966 182898 343450 183134
rect 343686 182898 374170 183134
rect 374406 182898 404890 183134
rect 405126 182898 435610 183134
rect 435846 182898 466330 183134
rect 466566 182898 497050 183134
rect 497286 182898 527770 183134
rect 528006 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 51610 165454
rect 51846 165218 82330 165454
rect 82566 165218 113050 165454
rect 113286 165218 143770 165454
rect 144006 165218 174490 165454
rect 174726 165218 205210 165454
rect 205446 165218 235930 165454
rect 236166 165218 266650 165454
rect 266886 165218 297370 165454
rect 297606 165218 328090 165454
rect 328326 165218 358810 165454
rect 359046 165218 389530 165454
rect 389766 165218 420250 165454
rect 420486 165218 450970 165454
rect 451206 165218 481690 165454
rect 481926 165218 512410 165454
rect 512646 165218 543130 165454
rect 543366 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 51610 165134
rect 51846 164898 82330 165134
rect 82566 164898 113050 165134
rect 113286 164898 143770 165134
rect 144006 164898 174490 165134
rect 174726 164898 205210 165134
rect 205446 164898 235930 165134
rect 236166 164898 266650 165134
rect 266886 164898 297370 165134
rect 297606 164898 328090 165134
rect 328326 164898 358810 165134
rect 359046 164898 389530 165134
rect 389766 164898 420250 165134
rect 420486 164898 450970 165134
rect 451206 164898 481690 165134
rect 481926 164898 512410 165134
rect 512646 164898 543130 165134
rect 543366 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 36250 147454
rect 36486 147218 66970 147454
rect 67206 147218 97690 147454
rect 97926 147218 128410 147454
rect 128646 147218 159130 147454
rect 159366 147218 189850 147454
rect 190086 147218 220570 147454
rect 220806 147218 251290 147454
rect 251526 147218 282010 147454
rect 282246 147218 312730 147454
rect 312966 147218 343450 147454
rect 343686 147218 374170 147454
rect 374406 147218 404890 147454
rect 405126 147218 435610 147454
rect 435846 147218 466330 147454
rect 466566 147218 497050 147454
rect 497286 147218 527770 147454
rect 528006 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 36250 147134
rect 36486 146898 66970 147134
rect 67206 146898 97690 147134
rect 97926 146898 128410 147134
rect 128646 146898 159130 147134
rect 159366 146898 189850 147134
rect 190086 146898 220570 147134
rect 220806 146898 251290 147134
rect 251526 146898 282010 147134
rect 282246 146898 312730 147134
rect 312966 146898 343450 147134
rect 343686 146898 374170 147134
rect 374406 146898 404890 147134
rect 405126 146898 435610 147134
rect 435846 146898 466330 147134
rect 466566 146898 497050 147134
rect 497286 146898 527770 147134
rect 528006 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 51610 129454
rect 51846 129218 82330 129454
rect 82566 129218 113050 129454
rect 113286 129218 143770 129454
rect 144006 129218 174490 129454
rect 174726 129218 205210 129454
rect 205446 129218 235930 129454
rect 236166 129218 266650 129454
rect 266886 129218 297370 129454
rect 297606 129218 328090 129454
rect 328326 129218 358810 129454
rect 359046 129218 389530 129454
rect 389766 129218 420250 129454
rect 420486 129218 450970 129454
rect 451206 129218 481690 129454
rect 481926 129218 512410 129454
rect 512646 129218 543130 129454
rect 543366 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 51610 129134
rect 51846 128898 82330 129134
rect 82566 128898 113050 129134
rect 113286 128898 143770 129134
rect 144006 128898 174490 129134
rect 174726 128898 205210 129134
rect 205446 128898 235930 129134
rect 236166 128898 266650 129134
rect 266886 128898 297370 129134
rect 297606 128898 328090 129134
rect 328326 128898 358810 129134
rect 359046 128898 389530 129134
rect 389766 128898 420250 129134
rect 420486 128898 450970 129134
rect 451206 128898 481690 129134
rect 481926 128898 512410 129134
rect 512646 128898 543130 129134
rect 543366 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 36250 111454
rect 36486 111218 66970 111454
rect 67206 111218 97690 111454
rect 97926 111218 128410 111454
rect 128646 111218 159130 111454
rect 159366 111218 189850 111454
rect 190086 111218 220570 111454
rect 220806 111218 251290 111454
rect 251526 111218 282010 111454
rect 282246 111218 312730 111454
rect 312966 111218 343450 111454
rect 343686 111218 374170 111454
rect 374406 111218 404890 111454
rect 405126 111218 435610 111454
rect 435846 111218 466330 111454
rect 466566 111218 497050 111454
rect 497286 111218 527770 111454
rect 528006 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 36250 111134
rect 36486 110898 66970 111134
rect 67206 110898 97690 111134
rect 97926 110898 128410 111134
rect 128646 110898 159130 111134
rect 159366 110898 189850 111134
rect 190086 110898 220570 111134
rect 220806 110898 251290 111134
rect 251526 110898 282010 111134
rect 282246 110898 312730 111134
rect 312966 110898 343450 111134
rect 343686 110898 374170 111134
rect 374406 110898 404890 111134
rect 405126 110898 435610 111134
rect 435846 110898 466330 111134
rect 466566 110898 497050 111134
rect 497286 110898 527770 111134
rect 528006 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 51610 93454
rect 51846 93218 82330 93454
rect 82566 93218 113050 93454
rect 113286 93218 143770 93454
rect 144006 93218 174490 93454
rect 174726 93218 205210 93454
rect 205446 93218 235930 93454
rect 236166 93218 266650 93454
rect 266886 93218 297370 93454
rect 297606 93218 328090 93454
rect 328326 93218 358810 93454
rect 359046 93218 389530 93454
rect 389766 93218 420250 93454
rect 420486 93218 450970 93454
rect 451206 93218 481690 93454
rect 481926 93218 512410 93454
rect 512646 93218 543130 93454
rect 543366 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 51610 93134
rect 51846 92898 82330 93134
rect 82566 92898 113050 93134
rect 113286 92898 143770 93134
rect 144006 92898 174490 93134
rect 174726 92898 205210 93134
rect 205446 92898 235930 93134
rect 236166 92898 266650 93134
rect 266886 92898 297370 93134
rect 297606 92898 328090 93134
rect 328326 92898 358810 93134
rect 359046 92898 389530 93134
rect 389766 92898 420250 93134
rect 420486 92898 450970 93134
rect 451206 92898 481690 93134
rect 481926 92898 512410 93134
rect 512646 92898 543130 93134
rect 543366 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 36250 75454
rect 36486 75218 66970 75454
rect 67206 75218 97690 75454
rect 97926 75218 128410 75454
rect 128646 75218 159130 75454
rect 159366 75218 189850 75454
rect 190086 75218 220570 75454
rect 220806 75218 251290 75454
rect 251526 75218 282010 75454
rect 282246 75218 312730 75454
rect 312966 75218 343450 75454
rect 343686 75218 374170 75454
rect 374406 75218 404890 75454
rect 405126 75218 435610 75454
rect 435846 75218 466330 75454
rect 466566 75218 497050 75454
rect 497286 75218 527770 75454
rect 528006 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 36250 75134
rect 36486 74898 66970 75134
rect 67206 74898 97690 75134
rect 97926 74898 128410 75134
rect 128646 74898 159130 75134
rect 159366 74898 189850 75134
rect 190086 74898 220570 75134
rect 220806 74898 251290 75134
rect 251526 74898 282010 75134
rect 282246 74898 312730 75134
rect 312966 74898 343450 75134
rect 343686 74898 374170 75134
rect 374406 74898 404890 75134
rect 405126 74898 435610 75134
rect 435846 74898 466330 75134
rect 466566 74898 497050 75134
rect 497286 74898 527770 75134
rect 528006 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 51610 57454
rect 51846 57218 82330 57454
rect 82566 57218 113050 57454
rect 113286 57218 143770 57454
rect 144006 57218 174490 57454
rect 174726 57218 205210 57454
rect 205446 57218 235930 57454
rect 236166 57218 266650 57454
rect 266886 57218 297370 57454
rect 297606 57218 328090 57454
rect 328326 57218 358810 57454
rect 359046 57218 389530 57454
rect 389766 57218 420250 57454
rect 420486 57218 450970 57454
rect 451206 57218 481690 57454
rect 481926 57218 512410 57454
rect 512646 57218 543130 57454
rect 543366 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 51610 57134
rect 51846 56898 82330 57134
rect 82566 56898 113050 57134
rect 113286 56898 143770 57134
rect 144006 56898 174490 57134
rect 174726 56898 205210 57134
rect 205446 56898 235930 57134
rect 236166 56898 266650 57134
rect 266886 56898 297370 57134
rect 297606 56898 328090 57134
rect 328326 56898 358810 57134
rect 359046 56898 389530 57134
rect 389766 56898 420250 57134
rect 420486 56898 450970 57134
rect 451206 56898 481690 57134
rect 481926 56898 512410 57134
rect 512646 56898 543130 57134
rect 543366 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 36250 39454
rect 36486 39218 66970 39454
rect 67206 39218 97690 39454
rect 97926 39218 128410 39454
rect 128646 39218 159130 39454
rect 159366 39218 189850 39454
rect 190086 39218 220570 39454
rect 220806 39218 251290 39454
rect 251526 39218 282010 39454
rect 282246 39218 312730 39454
rect 312966 39218 343450 39454
rect 343686 39218 374170 39454
rect 374406 39218 404890 39454
rect 405126 39218 435610 39454
rect 435846 39218 466330 39454
rect 466566 39218 497050 39454
rect 497286 39218 527770 39454
rect 528006 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 36250 39134
rect 36486 38898 66970 39134
rect 67206 38898 97690 39134
rect 97926 38898 128410 39134
rect 128646 38898 159130 39134
rect 159366 38898 189850 39134
rect 190086 38898 220570 39134
rect 220806 38898 251290 39134
rect 251526 38898 282010 39134
rect 282246 38898 312730 39134
rect 312966 38898 343450 39134
rect 343686 38898 374170 39134
rect 374406 38898 404890 39134
rect 405126 38898 435610 39134
rect 435846 38898 466330 39134
rect 466566 38898 497050 39134
rect 497286 38898 527770 39134
rect 528006 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1635763811
transform 1 0 32000 0 1 32000
box 474 0 519418 640000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 30000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 674000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 674000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 674000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 674000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 674000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 674000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 674000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 674000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 674000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 674000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 674000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 674000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 674000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 674000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 674000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 30000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 674000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 674000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 674000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 674000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 674000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 674000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 674000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 674000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 674000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 674000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 674000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 674000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 674000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 674000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 674000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 30000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 674000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 674000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 674000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 674000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 674000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 674000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 674000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 674000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 674000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 674000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 674000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 674000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 674000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 674000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 674000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 30000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 674000 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 674000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 674000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 674000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 674000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 674000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 674000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 674000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 674000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 674000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 674000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 674000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 674000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 674000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 674000 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 30000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 674000 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 674000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 674000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 674000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 674000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 674000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 674000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 674000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 674000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 674000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 674000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 674000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 674000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 674000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 30000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 674000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 674000 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 674000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 674000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 674000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 674000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 674000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 674000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 674000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 674000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 674000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 674000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 674000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 674000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 674000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 30000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 674000 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 674000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 674000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 674000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 674000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 674000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 674000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 674000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 674000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 674000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 674000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 674000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 674000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 674000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 30000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 674000 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 674000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 674000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 674000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 674000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 674000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 674000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 674000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 674000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 674000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 674000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 674000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 674000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 674000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
