magic
tech sky130A
magscale 1 2
timestamp 1635585791
<< locali >>
rect 307033 700111 307067 700485
rect 37289 697731 37323 699057
rect 42441 698411 42475 699057
rect 52377 697867 52411 699057
rect 67557 698003 67591 699057
rect 72801 698547 72835 699057
rect 82737 698139 82771 699057
rect 97917 698275 97951 699057
rect 103161 698751 103195 699057
rect 490941 698207 490975 698989
rect 495909 698683 495943 698989
rect 506029 698071 506063 698989
rect 511181 698615 511215 698989
rect 516149 698479 516183 698989
rect 521117 697935 521151 698989
rect 536389 697799 536423 698989
rect 546509 698343 546543 698989
rect 551477 697663 551511 698989
rect 566565 697595 566599 698989
rect 582389 33099 582423 702525
rect 582481 112863 582515 698377
rect 582573 126055 582607 697833
rect 582665 152711 582699 702321
rect 582757 165903 582791 697969
rect 582849 179231 582883 701097
rect 582941 192559 582975 698513
rect 583033 205751 583067 698105
rect 583125 232407 583159 701233
rect 583217 245599 583251 698241
rect 583309 272255 583343 698717
rect 583401 312103 583435 701641
rect 583493 325295 583527 701437
rect 583585 351951 583619 702661
rect 583677 418319 583711 701845
rect 583769 431647 583803 701709
rect 583861 537863 583895 703001
<< viali >>
rect 583861 703001 583895 703035
rect 583585 702661 583619 702695
rect 582389 702525 582423 702559
rect 307033 700485 307067 700519
rect 307033 700077 307067 700111
rect 37289 699057 37323 699091
rect 42441 699057 42475 699091
rect 42441 698377 42475 698411
rect 52377 699057 52411 699091
rect 67557 699057 67591 699091
rect 72801 699057 72835 699091
rect 72801 698513 72835 698547
rect 82737 699057 82771 699091
rect 97917 699057 97951 699091
rect 103161 699057 103195 699091
rect 103161 698717 103195 698751
rect 490941 698989 490975 699023
rect 97917 698241 97951 698275
rect 495909 698989 495943 699023
rect 495909 698649 495943 698683
rect 506029 698989 506063 699023
rect 490941 698173 490975 698207
rect 82737 698105 82771 698139
rect 511181 698989 511215 699023
rect 511181 698581 511215 698615
rect 516149 698989 516183 699023
rect 516149 698445 516183 698479
rect 521117 698989 521151 699023
rect 506029 698037 506063 698071
rect 67557 697969 67591 698003
rect 521117 697901 521151 697935
rect 536389 698989 536423 699023
rect 52377 697833 52411 697867
rect 546509 698989 546543 699023
rect 546509 698309 546543 698343
rect 551477 698989 551511 699023
rect 536389 697765 536423 697799
rect 37289 697697 37323 697731
rect 551477 697629 551511 697663
rect 566565 698989 566599 699023
rect 566565 697561 566599 697595
rect 582665 702321 582699 702355
rect 582481 698377 582515 698411
rect 582573 697833 582607 697867
rect 583401 701641 583435 701675
rect 583125 701233 583159 701267
rect 582849 701097 582883 701131
rect 582757 697969 582791 698003
rect 582941 698513 582975 698547
rect 583033 698105 583067 698139
rect 583309 698717 583343 698751
rect 583217 698241 583251 698275
rect 583493 701437 583527 701471
rect 583677 701845 583711 701879
rect 583769 701709 583803 701743
rect 583861 537829 583895 537863
rect 583769 431613 583803 431647
rect 583677 418285 583711 418319
rect 583585 351917 583619 351951
rect 583493 325261 583527 325295
rect 583401 312069 583435 312103
rect 583309 272221 583343 272255
rect 583217 245565 583251 245599
rect 583125 232373 583159 232407
rect 583033 205717 583067 205751
rect 582941 192525 582975 192559
rect 582849 179197 582883 179231
rect 582757 165869 582791 165903
rect 582665 152677 582699 152711
rect 582573 126021 582607 126055
rect 582481 112829 582515 112863
rect 582389 33065 582423 33099
<< metal1 >>
rect 6914 703808 6920 703860
rect 6972 703848 6978 703860
rect 581638 703848 581644 703860
rect 6972 703820 581644 703848
rect 6972 703808 6978 703820
rect 581638 703808 581644 703820
rect 581696 703808 581702 703860
rect 279326 703740 279332 703792
rect 279384 703780 279390 703792
rect 356054 703780 356060 703792
rect 279384 703752 356060 703780
rect 279384 703740 279390 703752
rect 356054 703740 356060 703752
rect 356112 703740 356118 703792
rect 238938 703672 238944 703724
rect 238996 703712 239002 703724
rect 316034 703712 316040 703724
rect 238996 703684 316040 703712
rect 238996 703672 239002 703684
rect 316034 703672 316040 703684
rect 316092 703672 316098 703724
rect 264146 703604 264152 703656
rect 264204 703644 264210 703656
rect 364242 703644 364248 703656
rect 264204 703616 364248 703644
rect 264204 703604 264210 703616
rect 364242 703604 364248 703616
rect 364300 703604 364306 703656
rect 249058 703536 249064 703588
rect 249116 703576 249122 703588
rect 410426 703576 410432 703588
rect 249116 703548 410432 703576
rect 249116 703536 249122 703548
rect 410426 703536 410432 703548
rect 410484 703536 410490 703588
rect 233878 703468 233884 703520
rect 233936 703508 233942 703520
rect 430022 703508 430028 703520
rect 233936 703480 430028 703508
rect 233936 703468 233942 703480
rect 430022 703468 430028 703480
rect 430080 703468 430086 703520
rect 218790 703400 218796 703452
rect 218848 703440 218854 703452
rect 581546 703440 581552 703452
rect 218848 703412 581552 703440
rect 218848 703400 218854 703412
rect 581546 703400 581552 703412
rect 581604 703400 581610 703452
rect 1486 703332 1492 703384
rect 1544 703372 1550 703384
rect 370130 703372 370136 703384
rect 1544 703344 370136 703372
rect 1544 703332 1550 703344
rect 370130 703332 370136 703344
rect 370188 703332 370194 703384
rect 203610 703264 203616 703316
rect 203668 703304 203674 703316
rect 582282 703304 582288 703316
rect 203668 703276 582288 703304
rect 203668 703264 203674 703276
rect 582282 703264 582288 703276
rect 582340 703264 582346 703316
rect 1670 703196 1676 703248
rect 1728 703236 1734 703248
rect 385310 703236 385316 703248
rect 1728 703208 385316 703236
rect 1728 703196 1734 703208
rect 385310 703196 385316 703208
rect 385368 703196 385374 703248
rect 188522 703128 188528 703180
rect 188580 703168 188586 703180
rect 582190 703168 582196 703180
rect 188580 703140 582196 703168
rect 188580 703128 188586 703140
rect 582190 703128 582196 703140
rect 582248 703128 582254 703180
rect 1762 703060 1768 703112
rect 1820 703100 1826 703112
rect 400398 703100 400404 703112
rect 1820 703072 400404 703100
rect 1820 703060 1826 703072
rect 400398 703060 400404 703072
rect 400456 703060 400462 703112
rect 178402 702992 178408 703044
rect 178460 703032 178466 703044
rect 583849 703035 583907 703041
rect 583849 703032 583861 703035
rect 178460 703004 583861 703032
rect 178460 702992 178466 703004
rect 583849 703001 583861 703004
rect 583895 703001 583907 703035
rect 583849 702995 583907 703001
rect 173342 702924 173348 702976
rect 173400 702964 173406 702976
rect 582098 702964 582104 702976
rect 173400 702936 582104 702964
rect 173400 702924 173406 702936
rect 582098 702924 582104 702936
rect 582156 702924 582162 702976
rect 1854 702856 1860 702908
rect 1912 702896 1918 702908
rect 415578 702896 415584 702908
rect 1912 702868 415584 702896
rect 1912 702856 1918 702868
rect 415578 702856 415584 702868
rect 415636 702856 415642 702908
rect 158254 702788 158260 702840
rect 158312 702828 158318 702840
rect 582006 702828 582012 702840
rect 158312 702800 582012 702828
rect 158312 702788 158318 702800
rect 582006 702788 582012 702800
rect 582064 702788 582070 702840
rect 2406 702720 2412 702772
rect 2464 702760 2470 702772
rect 445846 702760 445852 702772
rect 2464 702732 445852 702760
rect 2464 702720 2470 702732
rect 445846 702720 445852 702732
rect 445904 702720 445910 702772
rect 127986 702652 127992 702704
rect 128044 702692 128050 702704
rect 583573 702695 583631 702701
rect 583573 702692 583585 702695
rect 128044 702664 583585 702692
rect 128044 702652 128050 702664
rect 583573 702661 583585 702664
rect 583619 702661 583631 702695
rect 583573 702655 583631 702661
rect 22002 702584 22008 702636
rect 22060 702624 22066 702636
rect 581730 702624 581736 702636
rect 22060 702596 581736 702624
rect 22060 702584 22066 702596
rect 581730 702584 581736 702596
rect 581788 702584 581794 702636
rect 11882 702516 11888 702568
rect 11940 702556 11946 702568
rect 582377 702559 582435 702565
rect 582377 702556 582389 702559
rect 11940 702528 582389 702556
rect 11940 702516 11946 702528
rect 582377 702525 582389 702528
rect 582423 702525 582435 702559
rect 582377 702519 582435 702525
rect 270678 702448 270684 702500
rect 270736 702488 270742 702500
rect 314654 702488 314660 702500
rect 270736 702460 314660 702488
rect 270736 702448 270742 702460
rect 314654 702448 314660 702460
rect 314712 702448 314718 702500
rect 57330 702312 57336 702364
rect 57388 702352 57394 702364
rect 582653 702355 582711 702361
rect 582653 702352 582665 702355
rect 57388 702324 582665 702352
rect 57388 702312 57394 702324
rect 582653 702321 582665 702324
rect 582699 702321 582711 702355
rect 582653 702315 582711 702321
rect 243998 702244 244004 702296
rect 244056 702284 244062 702296
rect 320818 702284 320824 702296
rect 244056 702256 320824 702284
rect 244056 702244 244062 702256
rect 320818 702244 320824 702256
rect 320876 702244 320882 702296
rect 286962 702176 286968 702228
rect 287020 702216 287026 702228
rect 410518 702216 410524 702228
rect 287020 702188 410524 702216
rect 287020 702176 287026 702188
rect 410518 702176 410524 702188
rect 410576 702176 410582 702228
rect 168282 702108 168288 702160
rect 168340 702148 168346 702160
rect 336550 702148 336556 702160
rect 168340 702120 336556 702148
rect 168340 702108 168346 702120
rect 336550 702108 336556 702120
rect 336608 702108 336614 702160
rect 133046 702040 133052 702092
rect 133104 702080 133110 702092
rect 329834 702080 329840 702092
rect 133104 702052 329840 702080
rect 133104 702040 133110 702052
rect 329834 702040 329840 702052
rect 329892 702040 329898 702092
rect 332594 702040 332600 702092
rect 332652 702080 332658 702092
rect 380250 702080 380256 702092
rect 332652 702052 380256 702080
rect 332652 702040 332658 702052
rect 380250 702040 380256 702052
rect 380308 702040 380314 702092
rect 138014 701972 138020 702024
rect 138072 702012 138078 702024
rect 342070 702012 342076 702024
rect 138072 701984 342076 702012
rect 138072 701972 138078 701984
rect 342070 701972 342076 701984
rect 342128 701972 342134 702024
rect 266354 701904 266360 701956
rect 266412 701944 266418 701956
rect 481174 701944 481180 701956
rect 266412 701916 481180 701944
rect 266412 701904 266418 701916
rect 481174 701904 481180 701916
rect 481232 701904 481238 701956
rect 47210 701836 47216 701888
rect 47268 701876 47274 701888
rect 144362 701876 144368 701888
rect 47268 701848 144368 701876
rect 47268 701836 47274 701848
rect 144362 701836 144368 701848
rect 144420 701836 144426 701888
rect 153194 701836 153200 701888
rect 153252 701876 153258 701888
rect 583665 701879 583723 701885
rect 583665 701876 583677 701879
rect 153252 701848 583677 701876
rect 153252 701836 153258 701848
rect 583665 701845 583677 701848
rect 583711 701845 583723 701879
rect 583665 701839 583723 701845
rect 4706 701768 4712 701820
rect 4764 701808 4770 701820
rect 440786 701808 440792 701820
rect 4764 701780 440792 701808
rect 4764 701768 4770 701780
rect 440786 701768 440792 701780
rect 440844 701768 440850 701820
rect 32122 701700 32128 701752
rect 32180 701740 32186 701752
rect 132678 701740 132684 701752
rect 32180 701712 132684 701740
rect 32180 701700 32186 701712
rect 132678 701700 132684 701712
rect 132736 701700 132742 701752
rect 148134 701700 148140 701752
rect 148192 701740 148198 701752
rect 583757 701743 583815 701749
rect 583757 701740 583769 701743
rect 148192 701712 583769 701740
rect 148192 701700 148198 701712
rect 583757 701709 583769 701712
rect 583803 701709 583815 701743
rect 583757 701703 583815 701709
rect 122926 701632 122932 701684
rect 122984 701672 122990 701684
rect 583389 701675 583447 701681
rect 583389 701672 583401 701675
rect 122984 701644 583401 701672
rect 122984 701632 122990 701644
rect 583389 701641 583401 701644
rect 583435 701641 583447 701675
rect 583389 701635 583447 701641
rect 566 701564 572 701616
rect 624 701604 630 701616
rect 465994 701604 466000 701616
rect 624 701576 466000 701604
rect 624 701564 630 701576
rect 465994 701564 466000 701576
rect 466052 701564 466058 701616
rect 4890 701496 4896 701548
rect 4948 701536 4954 701548
rect 471054 701536 471060 701548
rect 4948 701508 471060 701536
rect 4948 701496 4954 701508
rect 471054 701496 471060 701508
rect 471112 701496 471118 701548
rect 117866 701428 117872 701480
rect 117924 701468 117930 701480
rect 583481 701471 583539 701477
rect 583481 701468 583493 701471
rect 117924 701440 583493 701468
rect 117924 701428 117930 701440
rect 583481 701437 583493 701440
rect 583527 701437 583539 701471
rect 583481 701431 583539 701437
rect 4798 701360 4804 701412
rect 4856 701400 4862 701412
rect 486234 701400 486240 701412
rect 4856 701372 486240 701400
rect 4856 701360 4862 701372
rect 486234 701360 486240 701372
rect 486292 701360 486298 701412
rect 92658 701292 92664 701344
rect 92716 701332 92722 701344
rect 581914 701332 581920 701344
rect 92716 701304 581920 701332
rect 92716 701292 92722 701304
rect 581914 701292 581920 701304
rect 581972 701292 581978 701344
rect 87598 701224 87604 701276
rect 87656 701264 87662 701276
rect 583113 701267 583171 701273
rect 583113 701264 583125 701267
rect 87656 701236 583125 701264
rect 87656 701224 87662 701236
rect 583113 701233 583125 701236
rect 583159 701233 583171 701267
rect 583113 701227 583171 701233
rect 4614 701156 4620 701208
rect 4672 701196 4678 701208
rect 501322 701196 501328 701208
rect 4672 701168 501328 701196
rect 4672 701156 4678 701168
rect 501322 701156 501328 701168
rect 501380 701156 501386 701208
rect 571978 701156 571984 701208
rect 572036 701196 572042 701208
rect 582558 701196 582564 701208
rect 572036 701168 582564 701196
rect 572036 701156 572042 701168
rect 582558 701156 582564 701168
rect 582616 701156 582622 701208
rect 77478 701088 77484 701140
rect 77536 701128 77542 701140
rect 582837 701131 582895 701137
rect 582837 701128 582849 701131
rect 77536 701100 582849 701128
rect 77536 701088 77542 701100
rect 582837 701097 582849 701100
rect 582883 701097 582895 701131
rect 582837 701091 582895 701097
rect 259178 701020 259184 701072
rect 259236 701060 259242 701072
rect 303522 701060 303528 701072
rect 259236 701032 303528 701060
rect 259236 701020 259242 701032
rect 303522 701020 303528 701032
rect 303580 701020 303586 701072
rect 554774 701020 554780 701072
rect 554832 701060 554838 701072
rect 577038 701060 577044 701072
rect 554832 701032 577044 701060
rect 554832 701020 554838 701032
rect 577038 701020 577044 701032
rect 577096 701020 577102 701072
rect 218974 700952 218980 701004
rect 219032 700992 219038 701004
rect 319714 700992 319720 701004
rect 219032 700964 319720 700992
rect 219032 700952 219038 700964
rect 319714 700952 319720 700964
rect 319772 700952 319778 701004
rect 356054 700952 356060 701004
rect 356112 700992 356118 701004
rect 364978 700992 364984 701004
rect 356112 700964 364984 700992
rect 356112 700952 356118 700964
rect 364978 700952 364984 700964
rect 365036 700952 365042 701004
rect 235166 700884 235172 700936
rect 235224 700924 235230 700936
rect 309594 700924 309600 700936
rect 235224 700896 309600 700924
rect 235224 700884 235230 700896
rect 309594 700884 309600 700896
rect 309652 700884 309658 700936
rect 316034 700884 316040 700936
rect 316092 700924 316098 700936
rect 527174 700924 527180 700936
rect 316092 700896 527180 700924
rect 316092 700884 316098 700896
rect 527174 700884 527180 700896
rect 527232 700884 527238 700936
rect 3786 700816 3792 700868
rect 3844 700856 3850 700868
rect 218054 700856 218060 700868
rect 3844 700828 218060 700856
rect 3844 700816 3850 700828
rect 218054 700816 218060 700828
rect 218112 700816 218118 700868
rect 254118 700816 254124 700868
rect 254176 700856 254182 700868
rect 462314 700856 462320 700868
rect 254176 700828 462320 700856
rect 254176 700816 254182 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 105446 700748 105452 700800
rect 105504 700788 105510 700800
rect 339862 700788 339868 700800
rect 105504 700760 339868 700788
rect 105504 700748 105510 700760
rect 339862 700748 339868 700760
rect 339920 700748 339926 700800
rect 342070 700748 342076 700800
rect 342128 700788 342134 700800
rect 580534 700788 580540 700800
rect 342128 700760 580540 700788
rect 342128 700748 342134 700760
rect 580534 700748 580540 700760
rect 580592 700748 580598 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 349982 700720 349988 700732
rect 89220 700692 349988 700720
rect 89220 700680 89226 700692
rect 349982 700680 349988 700692
rect 350040 700680 350046 700732
rect 364242 700680 364248 700732
rect 364300 700720 364306 700732
rect 429838 700720 429844 700732
rect 364300 700692 429844 700720
rect 364300 700680 364306 700692
rect 429838 700680 429844 700692
rect 429896 700680 429902 700732
rect 430022 700680 430028 700732
rect 430080 700720 430086 700732
rect 559650 700720 559656 700732
rect 430080 700692 559656 700720
rect 430080 700680 430086 700692
rect 559650 700680 559656 700692
rect 559708 700680 559714 700732
rect 4062 700612 4068 700664
rect 4120 700652 4126 700664
rect 266354 700652 266360 700664
rect 4120 700624 266360 700652
rect 4120 700612 4126 700624
rect 266354 700612 266360 700624
rect 266412 700612 266418 700664
rect 284386 700612 284392 700664
rect 284444 700652 284450 700664
rect 332502 700652 332508 700664
rect 284444 700624 332508 700652
rect 284444 700612 284450 700624
rect 332502 700612 332508 700624
rect 332560 700612 332566 700664
rect 336550 700612 336556 700664
rect 336608 700652 336614 700664
rect 580810 700652 580816 700664
rect 336608 700624 580816 700652
rect 336608 700612 336614 700624
rect 580810 700612 580816 700624
rect 580868 700612 580874 700664
rect 72970 700544 72976 700596
rect 73028 700584 73034 700596
rect 344922 700584 344928 700596
rect 73028 700556 344928 700584
rect 73028 700544 73034 700556
rect 344922 700544 344928 700556
rect 344980 700544 344986 700596
rect 410426 700544 410432 700596
rect 410484 700584 410490 700596
rect 494790 700584 494796 700596
rect 410484 700556 494796 700584
rect 410484 700544 410490 700556
rect 494790 700544 494796 700556
rect 494848 700544 494854 700596
rect 3234 700476 3240 700528
rect 3292 700516 3298 700528
rect 286962 700516 286968 700528
rect 3292 700488 286968 700516
rect 3292 700476 3298 700488
rect 286962 700476 286968 700488
rect 287020 700476 287026 700528
rect 294506 700476 294512 700528
rect 294564 700516 294570 700528
rect 300118 700516 300124 700528
rect 294564 700488 300124 700516
rect 294564 700476 294570 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 303522 700476 303528 700528
rect 303580 700516 303586 700528
rect 307021 700519 307079 700525
rect 307021 700516 307033 700519
rect 303580 700488 307033 700516
rect 303580 700476 303586 700488
rect 307021 700485 307033 700488
rect 307067 700485 307079 700519
rect 307021 700479 307079 700485
rect 329834 700476 329840 700528
rect 329892 700516 329898 700528
rect 580718 700516 580724 700528
rect 329892 700488 580724 700516
rect 329892 700476 329898 700488
rect 580718 700476 580724 700488
rect 580776 700476 580782 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 355042 700448 355048 700460
rect 40552 700420 355048 700448
rect 40552 700408 40558 700420
rect 355042 700408 355048 700420
rect 355100 700408 355106 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 365070 700380 365076 700392
rect 24360 700352 365076 700380
rect 24360 700340 24366 700352
rect 365070 700340 365076 700352
rect 365128 700340 365134 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 360010 700312 360016 700324
rect 8168 700284 360016 700312
rect 8168 700272 8174 700284
rect 360010 700272 360016 700284
rect 360068 700272 360074 700324
rect 137830 700204 137836 700256
rect 137888 700244 137894 700256
rect 329742 700244 329748 700256
rect 137888 700216 329748 700244
rect 137888 700204 137894 700216
rect 329742 700204 329748 700216
rect 329800 700204 329806 700256
rect 154114 700136 154120 700188
rect 154172 700176 154178 700188
rect 334802 700176 334808 700188
rect 154172 700148 334808 700176
rect 154172 700136 154178 700148
rect 334802 700136 334808 700148
rect 334860 700136 334866 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 270678 700108 270684 700120
rect 202840 700080 270684 700108
rect 202840 700068 202846 700080
rect 270678 700068 270684 700080
rect 270736 700068 270742 700120
rect 283834 700068 283840 700120
rect 283892 700108 283898 700120
rect 304534 700108 304540 700120
rect 283892 700080 304540 700108
rect 283892 700068 283898 700080
rect 304534 700068 304540 700080
rect 304592 700068 304598 700120
rect 307021 700111 307079 700117
rect 307021 700077 307033 700111
rect 307067 700108 307079 700111
rect 478506 700108 478512 700120
rect 307067 700080 478512 700108
rect 307067 700077 307079 700080
rect 307021 700071 307079 700077
rect 478506 700068 478512 700080
rect 478564 700068 478570 700120
rect 170306 700000 170312 700052
rect 170364 700040 170370 700052
rect 324774 700040 324780 700052
rect 170364 700012 324780 700040
rect 170364 700000 170370 700012
rect 324774 700000 324780 700012
rect 324832 700000 324838 700052
rect 274266 699932 274272 699984
rect 274324 699972 274330 699984
rect 413646 699972 413652 699984
rect 274324 699944 413652 699972
rect 274324 699932 274330 699944
rect 413646 699932 413652 699944
rect 413704 699932 413710 699984
rect 269206 699864 269212 699916
rect 269264 699904 269270 699916
rect 397454 699904 397460 699916
rect 269264 699876 397460 699904
rect 269264 699864 269270 699876
rect 397454 699864 397460 699876
rect 397512 699864 397518 699916
rect 289446 699796 289452 699848
rect 289504 699836 289510 699848
rect 348786 699836 348792 699848
rect 289504 699808 348792 699836
rect 289504 699796 289510 699808
rect 348786 699796 348792 699808
rect 348844 699796 348850 699848
rect 267642 699728 267648 699780
rect 267700 699768 267706 699780
rect 299474 699768 299480 699780
rect 267700 699740 299480 699768
rect 267700 699728 267706 699740
rect 299474 699728 299480 699740
rect 299532 699728 299538 699780
rect 320818 699728 320824 699780
rect 320876 699768 320882 699780
rect 543458 699768 543464 699780
rect 320876 699740 543464 699768
rect 320876 699728 320882 699740
rect 543458 699728 543464 699740
rect 543516 699728 543522 699780
rect 658 699660 664 699712
rect 716 699700 722 699712
rect 435726 699700 435732 699712
rect 716 699672 435732 699700
rect 716 699660 722 699672
rect 435726 699660 435732 699672
rect 435784 699660 435790 699712
rect 3694 699592 3700 699644
rect 3752 699632 3758 699644
rect 332594 699632 332600 699644
rect 3752 699604 332600 699632
rect 3752 699592 3758 699604
rect 332594 699592 332600 699604
rect 332652 699592 332658 699644
rect 229002 699524 229008 699576
rect 229060 699564 229066 699576
rect 579982 699564 579988 699576
rect 229060 699536 579988 699564
rect 229060 699524 229066 699536
rect 579982 699524 579988 699536
rect 580040 699524 580046 699576
rect 213822 699456 213828 699508
rect 213880 699496 213886 699508
rect 580074 699496 580080 699508
rect 213880 699468 580080 699496
rect 213880 699456 213886 699468
rect 580074 699456 580080 699468
rect 580132 699456 580138 699508
rect 144362 699388 144368 699440
rect 144420 699428 144426 699440
rect 580350 699428 580356 699440
rect 144420 699400 580356 699428
rect 144420 699388 144426 699400
rect 580350 699388 580356 699400
rect 580408 699388 580414 699440
rect 208946 699320 208952 699372
rect 209004 699360 209010 699372
rect 579062 699360 579068 699372
rect 209004 699332 579068 699360
rect 209004 699320 209010 699332
rect 579062 699320 579068 699332
rect 579120 699320 579126 699372
rect 1578 699252 1584 699304
rect 1636 699292 1642 699304
rect 374822 699292 374828 699304
rect 1636 699264 374828 699292
rect 1636 699252 1642 699264
rect 374822 699252 374828 699264
rect 374880 699252 374886 699304
rect 198734 699184 198740 699236
rect 198792 699224 198798 699236
rect 580166 699224 580172 699236
rect 198792 699196 580172 699224
rect 198792 699184 198798 699196
rect 580166 699184 580172 699196
rect 580224 699184 580230 699236
rect 3050 699116 3056 699168
rect 3108 699156 3114 699168
rect 395062 699156 395068 699168
rect 3108 699128 395068 699156
rect 3108 699116 3114 699128
rect 395062 699116 395068 699128
rect 395120 699116 395126 699168
rect 37274 699088 37280 699100
rect 37235 699060 37280 699088
rect 37274 699048 37280 699060
rect 37332 699048 37338 699100
rect 42426 699088 42432 699100
rect 42387 699060 42432 699088
rect 42426 699048 42432 699060
rect 42484 699048 42490 699100
rect 52362 699088 52368 699100
rect 52323 699060 52368 699088
rect 52362 699048 52368 699060
rect 52420 699048 52426 699100
rect 67542 699088 67548 699100
rect 67503 699060 67548 699088
rect 67542 699048 67548 699060
rect 67600 699048 67606 699100
rect 72786 699088 72792 699100
rect 72747 699060 72792 699088
rect 72786 699048 72792 699060
rect 72844 699048 72850 699100
rect 82722 699088 82728 699100
rect 82683 699060 82728 699088
rect 82722 699048 82728 699060
rect 82780 699048 82786 699100
rect 97902 699088 97908 699100
rect 97863 699060 97908 699088
rect 97902 699048 97908 699060
rect 97960 699048 97966 699100
rect 103146 699088 103152 699100
rect 103107 699060 103152 699088
rect 103146 699048 103152 699060
rect 103204 699048 103210 699100
rect 183554 699048 183560 699100
rect 183612 699088 183618 699100
rect 580902 699088 580908 699100
rect 183612 699060 580908 699088
rect 183612 699048 183618 699060
rect 580902 699048 580908 699060
rect 580960 699048 580966 699100
rect 750 698980 756 699032
rect 808 699020 814 699032
rect 405182 699020 405188 699032
rect 808 698992 405188 699020
rect 808 698980 814 698992
rect 405182 698980 405188 698992
rect 405240 698980 405246 699032
rect 420270 699020 420276 699032
rect 412606 698992 420276 699020
rect 2590 698912 2596 698964
rect 2648 698952 2654 698964
rect 412606 698952 412634 698992
rect 420270 698980 420276 698992
rect 420328 698980 420334 699032
rect 425238 699020 425244 699032
rect 422266 698992 425244 699020
rect 2648 698924 412634 698952
rect 2648 698912 2654 698924
rect 3142 698844 3148 698896
rect 3200 698884 3206 698896
rect 422266 698884 422294 698992
rect 425238 698980 425244 698992
rect 425296 698980 425302 699032
rect 455598 699020 455604 699032
rect 451246 698992 455604 699020
rect 3200 698856 422294 698884
rect 3200 698844 3206 698856
rect 3326 698776 3332 698828
rect 3384 698816 3390 698828
rect 451246 698816 451274 698992
rect 455598 698980 455604 698992
rect 455656 698980 455662 699032
rect 490926 699020 490932 699032
rect 490887 698992 490932 699020
rect 490926 698980 490932 698992
rect 490984 698980 490990 699032
rect 495894 699020 495900 699032
rect 495855 698992 495900 699020
rect 495894 698980 495900 698992
rect 495952 698980 495958 699032
rect 506014 699020 506020 699032
rect 505975 698992 506020 699020
rect 506014 698980 506020 698992
rect 506072 698980 506078 699032
rect 511166 699020 511172 699032
rect 511127 698992 511172 699020
rect 511166 698980 511172 698992
rect 511224 698980 511230 699032
rect 516134 699020 516140 699032
rect 516095 698992 516140 699020
rect 516134 698980 516140 698992
rect 516192 698980 516198 699032
rect 521102 699020 521108 699032
rect 521063 698992 521108 699020
rect 521102 698980 521108 698992
rect 521160 698980 521166 699032
rect 536374 699020 536380 699032
rect 536335 698992 536380 699020
rect 536374 698980 536380 698992
rect 536432 698980 536438 699032
rect 546494 699020 546500 699032
rect 546455 698992 546500 699020
rect 546494 698980 546500 698992
rect 546552 698980 546558 699032
rect 551462 699020 551468 699032
rect 551423 698992 551468 699020
rect 551462 698980 551468 698992
rect 551520 698980 551526 699032
rect 566550 699020 566556 699032
rect 566511 698992 566556 699020
rect 566550 698980 566556 698992
rect 566608 698980 566614 699032
rect 3384 698788 451274 698816
rect 3384 698776 3390 698788
rect 103149 698751 103207 698757
rect 103149 698717 103161 698751
rect 103195 698748 103207 698751
rect 583297 698751 583355 698757
rect 583297 698748 583309 698751
rect 103195 698720 583309 698748
rect 103195 698717 103207 698720
rect 103149 698711 103207 698717
rect 583297 698717 583309 698720
rect 583343 698717 583355 698751
rect 583297 698711 583355 698717
rect 2222 698640 2228 698692
rect 2280 698680 2286 698692
rect 495897 698683 495955 698689
rect 495897 698680 495909 698683
rect 2280 698652 495909 698680
rect 2280 698640 2286 698652
rect 495897 698649 495909 698652
rect 495943 698649 495955 698683
rect 495897 698643 495955 698649
rect 3878 698572 3884 698624
rect 3936 698612 3942 698624
rect 511169 698615 511227 698621
rect 511169 698612 511181 698615
rect 3936 698584 511181 698612
rect 3936 698572 3942 698584
rect 511169 698581 511181 698584
rect 511215 698581 511227 698615
rect 511169 698575 511227 698581
rect 72789 698547 72847 698553
rect 72789 698513 72801 698547
rect 72835 698544 72847 698547
rect 582929 698547 582987 698553
rect 582929 698544 582941 698547
rect 72835 698516 582941 698544
rect 72835 698513 72847 698516
rect 72789 698507 72847 698513
rect 582929 698513 582941 698516
rect 582975 698513 582987 698547
rect 582929 698507 582987 698513
rect 3970 698436 3976 698488
rect 4028 698476 4034 698488
rect 516137 698479 516195 698485
rect 516137 698476 516149 698479
rect 4028 698448 516149 698476
rect 4028 698436 4034 698448
rect 516137 698445 516149 698448
rect 516183 698445 516195 698479
rect 516137 698439 516195 698445
rect 42429 698411 42487 698417
rect 42429 698377 42441 698411
rect 42475 698408 42487 698411
rect 582469 698411 582527 698417
rect 582469 698408 582481 698411
rect 42475 698380 582481 698408
rect 42475 698377 42487 698380
rect 42429 698371 42487 698377
rect 582469 698377 582481 698380
rect 582515 698377 582527 698411
rect 582469 698371 582527 698377
rect 3602 698300 3608 698352
rect 3660 698340 3666 698352
rect 546497 698343 546555 698349
rect 546497 698340 546509 698343
rect 3660 698312 546509 698340
rect 3660 698300 3666 698312
rect 546497 698309 546509 698312
rect 546543 698309 546555 698343
rect 546497 698303 546555 698309
rect 97905 698275 97963 698281
rect 97905 698241 97917 698275
rect 97951 698272 97963 698275
rect 583205 698275 583263 698281
rect 583205 698272 583217 698275
rect 97951 698244 583217 698272
rect 97951 698241 97963 698244
rect 97905 698235 97963 698241
rect 583205 698241 583217 698244
rect 583251 698241 583263 698275
rect 583205 698235 583263 698241
rect 474 698164 480 698216
rect 532 698204 538 698216
rect 490929 698207 490987 698213
rect 490929 698204 490941 698207
rect 532 698176 490941 698204
rect 532 698164 538 698176
rect 490929 698173 490941 698176
rect 490975 698173 490987 698207
rect 490929 698167 490987 698173
rect 82725 698139 82783 698145
rect 82725 698105 82737 698139
rect 82771 698136 82783 698139
rect 583021 698139 583079 698145
rect 583021 698136 583033 698139
rect 82771 698108 583033 698136
rect 82771 698105 82783 698108
rect 82725 698099 82783 698105
rect 583021 698105 583033 698108
rect 583067 698105 583079 698139
rect 583021 698099 583079 698105
rect 382 698028 388 698080
rect 440 698068 446 698080
rect 506017 698071 506075 698077
rect 506017 698068 506029 698071
rect 440 698040 506029 698068
rect 440 698028 446 698040
rect 506017 698037 506029 698040
rect 506063 698037 506075 698071
rect 506017 698031 506075 698037
rect 67545 698003 67603 698009
rect 67545 697969 67557 698003
rect 67591 698000 67603 698003
rect 582745 698003 582803 698009
rect 582745 698000 582757 698003
rect 67591 697972 582757 698000
rect 67591 697969 67603 697972
rect 67545 697963 67603 697969
rect 582745 697969 582757 697972
rect 582791 697969 582803 698003
rect 582745 697963 582803 697969
rect 2130 697892 2136 697944
rect 2188 697932 2194 697944
rect 521105 697935 521163 697941
rect 521105 697932 521117 697935
rect 2188 697904 521117 697932
rect 2188 697892 2194 697904
rect 521105 697901 521117 697904
rect 521151 697901 521163 697935
rect 521105 697895 521163 697901
rect 52365 697867 52423 697873
rect 52365 697833 52377 697867
rect 52411 697864 52423 697867
rect 582561 697867 582619 697873
rect 582561 697864 582573 697867
rect 52411 697836 582573 697864
rect 52411 697833 52423 697836
rect 52365 697827 52423 697833
rect 582561 697833 582573 697836
rect 582607 697833 582619 697867
rect 582561 697827 582619 697833
rect 198 697756 204 697808
rect 256 697796 262 697808
rect 536377 697799 536435 697805
rect 536377 697796 536389 697799
rect 256 697768 536389 697796
rect 256 697756 262 697768
rect 536377 697765 536389 697768
rect 536423 697765 536435 697799
rect 536377 697759 536435 697765
rect 37277 697731 37335 697737
rect 37277 697697 37289 697731
rect 37323 697728 37335 697731
rect 581822 697728 581828 697740
rect 37323 697700 581828 697728
rect 37323 697697 37335 697700
rect 37277 697691 37335 697697
rect 581822 697688 581828 697700
rect 581880 697688 581886 697740
rect 106 697620 112 697672
rect 164 697660 170 697672
rect 551465 697663 551523 697669
rect 551465 697660 551477 697663
rect 164 697632 551477 697660
rect 164 697620 170 697632
rect 551465 697629 551477 697632
rect 551511 697629 551523 697663
rect 551465 697623 551523 697629
rect 14 697552 20 697604
rect 72 697592 78 697604
rect 566553 697595 566611 697601
rect 566553 697592 566565 697595
rect 72 697564 566565 697592
rect 72 697552 78 697564
rect 566553 697561 566565 697564
rect 566599 697561 566611 697595
rect 566553 697555 566611 697561
rect 3694 619556 3700 619608
rect 3752 619596 3758 619608
rect 4522 619596 4528 619608
rect 3752 619568 4528 619596
rect 3752 619556 3758 619568
rect 4522 619556 4528 619568
rect 4580 619556 4586 619608
rect 583386 537820 583392 537872
rect 583444 537860 583450 537872
rect 583849 537863 583907 537869
rect 583849 537860 583861 537863
rect 583444 537832 583861 537860
rect 583444 537820 583450 537832
rect 583849 537829 583861 537832
rect 583895 537829 583907 537863
rect 583849 537823 583907 537829
rect 3234 516128 3240 516180
rect 3292 516168 3298 516180
rect 4614 516168 4620 516180
rect 3292 516140 4620 516168
rect 3292 516128 3298 516140
rect 4614 516128 4620 516140
rect 4672 516128 4678 516180
rect 2774 462748 2780 462800
rect 2832 462788 2838 462800
rect 4706 462788 4712 462800
rect 2832 462760 4712 462788
rect 2832 462748 2838 462760
rect 4706 462748 4712 462760
rect 4764 462748 4770 462800
rect 583386 431604 583392 431656
rect 583444 431644 583450 431656
rect 583757 431647 583815 431653
rect 583757 431644 583769 431647
rect 583444 431616 583769 431644
rect 583444 431604 583450 431616
rect 583757 431613 583769 431616
rect 583803 431613 583815 431647
rect 583757 431607 583815 431613
rect 583386 418276 583392 418328
rect 583444 418316 583450 418328
rect 583665 418319 583723 418325
rect 583665 418316 583677 418319
rect 583444 418288 583677 418316
rect 583444 418276 583450 418288
rect 583665 418285 583677 418288
rect 583711 418285 583723 418319
rect 583665 418279 583723 418285
rect 583386 351908 583392 351960
rect 583444 351948 583450 351960
rect 583573 351951 583631 351957
rect 583573 351948 583585 351951
rect 583444 351920 583585 351948
rect 583444 351908 583450 351920
rect 583573 351917 583585 351920
rect 583619 351917 583631 351951
rect 583573 351911 583631 351917
rect 583386 325252 583392 325304
rect 583444 325292 583450 325304
rect 583481 325295 583539 325301
rect 583481 325292 583493 325295
rect 583444 325264 583493 325292
rect 583444 325252 583450 325264
rect 583481 325261 583493 325264
rect 583527 325261 583539 325295
rect 583481 325255 583539 325261
rect 583386 312100 583392 312112
rect 583347 312072 583392 312100
rect 583386 312060 583392 312072
rect 583444 312060 583450 312112
rect 2774 306212 2780 306264
rect 2832 306252 2838 306264
rect 4798 306252 4804 306264
rect 2832 306224 4804 306252
rect 2832 306212 2838 306224
rect 4798 306212 4804 306224
rect 4856 306212 4862 306264
rect 583294 272252 583300 272264
rect 583255 272224 583300 272252
rect 583294 272212 583300 272224
rect 583352 272212 583358 272264
rect 583202 245596 583208 245608
rect 583163 245568 583208 245596
rect 583202 245556 583208 245568
rect 583260 245556 583266 245608
rect 583110 232404 583116 232416
rect 583071 232376 583116 232404
rect 583110 232364 583116 232376
rect 583168 232364 583174 232416
rect 583018 205748 583024 205760
rect 582979 205720 583024 205748
rect 583018 205708 583024 205720
rect 583076 205708 583082 205760
rect 582926 192556 582932 192568
rect 582887 192528 582932 192556
rect 582926 192516 582932 192528
rect 582984 192516 582990 192568
rect 582834 179228 582840 179240
rect 582795 179200 582840 179228
rect 582834 179188 582840 179200
rect 582892 179188 582898 179240
rect 582742 165900 582748 165912
rect 582703 165872 582748 165900
rect 582742 165860 582748 165872
rect 582800 165860 582806 165912
rect 582650 152708 582656 152720
rect 582611 152680 582656 152708
rect 582650 152668 582656 152680
rect 582708 152668 582714 152720
rect 582561 126055 582619 126061
rect 582561 126021 582573 126055
rect 582607 126052 582619 126055
rect 582650 126052 582656 126064
rect 582607 126024 582656 126052
rect 582607 126021 582619 126024
rect 582561 126015 582619 126021
rect 582650 126012 582656 126024
rect 582708 126012 582714 126064
rect 582469 112863 582527 112869
rect 582469 112829 582481 112863
rect 582515 112860 582527 112863
rect 582650 112860 582656 112872
rect 582515 112832 582656 112860
rect 582515 112829 582527 112832
rect 582469 112823 582527 112829
rect 582650 112820 582656 112832
rect 582708 112820 582714 112872
rect 582377 33099 582435 33105
rect 582377 33065 582389 33099
rect 582423 33096 582435 33099
rect 582466 33096 582472 33108
rect 582423 33068 582472 33096
rect 582423 33065 582435 33068
rect 582377 33059 582435 33065
rect 582466 33056 582472 33068
rect 582524 33056 582530 33108
rect 3418 4088 3424 4140
rect 3476 4128 3482 4140
rect 582558 4128 582564 4140
rect 3476 4100 582564 4128
rect 3476 4088 3482 4100
rect 582558 4088 582564 4100
rect 582616 4088 582622 4140
rect 153010 4020 153016 4072
rect 153068 4060 153074 4072
rect 155402 4060 155408 4072
rect 153068 4032 155408 4060
rect 153068 4020 153074 4032
rect 155402 4020 155408 4032
rect 155460 4020 155466 4072
rect 155402 3884 155408 3936
rect 155460 3924 155466 3936
rect 157794 3924 157800 3936
rect 155460 3896 157800 3924
rect 155460 3884 155466 3896
rect 157794 3884 157800 3896
rect 157852 3884 157858 3936
rect 157794 3748 157800 3800
rect 157852 3788 157858 3800
rect 160094 3788 160100 3800
rect 157852 3760 160100 3788
rect 157852 3748 157858 3760
rect 160094 3748 160100 3760
rect 160152 3748 160158 3800
rect 66714 3680 66720 3732
rect 66772 3720 66778 3732
rect 70302 3720 70308 3732
rect 66772 3692 70308 3720
rect 66772 3680 66778 3692
rect 70302 3680 70308 3692
rect 70360 3680 70366 3732
rect 160094 3612 160100 3664
rect 160152 3652 160158 3664
rect 162486 3652 162492 3664
rect 160152 3624 162492 3652
rect 160152 3612 160158 3624
rect 162486 3612 162492 3624
rect 162544 3612 162550 3664
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 10778 3584 10784 3596
rect 6512 3556 10784 3584
rect 6512 3544 6518 3556
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 34790 3544 34796 3596
rect 34848 3584 34854 3596
rect 38746 3584 38752 3596
rect 34848 3556 38752 3584
rect 34848 3544 34854 3556
rect 38746 3544 38752 3556
rect 38804 3544 38810 3596
rect 54938 3544 54944 3596
rect 54996 3584 55002 3596
rect 58618 3584 58624 3596
rect 54996 3556 58624 3584
rect 54996 3544 55002 3556
rect 58618 3544 58624 3556
rect 58676 3544 58682 3596
rect 70302 3544 70308 3596
rect 70360 3584 70366 3596
rect 73798 3584 73804 3596
rect 70360 3556 73804 3584
rect 70360 3544 70366 3556
rect 73798 3544 73804 3556
rect 73856 3544 73862 3596
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 29454 3516 29460 3528
rect 25372 3488 29460 3516
rect 25372 3476 25378 3488
rect 29454 3476 29460 3488
rect 29512 3476 29518 3528
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 20070 3448 20076 3460
rect 15988 3420 20076 3448
rect 15988 3408 15994 3420
rect 20070 3408 20076 3420
rect 20128 3408 20134 3460
rect 45462 3408 45468 3460
rect 45520 3448 45526 3460
rect 49234 3448 49240 3460
rect 45520 3420 49240 3448
rect 45520 3408 45526 3420
rect 49234 3408 49240 3420
rect 49292 3408 49298 3460
rect 64322 3408 64328 3460
rect 64380 3448 64386 3460
rect 67910 3448 67916 3460
rect 64380 3420 67916 3448
rect 64380 3408 64386 3420
rect 67910 3408 67916 3420
rect 67968 3408 67974 3460
rect 73798 3408 73804 3460
rect 73856 3448 73862 3460
rect 77294 3448 77300 3460
rect 73856 3420 77300 3448
rect 73856 3408 73862 3420
rect 77294 3408 77300 3420
rect 77352 3408 77358 3460
rect 103330 3408 103336 3460
rect 103388 3448 103394 3460
rect 106458 3448 106464 3460
rect 103388 3420 106464 3448
rect 103388 3408 103394 3420
rect 106458 3408 106464 3420
rect 106516 3408 106522 3460
rect 46658 3136 46664 3188
rect 46716 3176 46722 3188
rect 50430 3176 50436 3188
rect 46716 3148 50436 3176
rect 46716 3136 46722 3148
rect 50430 3136 50436 3148
rect 50488 3136 50494 3188
rect 65518 3136 65524 3188
rect 65576 3176 65582 3188
rect 69106 3176 69112 3188
rect 65576 3148 69112 3176
rect 65576 3136 65582 3148
rect 69106 3136 69112 3148
rect 69164 3136 69170 3188
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 15470 3108 15476 3120
rect 11204 3080 15476 3108
rect 11204 3068 11210 3080
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 21266 3108 21272 3120
rect 17092 3080 21272 3108
rect 17092 3068 17098 3080
rect 21266 3068 21272 3080
rect 21324 3068 21330 3120
rect 28902 3068 28908 3120
rect 28960 3108 28966 3120
rect 32950 3108 32956 3120
rect 28960 3080 32956 3108
rect 28960 3068 28966 3080
rect 32950 3068 32956 3080
rect 33008 3068 33014 3120
rect 35986 3068 35992 3120
rect 36044 3108 36050 3120
rect 39942 3108 39948 3120
rect 36044 3080 39948 3108
rect 36044 3068 36050 3080
rect 39942 3068 39948 3080
rect 40000 3068 40006 3120
rect 40678 3068 40684 3120
rect 40736 3108 40742 3120
rect 44634 3108 44640 3120
rect 40736 3080 44640 3108
rect 40736 3068 40742 3080
rect 44634 3068 44640 3080
rect 44692 3068 44698 3120
rect 50154 3068 50160 3120
rect 50212 3108 50218 3120
rect 53926 3108 53932 3120
rect 50212 3080 53932 3108
rect 50212 3068 50218 3080
rect 53926 3068 53932 3080
rect 53984 3068 53990 3120
rect 135254 3068 135260 3120
rect 135312 3108 135318 3120
rect 137922 3108 137928 3120
rect 135312 3080 137928 3108
rect 135312 3068 135318 3080
rect 137922 3068 137928 3080
rect 137980 3068 137986 3120
rect 144730 3068 144736 3120
rect 144788 3108 144794 3120
rect 147306 3108 147312 3120
rect 144788 3080 147312 3108
rect 144788 3068 144794 3080
rect 147306 3068 147312 3080
rect 147364 3068 147370 3120
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 14274 3040 14280 3052
rect 10008 3012 14280 3040
rect 10008 3000 10014 3012
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 24762 3040 24768 3052
rect 20680 3012 24768 3040
rect 20680 3000 20686 3012
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 31754 3040 31760 3052
rect 27764 3012 31760 3040
rect 27764 3000 27770 3012
rect 31754 3000 31760 3012
rect 31812 3000 31818 3052
rect 32398 3000 32404 3052
rect 32456 3040 32462 3052
rect 36446 3040 36452 3052
rect 32456 3012 36452 3040
rect 32456 3000 32462 3012
rect 36446 3000 36452 3012
rect 36504 3000 36510 3052
rect 39574 3000 39580 3052
rect 39632 3040 39638 3052
rect 43438 3040 43444 3052
rect 39632 3012 43444 3040
rect 39632 3000 39638 3012
rect 43438 3000 43444 3012
rect 43496 3000 43502 3052
rect 48958 3000 48964 3052
rect 49016 3040 49022 3052
rect 52730 3040 52736 3052
rect 49016 3012 52736 3040
rect 49016 3000 49022 3012
rect 52730 3000 52736 3012
rect 52788 3000 52794 3052
rect 59630 3000 59636 3052
rect 59688 3040 59694 3052
rect 63310 3040 63316 3052
rect 59688 3012 63316 3040
rect 59688 3000 59694 3012
rect 63310 3000 63316 3012
rect 63368 3000 63374 3052
rect 69106 3000 69112 3052
rect 69164 3040 69170 3052
rect 72602 3040 72608 3052
rect 69164 3012 72608 3040
rect 69164 3000 69170 3012
rect 72602 3000 72608 3012
rect 72660 3000 72666 3052
rect 82078 3000 82084 3052
rect 82136 3040 82142 3052
rect 85482 3040 85488 3052
rect 82136 3012 85488 3040
rect 82136 3000 82142 3012
rect 85482 3000 85488 3012
rect 85540 3000 85546 3052
rect 106918 3000 106924 3052
rect 106976 3040 106982 3052
rect 109954 3040 109960 3052
rect 106976 3012 109960 3040
rect 106976 3000 106982 3012
rect 109954 3000 109960 3012
rect 110012 3000 110018 3052
rect 114002 3000 114008 3052
rect 114060 3040 114066 3052
rect 116946 3040 116952 3052
rect 114060 3012 116952 3040
rect 114060 3000 114066 3012
rect 116946 3000 116952 3012
rect 117004 3000 117010 3052
rect 128170 3000 128176 3052
rect 128228 3040 128234 3052
rect 130930 3040 130936 3052
rect 128228 3012 130936 3040
rect 128228 3000 128234 3012
rect 130930 3000 130936 3012
rect 130988 3000 130994 3052
rect 134150 3000 134156 3052
rect 134208 3040 134214 3052
rect 136818 3040 136824 3052
rect 134208 3012 136824 3040
rect 134208 3000 134214 3012
rect 136818 3000 136824 3012
rect 136876 3000 136882 3052
rect 143534 3000 143540 3052
rect 143592 3040 143598 3052
rect 146110 3040 146116 3052
rect 143592 3012 146116 3040
rect 143592 3000 143598 3012
rect 146110 3000 146116 3012
rect 146168 3000 146174 3052
rect 151814 3000 151820 3052
rect 151872 3040 151878 3052
rect 154298 3040 154304 3052
rect 151872 3012 154304 3040
rect 151872 3000 151878 3012
rect 154298 3000 154304 3012
rect 154356 3000 154362 3052
rect 4062 2932 4068 2984
rect 4120 2972 4126 2984
rect 8478 2972 8484 2984
rect 4120 2944 8484 2972
rect 4120 2932 4126 2944
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 13078 2972 13084 2984
rect 8812 2944 13084 2972
rect 8812 2932 8818 2944
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 18966 2972 18972 2984
rect 14792 2944 18972 2972
rect 14792 2932 14798 2944
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 21818 2932 21824 2984
rect 21876 2972 21882 2984
rect 25958 2972 25964 2984
rect 21876 2944 25964 2972
rect 21876 2932 21882 2944
rect 25958 2932 25964 2944
rect 26016 2932 26022 2984
rect 26510 2932 26516 2984
rect 26568 2972 26574 2984
rect 30558 2972 30564 2984
rect 26568 2944 30564 2972
rect 26568 2932 26574 2944
rect 30558 2932 30564 2944
rect 30616 2932 30622 2984
rect 33594 2932 33600 2984
rect 33652 2972 33658 2984
rect 37642 2972 37648 2984
rect 33652 2944 37648 2972
rect 33652 2932 33658 2944
rect 37642 2932 37648 2944
rect 37700 2932 37706 2984
rect 43070 2932 43076 2984
rect 43128 2972 43134 2984
rect 46934 2972 46940 2984
rect 43128 2944 46940 2972
rect 43128 2932 43134 2944
rect 46934 2932 46940 2944
rect 46992 2932 46998 2984
rect 51350 2932 51356 2984
rect 51408 2972 51414 2984
rect 55122 2972 55128 2984
rect 51408 2944 55128 2972
rect 51408 2932 51414 2944
rect 55122 2932 55128 2944
rect 55180 2932 55186 2984
rect 56042 2932 56048 2984
rect 56100 2972 56106 2984
rect 59814 2972 59820 2984
rect 56100 2944 59820 2972
rect 56100 2932 56106 2944
rect 59814 2932 59820 2944
rect 59872 2932 59878 2984
rect 60826 2932 60832 2984
rect 60884 2972 60890 2984
rect 64414 2972 64420 2984
rect 60884 2944 64420 2972
rect 60884 2932 60890 2944
rect 64414 2932 64420 2944
rect 64472 2932 64478 2984
rect 77386 2932 77392 2984
rect 77444 2972 77450 2984
rect 80790 2972 80796 2984
rect 77444 2944 80796 2972
rect 77444 2932 77450 2944
rect 80790 2932 80796 2944
rect 80848 2932 80854 2984
rect 80882 2932 80888 2984
rect 80940 2972 80946 2984
rect 84286 2972 84292 2984
rect 80940 2944 84292 2972
rect 80940 2932 80946 2944
rect 84286 2932 84292 2944
rect 84344 2932 84350 2984
rect 85666 2932 85672 2984
rect 85724 2972 85730 2984
rect 88978 2972 88984 2984
rect 85724 2944 88984 2972
rect 85724 2932 85730 2944
rect 88978 2932 88984 2944
rect 89036 2932 89042 2984
rect 89162 2932 89168 2984
rect 89220 2972 89226 2984
rect 92474 2972 92480 2984
rect 89220 2944 92480 2972
rect 89220 2932 89226 2944
rect 92474 2932 92480 2944
rect 92532 2932 92538 2984
rect 92750 2932 92756 2984
rect 92808 2972 92814 2984
rect 95970 2972 95976 2984
rect 92808 2944 95976 2972
rect 92808 2932 92814 2944
rect 95970 2932 95976 2944
rect 96028 2932 96034 2984
rect 96246 2932 96252 2984
rect 96304 2972 96310 2984
rect 99466 2972 99472 2984
rect 96304 2944 99472 2972
rect 96304 2932 96310 2944
rect 99466 2932 99472 2944
rect 99524 2932 99530 2984
rect 99834 2932 99840 2984
rect 99892 2972 99898 2984
rect 102962 2972 102968 2984
rect 99892 2944 102968 2972
rect 99892 2932 99898 2944
rect 102962 2932 102968 2944
rect 103020 2932 103026 2984
rect 108114 2932 108120 2984
rect 108172 2972 108178 2984
rect 111150 2972 111156 2984
rect 108172 2944 111156 2972
rect 108172 2932 108178 2944
rect 111150 2932 111156 2944
rect 111208 2932 111214 2984
rect 111610 2932 111616 2984
rect 111668 2972 111674 2984
rect 114646 2972 114652 2984
rect 111668 2944 114652 2972
rect 111668 2932 111674 2944
rect 114646 2932 114652 2944
rect 114704 2932 114710 2984
rect 117590 2932 117596 2984
rect 117648 2972 117654 2984
rect 120442 2972 120448 2984
rect 117648 2944 120448 2972
rect 117648 2932 117654 2944
rect 120442 2932 120448 2944
rect 120500 2932 120506 2984
rect 121086 2932 121092 2984
rect 121144 2972 121150 2984
rect 123938 2972 123944 2984
rect 121144 2944 123944 2972
rect 121144 2932 121150 2944
rect 123938 2932 123944 2944
rect 123996 2932 124002 2984
rect 124674 2932 124680 2984
rect 124732 2972 124738 2984
rect 127434 2972 127440 2984
rect 124732 2944 127440 2972
rect 124732 2932 124738 2944
rect 127434 2932 127440 2944
rect 127492 2932 127498 2984
rect 129366 2932 129372 2984
rect 129424 2972 129430 2984
rect 132126 2972 132132 2984
rect 129424 2944 132132 2972
rect 129424 2932 129430 2944
rect 132126 2932 132132 2944
rect 132184 2932 132190 2984
rect 132954 2932 132960 2984
rect 133012 2972 133018 2984
rect 135622 2972 135628 2984
rect 133012 2944 135628 2972
rect 133012 2932 133018 2944
rect 135622 2932 135628 2944
rect 135680 2932 135686 2984
rect 138842 2932 138848 2984
rect 138900 2972 138906 2984
rect 141418 2972 141424 2984
rect 138900 2944 141424 2972
rect 138900 2932 138906 2944
rect 141418 2932 141424 2944
rect 141476 2932 141482 2984
rect 142430 2932 142436 2984
rect 142488 2972 142494 2984
rect 144914 2972 144920 2984
rect 142488 2944 144920 2972
rect 142488 2932 142494 2944
rect 144914 2932 144920 2944
rect 144972 2932 144978 2984
rect 148318 2932 148324 2984
rect 148376 2972 148382 2984
rect 150802 2972 150808 2984
rect 148376 2944 150808 2972
rect 148376 2932 148382 2944
rect 150802 2932 150808 2944
rect 150860 2932 150866 2984
rect 154206 2932 154212 2984
rect 154264 2972 154270 2984
rect 156598 2972 156604 2984
rect 154264 2944 156604 2972
rect 154264 2932 154270 2944
rect 156598 2932 156604 2944
rect 156656 2932 156662 2984
rect 158990 2932 158996 2984
rect 159048 2972 159054 2984
rect 161290 2972 161296 2984
rect 159048 2944 161296 2972
rect 159048 2932 159054 2944
rect 161290 2932 161296 2944
rect 161348 2932 161354 2984
rect 162486 2932 162492 2984
rect 162544 2972 162550 2984
rect 164786 2972 164792 2984
rect 162544 2944 164792 2972
rect 162544 2932 162550 2944
rect 164786 2932 164792 2944
rect 164844 2932 164850 2984
rect 167178 2932 167184 2984
rect 167236 2972 167242 2984
rect 169478 2972 169484 2984
rect 167236 2944 169484 2972
rect 167236 2932 167242 2944
rect 169478 2932 169484 2944
rect 169536 2932 169542 2984
rect 174262 2932 174268 2984
rect 174320 2972 174326 2984
rect 176470 2972 176476 2984
rect 174320 2944 176476 2972
rect 174320 2932 174326 2944
rect 176470 2932 176476 2944
rect 176528 2932 176534 2984
rect 177850 2932 177856 2984
rect 177908 2972 177914 2984
rect 179966 2972 179972 2984
rect 177908 2944 179972 2972
rect 177908 2932 177914 2944
rect 179966 2932 179972 2944
rect 180024 2932 180030 2984
rect 181438 2932 181444 2984
rect 181496 2972 181502 2984
rect 183462 2972 183468 2984
rect 181496 2944 183468 2972
rect 181496 2932 181502 2944
rect 183462 2932 183468 2944
rect 183520 2932 183526 2984
rect 192018 2932 192024 2984
rect 192076 2972 192082 2984
rect 193950 2972 193956 2984
rect 192076 2944 193956 2972
rect 192076 2932 192082 2944
rect 193950 2932 193956 2944
rect 194008 2932 194014 2984
rect 199102 2932 199108 2984
rect 199160 2972 199166 2984
rect 200942 2972 200948 2984
rect 199160 2944 200948 2972
rect 199160 2932 199166 2944
rect 200942 2932 200948 2944
rect 201000 2932 201006 2984
rect 202690 2932 202696 2984
rect 202748 2972 202754 2984
rect 204438 2972 204444 2984
rect 202748 2944 204444 2972
rect 202748 2932 202754 2944
rect 204438 2932 204444 2944
rect 204496 2932 204502 2984
rect 206186 2932 206192 2984
rect 206244 2972 206250 2984
rect 207934 2972 207940 2984
rect 206244 2944 207940 2972
rect 206244 2932 206250 2944
rect 207934 2932 207940 2944
rect 207992 2932 207998 2984
rect 209774 2932 209780 2984
rect 209832 2972 209838 2984
rect 211430 2972 211436 2984
rect 209832 2944 211436 2972
rect 209832 2932 209838 2944
rect 211430 2932 211436 2944
rect 211488 2932 211494 2984
rect 215662 2932 215668 2984
rect 215720 2972 215726 2984
rect 217318 2972 217324 2984
rect 215720 2944 217324 2972
rect 215720 2932 215726 2944
rect 217318 2932 217324 2944
rect 217376 2932 217382 2984
rect 226334 2932 226340 2984
rect 226392 2972 226398 2984
rect 227806 2972 227812 2984
rect 226392 2944 227812 2972
rect 226392 2932 226398 2944
rect 227806 2932 227812 2944
rect 227864 2932 227870 2984
rect 229830 2932 229836 2984
rect 229888 2972 229894 2984
rect 231302 2972 231308 2984
rect 229888 2944 231308 2972
rect 229888 2932 229894 2944
rect 231302 2932 231308 2944
rect 231360 2932 231366 2984
rect 233418 2932 233424 2984
rect 233476 2972 233482 2984
rect 234798 2972 234804 2984
rect 233476 2944 234804 2972
rect 233476 2932 233482 2944
rect 234798 2932 234804 2944
rect 234856 2932 234862 2984
rect 238110 2932 238116 2984
rect 238168 2972 238174 2984
rect 239398 2972 239404 2984
rect 238168 2944 239404 2972
rect 238168 2932 238174 2944
rect 239398 2932 239404 2944
rect 239456 2932 239462 2984
rect 241698 2932 241704 2984
rect 241756 2972 241762 2984
rect 242986 2972 242992 2984
rect 241756 2944 242992 2972
rect 241756 2932 241762 2944
rect 242986 2932 242992 2944
rect 243044 2932 243050 2984
rect 246390 2932 246396 2984
rect 246448 2972 246454 2984
rect 247586 2972 247592 2984
rect 246448 2944 247592 2972
rect 246448 2932 246454 2944
rect 247586 2932 247592 2944
rect 247644 2932 247650 2984
rect 248874 2932 248880 2984
rect 248932 2972 248938 2984
rect 249978 2972 249984 2984
rect 248932 2944 249984 2972
rect 248932 2932 248938 2944
rect 249978 2932 249984 2944
rect 250036 2932 250042 2984
rect 252370 2932 252376 2984
rect 252428 2972 252434 2984
rect 253474 2972 253480 2984
rect 252428 2944 253480 2972
rect 252428 2932 252434 2944
rect 253474 2932 253480 2944
rect 253532 2932 253538 2984
rect 570782 2932 570788 2984
rect 570840 2972 570846 2984
rect 573910 2972 573916 2984
rect 570840 2944 573916 2972
rect 570840 2932 570846 2944
rect 573910 2932 573916 2944
rect 573968 2932 573974 2984
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 7282 2904 7288 2916
rect 2924 2876 7288 2904
rect 2924 2864 2930 2876
rect 7282 2864 7288 2876
rect 7340 2864 7346 2916
rect 12342 2864 12348 2916
rect 12400 2904 12406 2916
rect 16482 2904 16488 2916
rect 12400 2876 16488 2904
rect 12400 2864 12406 2876
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 23566 2904 23572 2916
rect 19484 2876 23572 2904
rect 19484 2864 19490 2876
rect 23566 2864 23572 2876
rect 23624 2864 23630 2916
rect 24210 2864 24216 2916
rect 24268 2904 24274 2916
rect 28258 2904 28264 2916
rect 24268 2876 28264 2904
rect 24268 2864 24274 2876
rect 28258 2864 28264 2876
rect 28316 2864 28322 2916
rect 30098 2864 30104 2916
rect 30156 2904 30162 2916
rect 34146 2904 34152 2916
rect 30156 2876 34152 2904
rect 30156 2864 30162 2876
rect 34146 2864 34152 2876
rect 34204 2864 34210 2916
rect 37182 2864 37188 2916
rect 37240 2904 37246 2916
rect 41138 2904 41144 2916
rect 37240 2876 41144 2904
rect 37240 2864 37246 2876
rect 41138 2864 41144 2876
rect 41196 2864 41202 2916
rect 41874 2864 41880 2916
rect 41932 2904 41938 2916
rect 45738 2904 45744 2916
rect 41932 2876 45744 2904
rect 41932 2864 41938 2876
rect 45738 2864 45744 2876
rect 45796 2864 45802 2916
rect 47854 2864 47860 2916
rect 47912 2904 47918 2916
rect 51626 2904 51632 2916
rect 47912 2876 51632 2904
rect 47912 2864 47918 2876
rect 51626 2864 51632 2876
rect 51684 2864 51690 2916
rect 53742 2864 53748 2916
rect 53800 2904 53806 2916
rect 57422 2904 57428 2916
rect 53800 2876 57428 2904
rect 53800 2864 53806 2876
rect 57422 2864 57428 2876
rect 57480 2864 57486 2916
rect 58434 2864 58440 2916
rect 58492 2904 58498 2916
rect 62114 2904 62120 2916
rect 58492 2876 62120 2904
rect 58492 2864 58498 2876
rect 62114 2864 62120 2876
rect 62172 2864 62178 2916
rect 63218 2864 63224 2916
rect 63276 2904 63282 2916
rect 66806 2904 66812 2916
rect 63276 2876 66812 2904
rect 63276 2864 63282 2876
rect 66806 2864 66812 2876
rect 66864 2864 66870 2916
rect 72602 2864 72608 2916
rect 72660 2904 72666 2916
rect 76098 2904 76104 2916
rect 72660 2876 76104 2904
rect 72660 2864 72666 2876
rect 76098 2864 76104 2876
rect 76156 2864 76162 2916
rect 76190 2864 76196 2916
rect 76248 2904 76254 2916
rect 79594 2904 79600 2916
rect 76248 2876 79600 2904
rect 76248 2864 76254 2876
rect 79594 2864 79600 2876
rect 79652 2864 79658 2916
rect 79686 2864 79692 2916
rect 79744 2904 79750 2916
rect 83090 2904 83096 2916
rect 79744 2876 83096 2904
rect 79744 2864 79750 2876
rect 83090 2864 83096 2876
rect 83148 2864 83154 2916
rect 84470 2864 84476 2916
rect 84528 2904 84534 2916
rect 87782 2904 87788 2916
rect 84528 2876 87788 2904
rect 84528 2864 84534 2876
rect 87782 2864 87788 2876
rect 87840 2864 87846 2916
rect 87966 2864 87972 2916
rect 88024 2904 88030 2916
rect 91278 2904 91284 2916
rect 88024 2876 91284 2904
rect 88024 2864 88030 2876
rect 91278 2864 91284 2876
rect 91336 2864 91342 2916
rect 91554 2864 91560 2916
rect 91612 2904 91618 2916
rect 94774 2904 94780 2916
rect 91612 2876 94780 2904
rect 91612 2864 91618 2876
rect 94774 2864 94780 2876
rect 94832 2864 94838 2916
rect 95142 2864 95148 2916
rect 95200 2904 95206 2916
rect 98270 2904 98276 2916
rect 95200 2876 98276 2904
rect 95200 2864 95206 2876
rect 98270 2864 98276 2876
rect 98328 2864 98334 2916
rect 98638 2864 98644 2916
rect 98696 2904 98702 2916
rect 101766 2904 101772 2916
rect 98696 2876 101772 2904
rect 98696 2864 98702 2876
rect 101766 2864 101772 2876
rect 101824 2864 101830 2916
rect 102226 2864 102232 2916
rect 102284 2904 102290 2916
rect 105262 2904 105268 2916
rect 102284 2876 105268 2904
rect 102284 2864 102290 2876
rect 105262 2864 105268 2876
rect 105320 2864 105326 2916
rect 105722 2864 105728 2916
rect 105780 2904 105786 2916
rect 108758 2904 108764 2916
rect 105780 2876 108764 2904
rect 105780 2864 105786 2876
rect 108758 2864 108764 2876
rect 108816 2864 108822 2916
rect 110506 2864 110512 2916
rect 110564 2904 110570 2916
rect 113450 2904 113456 2916
rect 110564 2876 113456 2904
rect 110564 2864 110570 2876
rect 113450 2864 113456 2876
rect 113508 2864 113514 2916
rect 115750 2904 115756 2916
rect 114296 2876 115756 2904
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 1728 2808 4200 2836
rect 1728 2796 1734 2808
rect 4172 2768 4200 2808
rect 5258 2796 5264 2848
rect 5316 2836 5322 2848
rect 5316 2808 6914 2836
rect 5316 2796 5322 2808
rect 6086 2768 6092 2780
rect 4172 2740 6092 2768
rect 6086 2728 6092 2740
rect 6144 2728 6150 2780
rect 6886 2768 6914 2808
rect 7650 2796 7656 2848
rect 7708 2836 7714 2848
rect 11974 2836 11980 2848
rect 7708 2808 11980 2836
rect 7708 2796 7714 2808
rect 11974 2796 11980 2808
rect 12032 2796 12038 2848
rect 13538 2796 13544 2848
rect 13596 2836 13602 2848
rect 17770 2836 17776 2848
rect 13596 2808 17776 2836
rect 13596 2796 13602 2808
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18230 2796 18236 2848
rect 18288 2836 18294 2848
rect 22462 2836 22468 2848
rect 18288 2808 22468 2836
rect 18288 2796 18294 2808
rect 22462 2796 22468 2808
rect 22520 2796 22526 2848
rect 23014 2796 23020 2848
rect 23072 2836 23078 2848
rect 27062 2836 27068 2848
rect 23072 2808 27068 2836
rect 23072 2796 23078 2808
rect 27062 2796 27068 2808
rect 27120 2796 27126 2848
rect 31294 2796 31300 2848
rect 31352 2836 31358 2848
rect 35250 2836 35256 2848
rect 31352 2808 35256 2836
rect 31352 2796 31358 2808
rect 35250 2796 35256 2808
rect 35308 2796 35314 2848
rect 38378 2796 38384 2848
rect 38436 2836 38442 2848
rect 42242 2836 42248 2848
rect 38436 2808 42248 2836
rect 38436 2796 38442 2808
rect 42242 2796 42248 2808
rect 42300 2796 42306 2848
rect 44266 2796 44272 2848
rect 44324 2836 44330 2848
rect 48130 2836 48136 2848
rect 44324 2808 48136 2836
rect 44324 2796 44330 2808
rect 48130 2796 48136 2808
rect 48188 2796 48194 2848
rect 52546 2796 52552 2848
rect 52604 2836 52610 2848
rect 56226 2836 56232 2848
rect 52604 2808 56232 2836
rect 52604 2796 52610 2808
rect 56226 2796 56232 2808
rect 56284 2796 56290 2848
rect 57238 2796 57244 2848
rect 57296 2836 57302 2848
rect 60918 2836 60924 2848
rect 57296 2808 60924 2836
rect 57296 2796 57302 2808
rect 60918 2796 60924 2808
rect 60976 2796 60982 2848
rect 62022 2796 62028 2848
rect 62080 2836 62086 2848
rect 65610 2836 65616 2848
rect 62080 2808 65616 2836
rect 62080 2796 62086 2808
rect 65610 2796 65616 2808
rect 65668 2796 65674 2848
rect 67910 2796 67916 2848
rect 67968 2836 67974 2848
rect 71406 2836 71412 2848
rect 67968 2808 71412 2836
rect 67968 2796 67974 2808
rect 71406 2796 71412 2808
rect 71464 2796 71470 2848
rect 71498 2796 71504 2848
rect 71556 2836 71562 2848
rect 74902 2836 74908 2848
rect 71556 2808 74908 2836
rect 71556 2796 71562 2808
rect 74902 2796 74908 2808
rect 74960 2796 74966 2848
rect 74994 2796 75000 2848
rect 75052 2836 75058 2848
rect 78398 2836 78404 2848
rect 75052 2808 78404 2836
rect 75052 2796 75058 2808
rect 78398 2796 78404 2808
rect 78456 2796 78462 2848
rect 78582 2796 78588 2848
rect 78640 2836 78646 2848
rect 81894 2836 81900 2848
rect 78640 2808 81900 2836
rect 78640 2796 78646 2808
rect 81894 2796 81900 2808
rect 81952 2796 81958 2848
rect 83274 2796 83280 2848
rect 83332 2836 83338 2848
rect 86586 2836 86592 2848
rect 83332 2808 86592 2836
rect 83332 2796 83338 2808
rect 86586 2796 86592 2808
rect 86644 2796 86650 2848
rect 86862 2796 86868 2848
rect 86920 2836 86926 2848
rect 90082 2836 90088 2848
rect 86920 2808 90088 2836
rect 86920 2796 86926 2808
rect 90082 2796 90088 2808
rect 90140 2796 90146 2848
rect 90358 2796 90364 2848
rect 90416 2836 90422 2848
rect 93578 2836 93584 2848
rect 90416 2808 93584 2836
rect 90416 2796 90422 2808
rect 93578 2796 93584 2808
rect 93636 2796 93642 2848
rect 93946 2796 93952 2848
rect 94004 2836 94010 2848
rect 97074 2836 97080 2848
rect 94004 2808 97080 2836
rect 94004 2796 94010 2808
rect 97074 2796 97080 2808
rect 97132 2796 97138 2848
rect 97442 2796 97448 2848
rect 97500 2836 97506 2848
rect 100570 2836 100576 2848
rect 97500 2808 100576 2836
rect 97500 2796 97506 2808
rect 100570 2796 100576 2808
rect 100628 2796 100634 2848
rect 101030 2796 101036 2848
rect 101088 2836 101094 2848
rect 104066 2836 104072 2848
rect 101088 2808 104072 2836
rect 101088 2796 101094 2808
rect 104066 2796 104072 2808
rect 104124 2796 104130 2848
rect 104526 2796 104532 2848
rect 104584 2836 104590 2848
rect 107562 2836 107568 2848
rect 104584 2808 107568 2836
rect 104584 2796 104590 2808
rect 107562 2796 107568 2808
rect 107620 2796 107626 2848
rect 109310 2796 109316 2848
rect 109368 2836 109374 2848
rect 112254 2836 112260 2848
rect 109368 2808 112260 2836
rect 109368 2796 109374 2808
rect 112254 2796 112260 2808
rect 112312 2796 112318 2848
rect 112806 2796 112812 2848
rect 112864 2836 112870 2848
rect 114296 2836 114324 2876
rect 115750 2864 115756 2876
rect 115808 2864 115814 2916
rect 116394 2864 116400 2916
rect 116452 2904 116458 2916
rect 119246 2904 119252 2916
rect 116452 2876 119252 2904
rect 116452 2864 116458 2876
rect 119246 2864 119252 2876
rect 119304 2864 119310 2916
rect 119890 2864 119896 2916
rect 119948 2904 119954 2916
rect 122742 2904 122748 2916
rect 119948 2876 122748 2904
rect 119948 2864 119954 2876
rect 122742 2864 122748 2876
rect 122800 2864 122806 2916
rect 123478 2864 123484 2916
rect 123536 2904 123542 2916
rect 126238 2904 126244 2916
rect 123536 2876 126244 2904
rect 123536 2864 123542 2876
rect 126238 2864 126244 2876
rect 126296 2864 126302 2916
rect 126974 2864 126980 2916
rect 127032 2904 127038 2916
rect 129734 2904 129740 2916
rect 127032 2876 129740 2904
rect 127032 2864 127038 2876
rect 129734 2864 129740 2876
rect 129792 2864 129798 2916
rect 131758 2864 131764 2916
rect 131816 2904 131822 2916
rect 134426 2904 134432 2916
rect 131816 2876 134432 2904
rect 131816 2864 131822 2876
rect 134426 2864 134432 2876
rect 134484 2864 134490 2916
rect 137646 2864 137652 2916
rect 137704 2904 137710 2916
rect 140314 2904 140320 2916
rect 137704 2876 140320 2904
rect 137704 2864 137710 2876
rect 140314 2864 140320 2876
rect 140372 2864 140378 2916
rect 141234 2864 141240 2916
rect 141292 2904 141298 2916
rect 143810 2904 143816 2916
rect 141292 2876 143816 2904
rect 141292 2864 141298 2876
rect 143810 2864 143816 2876
rect 143868 2864 143874 2916
rect 147122 2864 147128 2916
rect 147180 2904 147186 2916
rect 149606 2904 149612 2916
rect 147180 2876 149612 2904
rect 147180 2864 147186 2876
rect 149606 2864 149612 2876
rect 149664 2864 149670 2916
rect 150618 2864 150624 2916
rect 150676 2904 150682 2916
rect 153102 2904 153108 2916
rect 150676 2876 153108 2904
rect 150676 2864 150682 2876
rect 153102 2864 153108 2876
rect 153160 2864 153166 2916
rect 163682 2864 163688 2916
rect 163740 2904 163746 2916
rect 165982 2904 165988 2916
rect 163740 2876 165988 2904
rect 163740 2864 163746 2876
rect 165982 2864 165988 2876
rect 166040 2864 166046 2916
rect 166074 2864 166080 2916
rect 166132 2904 166138 2916
rect 168282 2904 168288 2916
rect 166132 2876 168288 2904
rect 166132 2864 166138 2876
rect 168282 2864 168288 2876
rect 168340 2864 168346 2916
rect 169570 2864 169576 2916
rect 169628 2904 169634 2916
rect 171778 2904 171784 2916
rect 169628 2876 171784 2904
rect 169628 2864 169634 2876
rect 171778 2864 171784 2876
rect 171836 2864 171842 2916
rect 172974 2904 172980 2916
rect 171888 2876 172980 2904
rect 112864 2808 114324 2836
rect 112864 2796 112870 2808
rect 115198 2796 115204 2848
rect 115256 2836 115262 2848
rect 118142 2836 118148 2848
rect 115256 2808 118148 2836
rect 115256 2796 115262 2808
rect 118142 2796 118148 2808
rect 118200 2796 118206 2848
rect 118786 2796 118792 2848
rect 118844 2836 118850 2848
rect 121638 2836 121644 2848
rect 118844 2808 121644 2836
rect 118844 2796 118850 2808
rect 121638 2796 121644 2808
rect 121696 2796 121702 2848
rect 122282 2796 122288 2848
rect 122340 2836 122346 2848
rect 125134 2836 125140 2848
rect 122340 2808 125140 2836
rect 122340 2796 122346 2808
rect 125134 2796 125140 2808
rect 125192 2796 125198 2848
rect 125870 2796 125876 2848
rect 125928 2836 125934 2848
rect 128630 2836 128636 2848
rect 125928 2808 128636 2836
rect 125928 2796 125934 2808
rect 128630 2796 128636 2808
rect 128688 2796 128694 2848
rect 130562 2796 130568 2848
rect 130620 2836 130626 2848
rect 133230 2836 133236 2848
rect 130620 2808 133236 2836
rect 130620 2796 130626 2808
rect 133230 2796 133236 2808
rect 133288 2796 133294 2848
rect 136450 2796 136456 2848
rect 136508 2836 136514 2848
rect 139118 2836 139124 2848
rect 136508 2808 139124 2836
rect 136508 2796 136514 2808
rect 139118 2796 139124 2808
rect 139176 2796 139182 2848
rect 140038 2796 140044 2848
rect 140096 2836 140102 2848
rect 142614 2836 142620 2848
rect 140096 2808 142620 2836
rect 140096 2796 140102 2808
rect 142614 2796 142620 2808
rect 142672 2796 142678 2848
rect 145926 2796 145932 2848
rect 145984 2836 145990 2848
rect 148410 2836 148416 2848
rect 145984 2808 148416 2836
rect 145984 2796 145990 2808
rect 148410 2796 148416 2808
rect 148468 2796 148474 2848
rect 149514 2796 149520 2848
rect 149572 2836 149578 2848
rect 151906 2836 151912 2848
rect 149572 2808 151912 2836
rect 149572 2796 149578 2808
rect 151906 2796 151912 2808
rect 151964 2796 151970 2848
rect 156598 2796 156604 2848
rect 156656 2836 156662 2848
rect 158898 2836 158904 2848
rect 156656 2808 158904 2836
rect 156656 2796 156662 2808
rect 158898 2796 158904 2808
rect 158956 2796 158962 2848
rect 161290 2796 161296 2848
rect 161348 2836 161354 2848
rect 163590 2836 163596 2848
rect 161348 2808 163596 2836
rect 161348 2796 161354 2808
rect 163590 2796 163596 2808
rect 163648 2796 163654 2848
rect 164878 2796 164884 2848
rect 164936 2836 164942 2848
rect 167086 2836 167092 2848
rect 164936 2808 167092 2836
rect 164936 2796 164942 2808
rect 167086 2796 167092 2808
rect 167144 2796 167150 2848
rect 168374 2796 168380 2848
rect 168432 2836 168438 2848
rect 170582 2836 170588 2848
rect 168432 2808 170588 2836
rect 168432 2796 168438 2808
rect 170582 2796 170588 2808
rect 170640 2796 170646 2848
rect 170766 2796 170772 2848
rect 170824 2836 170830 2848
rect 171888 2836 171916 2876
rect 172974 2864 172980 2876
rect 173032 2864 173038 2916
rect 173158 2864 173164 2916
rect 173216 2904 173222 2916
rect 175274 2904 175280 2916
rect 173216 2876 175280 2904
rect 173216 2864 173222 2876
rect 175274 2864 175280 2876
rect 175332 2864 175338 2916
rect 176654 2864 176660 2916
rect 176712 2904 176718 2916
rect 178770 2904 178776 2916
rect 176712 2876 178776 2904
rect 176712 2864 176718 2876
rect 178770 2864 178776 2876
rect 178828 2864 178834 2916
rect 180242 2864 180248 2916
rect 180300 2904 180306 2916
rect 182266 2904 182272 2916
rect 180300 2876 182272 2904
rect 180300 2864 180306 2876
rect 182266 2864 182272 2876
rect 182324 2864 182330 2916
rect 183738 2864 183744 2916
rect 183796 2904 183802 2916
rect 185762 2904 185768 2916
rect 183796 2876 185768 2904
rect 183796 2864 183802 2876
rect 185762 2864 185768 2876
rect 185820 2864 185826 2916
rect 186130 2864 186136 2916
rect 186188 2904 186194 2916
rect 188154 2904 188160 2916
rect 186188 2876 188160 2904
rect 186188 2864 186194 2876
rect 188154 2864 188160 2876
rect 188212 2864 188218 2916
rect 188522 2864 188528 2916
rect 188580 2904 188586 2916
rect 190454 2904 190460 2916
rect 188580 2876 190460 2904
rect 188580 2864 188586 2876
rect 190454 2864 190460 2876
rect 190512 2864 190518 2916
rect 191650 2904 191656 2916
rect 190748 2876 191656 2904
rect 170824 2808 171916 2836
rect 170824 2796 170830 2808
rect 171962 2796 171968 2848
rect 172020 2836 172026 2848
rect 174078 2836 174084 2848
rect 172020 2808 174084 2836
rect 172020 2796 172026 2808
rect 174078 2796 174084 2808
rect 174136 2796 174142 2848
rect 175458 2796 175464 2848
rect 175516 2836 175522 2848
rect 177574 2836 177580 2848
rect 175516 2808 177580 2836
rect 175516 2796 175522 2808
rect 177574 2796 177580 2808
rect 177632 2796 177638 2848
rect 179046 2796 179052 2848
rect 179104 2836 179110 2848
rect 181070 2836 181076 2848
rect 179104 2808 181076 2836
rect 179104 2796 179110 2808
rect 181070 2796 181076 2808
rect 181128 2796 181134 2848
rect 182542 2796 182548 2848
rect 182600 2836 182606 2848
rect 184566 2836 184572 2848
rect 182600 2808 184572 2836
rect 182600 2796 182606 2808
rect 184566 2796 184572 2808
rect 184624 2796 184630 2848
rect 184934 2796 184940 2848
rect 184992 2836 184998 2848
rect 186958 2836 186964 2848
rect 184992 2808 186964 2836
rect 184992 2796 184998 2808
rect 186958 2796 186964 2808
rect 187016 2796 187022 2848
rect 187326 2796 187332 2848
rect 187384 2836 187390 2848
rect 189258 2836 189264 2848
rect 187384 2808 189264 2836
rect 187384 2796 187390 2808
rect 189258 2796 189264 2808
rect 189316 2796 189322 2848
rect 189718 2796 189724 2848
rect 189776 2836 189782 2848
rect 190748 2836 190776 2876
rect 191650 2864 191656 2876
rect 191708 2864 191714 2916
rect 193214 2864 193220 2916
rect 193272 2904 193278 2916
rect 195146 2904 195152 2916
rect 193272 2876 195152 2904
rect 193272 2864 193278 2876
rect 195146 2864 195152 2876
rect 195204 2864 195210 2916
rect 195606 2864 195612 2916
rect 195664 2904 195670 2916
rect 197446 2904 197452 2916
rect 195664 2876 197452 2904
rect 195664 2864 195670 2876
rect 197446 2864 197452 2876
rect 197504 2864 197510 2916
rect 197906 2864 197912 2916
rect 197964 2904 197970 2916
rect 199746 2904 199752 2916
rect 197964 2876 199752 2904
rect 197964 2864 197970 2876
rect 199746 2864 199752 2876
rect 199804 2864 199810 2916
rect 200298 2864 200304 2916
rect 200356 2904 200362 2916
rect 202138 2904 202144 2916
rect 200356 2876 202144 2904
rect 200356 2864 200362 2876
rect 202138 2864 202144 2876
rect 202196 2864 202202 2916
rect 203886 2864 203892 2916
rect 203944 2904 203950 2916
rect 205634 2904 205640 2916
rect 203944 2876 205640 2904
rect 203944 2864 203950 2876
rect 205634 2864 205640 2876
rect 205692 2864 205698 2916
rect 207382 2864 207388 2916
rect 207440 2904 207446 2916
rect 209130 2904 209136 2916
rect 207440 2876 209136 2904
rect 207440 2864 207446 2876
rect 209130 2864 209136 2876
rect 209188 2864 209194 2916
rect 210970 2864 210976 2916
rect 211028 2904 211034 2916
rect 212626 2904 212632 2916
rect 211028 2876 212632 2904
rect 211028 2864 211034 2876
rect 212626 2864 212632 2876
rect 212684 2864 212690 2916
rect 213362 2864 213368 2916
rect 213420 2904 213426 2916
rect 214926 2904 214932 2916
rect 213420 2876 214932 2904
rect 213420 2864 213426 2876
rect 214926 2864 214932 2876
rect 214984 2864 214990 2916
rect 216858 2864 216864 2916
rect 216916 2904 216922 2916
rect 218422 2904 218428 2916
rect 216916 2876 218428 2904
rect 216916 2864 216922 2876
rect 218422 2864 218428 2876
rect 218480 2864 218486 2916
rect 219250 2864 219256 2916
rect 219308 2904 219314 2916
rect 220814 2904 220820 2916
rect 219308 2876 220820 2904
rect 219308 2864 219314 2876
rect 220814 2864 220820 2876
rect 220872 2864 220878 2916
rect 221550 2864 221556 2916
rect 221608 2904 221614 2916
rect 223114 2904 223120 2916
rect 221608 2876 223120 2904
rect 221608 2864 221614 2876
rect 223114 2864 223120 2876
rect 223172 2864 223178 2916
rect 223942 2864 223948 2916
rect 224000 2904 224006 2916
rect 225414 2904 225420 2916
rect 224000 2876 225420 2904
rect 224000 2864 224006 2876
rect 225414 2864 225420 2876
rect 225472 2864 225478 2916
rect 227530 2864 227536 2916
rect 227588 2904 227594 2916
rect 228910 2904 228916 2916
rect 227588 2876 228916 2904
rect 227588 2864 227594 2876
rect 228910 2864 228916 2876
rect 228968 2864 228974 2916
rect 231026 2864 231032 2916
rect 231084 2904 231090 2916
rect 232406 2904 232412 2916
rect 231084 2876 232412 2904
rect 231084 2864 231090 2876
rect 232406 2864 232412 2876
rect 232464 2864 232470 2916
rect 234614 2864 234620 2916
rect 234672 2904 234678 2916
rect 235902 2904 235908 2916
rect 234672 2876 235908 2904
rect 234672 2864 234678 2876
rect 235902 2864 235908 2876
rect 235960 2864 235966 2916
rect 237006 2864 237012 2916
rect 237064 2904 237070 2916
rect 238294 2904 238300 2916
rect 237064 2876 238300 2904
rect 237064 2864 237070 2876
rect 238294 2864 238300 2876
rect 238352 2864 238358 2916
rect 240502 2864 240508 2916
rect 240560 2904 240566 2916
rect 241790 2904 241796 2916
rect 240560 2876 241796 2904
rect 240560 2864 240566 2876
rect 241790 2864 241796 2876
rect 241848 2864 241854 2916
rect 245194 2864 245200 2916
rect 245252 2904 245258 2916
rect 246482 2904 246488 2916
rect 245252 2876 246488 2904
rect 245252 2864 245258 2876
rect 246482 2864 246488 2876
rect 246540 2864 246546 2916
rect 540422 2864 540428 2916
rect 540480 2904 540486 2916
rect 543182 2904 543188 2916
rect 540480 2876 543188 2904
rect 540480 2864 540486 2876
rect 543182 2864 543188 2876
rect 543240 2864 543246 2916
rect 547414 2864 547420 2916
rect 547472 2904 547478 2916
rect 550266 2904 550272 2916
rect 547472 2876 550272 2904
rect 547472 2864 547478 2876
rect 550266 2864 550272 2876
rect 550324 2864 550330 2916
rect 553394 2864 553400 2916
rect 553452 2904 553458 2916
rect 556154 2904 556160 2916
rect 553452 2876 556160 2904
rect 553452 2864 553458 2876
rect 556154 2864 556160 2876
rect 556212 2864 556218 2916
rect 561674 2864 561680 2916
rect 561732 2904 561738 2916
rect 564434 2904 564440 2916
rect 561732 2876 564440 2904
rect 561732 2864 561738 2876
rect 564434 2864 564440 2876
rect 564492 2864 564498 2916
rect 568574 2864 568580 2916
rect 568632 2904 568638 2916
rect 571518 2904 571524 2916
rect 568632 2876 571524 2904
rect 568632 2864 568638 2876
rect 571518 2864 571524 2876
rect 571576 2864 571582 2916
rect 189776 2808 190776 2836
rect 189776 2796 189782 2808
rect 190822 2796 190828 2848
rect 190880 2836 190886 2848
rect 192754 2836 192760 2848
rect 190880 2808 192760 2836
rect 190880 2796 190886 2808
rect 192754 2796 192760 2808
rect 192812 2796 192818 2848
rect 194410 2796 194416 2848
rect 194468 2836 194474 2848
rect 196250 2836 196256 2848
rect 194468 2808 196256 2836
rect 194468 2796 194474 2808
rect 196250 2796 196256 2808
rect 196308 2796 196314 2848
rect 196802 2796 196808 2848
rect 196860 2836 196866 2848
rect 198642 2836 198648 2848
rect 196860 2808 198648 2836
rect 196860 2796 196866 2808
rect 198642 2796 198648 2808
rect 198700 2796 198706 2848
rect 201494 2796 201500 2848
rect 201552 2836 201558 2848
rect 203242 2836 203248 2848
rect 201552 2808 203248 2836
rect 201552 2796 201558 2808
rect 203242 2796 203248 2808
rect 203300 2796 203306 2848
rect 205082 2796 205088 2848
rect 205140 2836 205146 2848
rect 206738 2836 206744 2848
rect 205140 2808 206744 2836
rect 205140 2796 205146 2808
rect 206738 2796 206744 2808
rect 206796 2796 206802 2848
rect 208578 2796 208584 2848
rect 208636 2836 208642 2848
rect 210234 2836 210240 2848
rect 208636 2808 210240 2836
rect 208636 2796 208642 2808
rect 210234 2796 210240 2808
rect 210292 2796 210298 2848
rect 212166 2796 212172 2848
rect 212224 2836 212230 2848
rect 213730 2836 213736 2848
rect 212224 2808 213736 2836
rect 212224 2796 212230 2808
rect 213730 2796 213736 2808
rect 213788 2796 213794 2848
rect 214466 2796 214472 2848
rect 214524 2836 214530 2848
rect 216122 2836 216128 2848
rect 214524 2808 216128 2836
rect 214524 2796 214530 2808
rect 216122 2796 216128 2808
rect 216180 2796 216186 2848
rect 218054 2796 218060 2848
rect 218112 2836 218118 2848
rect 219618 2836 219624 2848
rect 218112 2808 219624 2836
rect 218112 2796 218118 2808
rect 219618 2796 219624 2808
rect 219676 2796 219682 2848
rect 220446 2796 220452 2848
rect 220504 2836 220510 2848
rect 221918 2836 221924 2848
rect 220504 2808 221924 2836
rect 220504 2796 220510 2808
rect 221918 2796 221924 2808
rect 221976 2796 221982 2848
rect 222746 2796 222752 2848
rect 222804 2836 222810 2848
rect 224310 2836 224316 2848
rect 222804 2808 224316 2836
rect 222804 2796 222810 2808
rect 224310 2796 224316 2808
rect 224368 2796 224374 2848
rect 225138 2796 225144 2848
rect 225196 2836 225202 2848
rect 226610 2836 226616 2848
rect 225196 2808 226616 2836
rect 225196 2796 225202 2808
rect 226610 2796 226616 2808
rect 226668 2796 226674 2848
rect 228726 2796 228732 2848
rect 228784 2836 228790 2848
rect 230106 2836 230112 2848
rect 228784 2808 230112 2836
rect 228784 2796 228790 2808
rect 230106 2796 230112 2808
rect 230164 2796 230170 2848
rect 232222 2796 232228 2848
rect 232280 2836 232286 2848
rect 233602 2836 233608 2848
rect 232280 2808 233608 2836
rect 232280 2796 232286 2808
rect 233602 2796 233608 2808
rect 233660 2796 233666 2848
rect 235810 2796 235816 2848
rect 235868 2836 235874 2848
rect 237098 2836 237104 2848
rect 235868 2808 237104 2836
rect 235868 2796 235874 2808
rect 237098 2796 237104 2808
rect 237156 2796 237162 2848
rect 239306 2796 239312 2848
rect 239364 2836 239370 2848
rect 240594 2836 240600 2848
rect 239364 2808 240600 2836
rect 239364 2796 239370 2808
rect 240594 2796 240600 2808
rect 240652 2796 240658 2848
rect 242894 2796 242900 2848
rect 242952 2836 242958 2848
rect 244090 2836 244096 2848
rect 242952 2808 244096 2836
rect 242952 2796 242958 2808
rect 244090 2796 244096 2808
rect 244148 2796 244154 2848
rect 244182 2796 244188 2848
rect 244240 2836 244246 2848
rect 245286 2836 245292 2848
rect 244240 2808 245292 2836
rect 244240 2796 244246 2808
rect 245286 2796 245292 2808
rect 245344 2796 245350 2848
rect 247586 2796 247592 2848
rect 247644 2836 247650 2848
rect 248782 2836 248788 2848
rect 247644 2808 248788 2836
rect 247644 2796 247650 2808
rect 248782 2796 248788 2808
rect 248840 2796 248846 2848
rect 249978 2796 249984 2848
rect 250036 2836 250042 2848
rect 251082 2836 251088 2848
rect 250036 2808 251088 2836
rect 250036 2796 250042 2808
rect 251082 2796 251088 2808
rect 251140 2796 251146 2848
rect 253474 2796 253480 2848
rect 253532 2836 253538 2848
rect 254578 2836 254584 2848
rect 253532 2808 254584 2836
rect 253532 2796 253538 2808
rect 254578 2796 254584 2808
rect 254636 2796 254642 2848
rect 254670 2796 254676 2848
rect 254728 2836 254734 2848
rect 255774 2836 255780 2848
rect 254728 2808 255780 2836
rect 254728 2796 254734 2808
rect 255774 2796 255780 2808
rect 255832 2796 255838 2848
rect 255866 2796 255872 2848
rect 255924 2836 255930 2848
rect 256970 2836 256976 2848
rect 255924 2808 256976 2836
rect 255924 2796 255930 2808
rect 256970 2796 256976 2808
rect 257028 2796 257034 2848
rect 257062 2796 257068 2848
rect 257120 2836 257126 2848
rect 258074 2836 258080 2848
rect 257120 2808 258080 2836
rect 257120 2796 257126 2808
rect 258074 2796 258080 2808
rect 258132 2796 258138 2848
rect 259454 2796 259460 2848
rect 259512 2836 259518 2848
rect 260466 2836 260472 2848
rect 259512 2808 260472 2836
rect 259512 2796 259518 2808
rect 260466 2796 260472 2808
rect 260524 2796 260530 2848
rect 260650 2796 260656 2848
rect 260708 2836 260714 2848
rect 261570 2836 261576 2848
rect 260708 2808 261576 2836
rect 260708 2796 260714 2808
rect 261570 2796 261576 2808
rect 261628 2796 261634 2848
rect 261754 2796 261760 2848
rect 261812 2836 261818 2848
rect 262766 2836 262772 2848
rect 261812 2808 262772 2836
rect 261812 2796 261818 2808
rect 262766 2796 262772 2808
rect 262824 2796 262830 2848
rect 262950 2796 262956 2848
rect 263008 2836 263014 2848
rect 263962 2836 263968 2848
rect 263008 2808 263968 2836
rect 263008 2796 263014 2808
rect 263962 2796 263968 2808
rect 264020 2796 264026 2848
rect 264146 2796 264152 2848
rect 264204 2836 264210 2848
rect 265066 2836 265072 2848
rect 264204 2808 265072 2836
rect 264204 2796 264210 2808
rect 265066 2796 265072 2808
rect 265124 2796 265130 2848
rect 266538 2796 266544 2848
rect 266596 2836 266602 2848
rect 267458 2836 267464 2848
rect 266596 2808 267464 2836
rect 266596 2796 266602 2808
rect 267458 2796 267464 2808
rect 267516 2796 267522 2848
rect 267734 2796 267740 2848
rect 267792 2836 267798 2848
rect 268654 2836 268660 2848
rect 267792 2808 268660 2836
rect 267792 2796 267798 2808
rect 268654 2796 268660 2808
rect 268712 2796 268718 2848
rect 268838 2796 268844 2848
rect 268896 2836 268902 2848
rect 269758 2836 269764 2848
rect 268896 2808 269764 2836
rect 268896 2796 268902 2808
rect 269758 2796 269764 2808
rect 269816 2796 269822 2848
rect 270034 2796 270040 2848
rect 270092 2836 270098 2848
rect 270954 2836 270960 2848
rect 270092 2808 270960 2836
rect 270092 2796 270098 2808
rect 270954 2796 270960 2808
rect 271012 2796 271018 2848
rect 271230 2796 271236 2848
rect 271288 2836 271294 2848
rect 272150 2836 272156 2848
rect 271288 2808 272156 2836
rect 271288 2796 271294 2808
rect 272150 2796 272156 2808
rect 272208 2796 272214 2848
rect 272426 2796 272432 2848
rect 272484 2836 272490 2848
rect 273254 2836 273260 2848
rect 272484 2808 273260 2836
rect 272484 2796 272490 2808
rect 273254 2796 273260 2808
rect 273312 2796 273318 2848
rect 273622 2796 273628 2848
rect 273680 2836 273686 2848
rect 274450 2836 274456 2848
rect 273680 2808 274456 2836
rect 273680 2796 273686 2808
rect 274450 2796 274456 2808
rect 274508 2796 274514 2848
rect 274818 2796 274824 2848
rect 274876 2836 274882 2848
rect 275646 2836 275652 2848
rect 274876 2808 275652 2836
rect 274876 2796 274882 2808
rect 275646 2796 275652 2808
rect 275704 2796 275710 2848
rect 277118 2796 277124 2848
rect 277176 2836 277182 2848
rect 277946 2836 277952 2848
rect 277176 2808 277952 2836
rect 277176 2796 277182 2808
rect 277946 2796 277952 2808
rect 278004 2796 278010 2848
rect 278314 2796 278320 2848
rect 278372 2836 278378 2848
rect 279142 2836 279148 2848
rect 278372 2808 279148 2836
rect 278372 2796 278378 2808
rect 279142 2796 279148 2808
rect 279200 2796 279206 2848
rect 279510 2796 279516 2848
rect 279568 2836 279574 2848
rect 280246 2836 280252 2848
rect 279568 2808 280252 2836
rect 279568 2796 279574 2808
rect 280246 2796 280252 2808
rect 280304 2796 280310 2848
rect 280706 2796 280712 2848
rect 280764 2836 280770 2848
rect 281442 2836 281448 2848
rect 280764 2808 281448 2836
rect 280764 2796 280770 2808
rect 281442 2796 281448 2808
rect 281500 2796 281506 2848
rect 281902 2796 281908 2848
rect 281960 2836 281966 2848
rect 282638 2836 282644 2848
rect 281960 2808 282644 2836
rect 281960 2796 281966 2808
rect 282638 2796 282644 2808
rect 282696 2796 282702 2848
rect 284294 2796 284300 2848
rect 284352 2836 284358 2848
rect 284938 2836 284944 2848
rect 284352 2808 284944 2836
rect 284352 2796 284358 2808
rect 284938 2796 284944 2808
rect 284996 2796 285002 2848
rect 285398 2796 285404 2848
rect 285456 2836 285462 2848
rect 286134 2836 286140 2848
rect 285456 2808 286140 2836
rect 285456 2796 285462 2808
rect 286134 2796 286140 2808
rect 286192 2796 286198 2848
rect 286594 2796 286600 2848
rect 286652 2836 286658 2848
rect 287238 2836 287244 2848
rect 286652 2808 287244 2836
rect 286652 2796 286658 2808
rect 287238 2796 287244 2808
rect 287296 2796 287302 2848
rect 287790 2796 287796 2848
rect 287848 2836 287854 2848
rect 288434 2836 288440 2848
rect 287848 2808 288440 2836
rect 287848 2796 287854 2808
rect 288434 2796 288440 2808
rect 288492 2796 288498 2848
rect 288986 2796 288992 2848
rect 289044 2836 289050 2848
rect 289630 2836 289636 2848
rect 289044 2808 289636 2836
rect 289044 2796 289050 2808
rect 289630 2796 289636 2808
rect 289688 2796 289694 2848
rect 291378 2796 291384 2848
rect 291436 2836 291442 2848
rect 291930 2836 291936 2848
rect 291436 2808 291936 2836
rect 291436 2796 291442 2808
rect 291930 2796 291936 2808
rect 291988 2796 291994 2848
rect 292574 2796 292580 2848
rect 292632 2836 292638 2848
rect 293126 2836 293132 2848
rect 292632 2808 293132 2836
rect 292632 2796 292638 2808
rect 293126 2796 293132 2808
rect 293184 2796 293190 2848
rect 293678 2796 293684 2848
rect 293736 2836 293742 2848
rect 294322 2836 294328 2848
rect 293736 2808 294328 2836
rect 293736 2796 293742 2808
rect 294322 2796 294328 2808
rect 294380 2796 294386 2848
rect 294874 2796 294880 2848
rect 294932 2836 294938 2848
rect 295426 2836 295432 2848
rect 294932 2808 295432 2836
rect 294932 2796 294938 2808
rect 295426 2796 295432 2808
rect 295484 2796 295490 2848
rect 296070 2796 296076 2848
rect 296128 2836 296134 2848
rect 296622 2836 296628 2848
rect 296128 2808 296628 2836
rect 296128 2796 296134 2808
rect 296622 2796 296628 2808
rect 296680 2796 296686 2848
rect 298462 2796 298468 2848
rect 298520 2836 298526 2848
rect 298922 2836 298928 2848
rect 298520 2808 298928 2836
rect 298520 2796 298526 2808
rect 298922 2796 298928 2808
rect 298980 2796 298986 2848
rect 299658 2796 299664 2848
rect 299716 2836 299722 2848
rect 300118 2836 300124 2848
rect 299716 2808 300124 2836
rect 299716 2796 299722 2808
rect 300118 2796 300124 2808
rect 300176 2796 300182 2848
rect 300762 2796 300768 2848
rect 300820 2836 300826 2848
rect 301314 2836 301320 2848
rect 300820 2808 301320 2836
rect 300820 2796 300826 2808
rect 301314 2796 301320 2808
rect 301372 2796 301378 2848
rect 301958 2796 301964 2848
rect 302016 2836 302022 2848
rect 302418 2836 302424 2848
rect 302016 2808 302424 2836
rect 302016 2796 302022 2808
rect 302418 2796 302424 2808
rect 302476 2796 302482 2848
rect 303154 2796 303160 2848
rect 303212 2836 303218 2848
rect 303614 2836 303620 2848
rect 303212 2808 303620 2836
rect 303212 2796 303218 2808
rect 303614 2796 303620 2808
rect 303672 2796 303678 2848
rect 368934 2796 368940 2848
rect 368992 2836 368998 2848
rect 369394 2836 369400 2848
rect 368992 2808 369400 2836
rect 368992 2796 368998 2808
rect 369394 2796 369400 2808
rect 369452 2796 369458 2848
rect 370130 2796 370136 2848
rect 370188 2836 370194 2848
rect 370590 2836 370596 2848
rect 370188 2808 370596 2836
rect 370188 2796 370194 2808
rect 370590 2796 370596 2808
rect 370648 2796 370654 2848
rect 375926 2796 375932 2848
rect 375984 2836 375990 2848
rect 376478 2836 376484 2848
rect 375984 2808 376484 2836
rect 375984 2796 375990 2808
rect 376478 2796 376484 2808
rect 376536 2796 376542 2848
rect 377122 2796 377128 2848
rect 377180 2836 377186 2848
rect 377674 2836 377680 2848
rect 377180 2808 377680 2836
rect 377180 2796 377186 2808
rect 377674 2796 377680 2808
rect 377732 2796 377738 2848
rect 382918 2796 382924 2848
rect 382976 2836 382982 2848
rect 383562 2836 383568 2848
rect 382976 2808 383568 2836
rect 382976 2796 382982 2808
rect 383562 2796 383568 2808
rect 383620 2796 383626 2848
rect 384114 2796 384120 2848
rect 384172 2836 384178 2848
rect 384758 2836 384764 2848
rect 384172 2808 384764 2836
rect 384172 2796 384178 2808
rect 384758 2796 384764 2808
rect 384816 2796 384822 2848
rect 386414 2796 386420 2848
rect 386472 2836 386478 2848
rect 387150 2836 387156 2848
rect 386472 2808 387156 2836
rect 386472 2796 386478 2808
rect 387150 2796 387156 2808
rect 387208 2796 387214 2848
rect 391106 2796 391112 2848
rect 391164 2836 391170 2848
rect 391842 2836 391848 2848
rect 391164 2808 391848 2836
rect 391164 2796 391170 2808
rect 391842 2796 391848 2808
rect 391900 2796 391906 2848
rect 393406 2796 393412 2848
rect 393464 2836 393470 2848
rect 394234 2836 394240 2848
rect 393464 2808 394240 2836
rect 393464 2796 393470 2808
rect 394234 2796 394240 2808
rect 394292 2796 394298 2848
rect 400490 2796 400496 2848
rect 400548 2836 400554 2848
rect 401318 2836 401324 2848
rect 400548 2808 401324 2836
rect 400548 2796 400554 2808
rect 401318 2796 401324 2808
rect 401376 2796 401382 2848
rect 401594 2796 401600 2848
rect 401652 2836 401658 2848
rect 402514 2836 402520 2848
rect 401652 2808 402520 2836
rect 401652 2796 401658 2808
rect 402514 2796 402520 2808
rect 402572 2796 402578 2848
rect 407482 2796 407488 2848
rect 407540 2836 407546 2848
rect 408402 2836 408408 2848
rect 407540 2808 408408 2836
rect 407540 2796 407546 2808
rect 408402 2796 408408 2808
rect 408460 2796 408466 2848
rect 408586 2796 408592 2848
rect 408644 2836 408650 2848
rect 409598 2836 409604 2848
rect 408644 2808 409604 2836
rect 408644 2796 408650 2808
rect 409598 2796 409604 2808
rect 409656 2796 409662 2848
rect 415578 2796 415584 2848
rect 415636 2836 415642 2848
rect 416682 2836 416688 2848
rect 415636 2808 416688 2836
rect 415636 2796 415642 2808
rect 416682 2796 416688 2808
rect 416740 2796 416746 2848
rect 431954 2796 431960 2848
rect 432012 2836 432018 2848
rect 433242 2836 433248 2848
rect 432012 2808 433248 2836
rect 432012 2796 432018 2808
rect 433242 2796 433248 2808
rect 433300 2796 433306 2848
rect 472250 2836 472256 2848
rect 470566 2808 472256 2836
rect 9582 2768 9588 2780
rect 6886 2740 9588 2768
rect 9582 2728 9588 2740
rect 9640 2728 9646 2780
rect 470410 2728 470416 2780
rect 470468 2768 470474 2780
rect 470566 2768 470594 2808
rect 472250 2796 472256 2808
rect 472308 2796 472314 2848
rect 480530 2836 480536 2848
rect 480226 2808 480536 2836
rect 470468 2740 470594 2768
rect 470468 2728 470474 2740
rect 478598 2728 478604 2780
rect 478656 2768 478662 2780
rect 480226 2768 480254 2808
rect 480530 2796 480536 2808
rect 480588 2796 480594 2848
rect 487614 2836 487620 2848
rect 487080 2808 487620 2836
rect 478656 2740 480254 2768
rect 478656 2728 478662 2740
rect 485590 2728 485596 2780
rect 485648 2768 485654 2780
rect 487080 2768 487108 2808
rect 487614 2796 487620 2808
rect 487672 2796 487678 2848
rect 492674 2796 492680 2848
rect 492732 2836 492738 2848
rect 494698 2836 494704 2848
rect 492732 2808 494704 2836
rect 492732 2796 492738 2808
rect 494698 2796 494704 2808
rect 494756 2796 494762 2848
rect 495894 2836 495900 2848
rect 495360 2808 495900 2836
rect 485648 2740 487108 2768
rect 485648 2728 485654 2740
rect 493778 2728 493784 2780
rect 493836 2768 493842 2780
rect 495360 2768 495388 2808
rect 495894 2796 495900 2808
rect 495952 2796 495958 2848
rect 502978 2836 502984 2848
rect 502260 2808 502984 2836
rect 493836 2740 495388 2768
rect 493836 2728 493842 2740
rect 500770 2728 500776 2780
rect 500828 2768 500834 2780
rect 502260 2768 502288 2808
rect 502978 2796 502984 2808
rect 503036 2796 503042 2848
rect 505370 2836 505376 2848
rect 505020 2808 505376 2836
rect 500828 2740 502288 2768
rect 500828 2728 500834 2740
rect 503162 2728 503168 2780
rect 503220 2768 503226 2780
rect 505020 2768 505048 2808
rect 505370 2796 505376 2808
rect 505428 2796 505434 2848
rect 507854 2796 507860 2848
rect 507912 2836 507918 2848
rect 510062 2836 510068 2848
rect 507912 2808 510068 2836
rect 507912 2796 507918 2808
rect 510062 2796 510068 2808
rect 510120 2796 510126 2848
rect 512454 2836 512460 2848
rect 511920 2808 512460 2836
rect 503220 2740 505048 2768
rect 503220 2728 503226 2740
rect 510154 2728 510160 2780
rect 510212 2768 510218 2780
rect 511920 2768 511948 2808
rect 512454 2796 512460 2808
rect 512512 2796 512518 2848
rect 518342 2836 518348 2848
rect 517072 2808 518348 2836
rect 510212 2740 511948 2768
rect 510212 2728 510218 2740
rect 515950 2728 515956 2780
rect 516008 2768 516014 2780
rect 517072 2768 517100 2808
rect 518342 2796 518348 2808
rect 518400 2796 518406 2848
rect 519538 2836 519544 2848
rect 518866 2808 519544 2836
rect 516008 2740 517100 2768
rect 516008 2728 516014 2740
rect 517146 2728 517152 2780
rect 517204 2768 517210 2780
rect 518866 2768 518894 2808
rect 519538 2796 519544 2808
rect 519596 2796 519602 2848
rect 521838 2836 521844 2848
rect 521580 2808 521844 2836
rect 517204 2740 518894 2768
rect 517204 2728 517210 2740
rect 519446 2728 519452 2780
rect 519504 2768 519510 2780
rect 521580 2768 521608 2808
rect 521838 2796 521844 2808
rect 521896 2796 521902 2848
rect 523034 2796 523040 2848
rect 523092 2836 523098 2848
rect 525426 2836 525432 2848
rect 523092 2808 525432 2836
rect 523092 2796 523098 2808
rect 525426 2796 525432 2808
rect 525484 2796 525490 2848
rect 526622 2836 526628 2848
rect 525720 2808 526628 2836
rect 519504 2740 521608 2768
rect 519504 2728 519510 2740
rect 524138 2728 524144 2780
rect 524196 2768 524202 2780
rect 525720 2768 525748 2808
rect 526622 2796 526628 2808
rect 526680 2796 526686 2848
rect 527818 2836 527824 2848
rect 527008 2808 527824 2836
rect 524196 2740 525748 2768
rect 524196 2728 524202 2740
rect 525242 2660 525248 2712
rect 525300 2700 525306 2712
rect 527008 2700 527036 2808
rect 527818 2796 527824 2808
rect 527876 2796 527882 2848
rect 533706 2836 533712 2848
rect 532620 2808 533712 2836
rect 531130 2728 531136 2780
rect 531188 2768 531194 2780
rect 532620 2768 532648 2808
rect 533706 2796 533712 2808
rect 533764 2796 533770 2848
rect 534902 2836 534908 2848
rect 534000 2808 534908 2836
rect 531188 2740 532648 2768
rect 531188 2728 531194 2740
rect 525300 2672 527036 2700
rect 525300 2660 525306 2672
rect 532326 2660 532332 2712
rect 532384 2700 532390 2712
rect 534000 2700 534028 2808
rect 534902 2796 534908 2808
rect 534960 2796 534966 2848
rect 537202 2836 537208 2848
rect 536760 2808 537208 2836
rect 534626 2728 534632 2780
rect 534684 2768 534690 2780
rect 536760 2768 536788 2808
rect 537202 2796 537208 2808
rect 537260 2796 537266 2848
rect 538214 2796 538220 2848
rect 538272 2836 538278 2848
rect 540790 2836 540796 2848
rect 538272 2808 540796 2836
rect 538272 2796 538278 2808
rect 540790 2796 540796 2808
rect 540848 2796 540854 2848
rect 541986 2836 541992 2848
rect 540900 2808 541992 2836
rect 534684 2740 536788 2768
rect 534684 2728 534690 2740
rect 539318 2728 539324 2780
rect 539376 2768 539382 2780
rect 540900 2768 540928 2808
rect 541986 2796 541992 2808
rect 542044 2796 542050 2848
rect 544378 2836 544384 2848
rect 542740 2808 544384 2836
rect 539376 2740 540928 2768
rect 539376 2728 539382 2740
rect 541618 2728 541624 2780
rect 541676 2768 541682 2780
rect 542740 2768 542768 2808
rect 544378 2796 544384 2808
rect 544436 2796 544442 2848
rect 545482 2836 545488 2848
rect 545040 2808 545488 2836
rect 541676 2740 542768 2768
rect 541676 2728 541682 2740
rect 542814 2728 542820 2780
rect 542872 2768 542878 2780
rect 545040 2768 545068 2808
rect 545482 2796 545488 2808
rect 545540 2796 545546 2848
rect 549070 2836 549076 2848
rect 547846 2808 549076 2836
rect 542872 2740 545068 2768
rect 542872 2728 542878 2740
rect 546310 2728 546316 2780
rect 546368 2768 546374 2780
rect 547846 2768 547874 2808
rect 549070 2796 549076 2808
rect 549128 2796 549134 2848
rect 551462 2836 551468 2848
rect 550560 2808 551468 2836
rect 546368 2740 547874 2768
rect 546368 2728 546374 2740
rect 548610 2728 548616 2780
rect 548668 2768 548674 2780
rect 550560 2768 550588 2808
rect 551462 2796 551468 2808
rect 551520 2796 551526 2848
rect 552658 2836 552664 2848
rect 551940 2808 552664 2836
rect 548668 2740 550588 2768
rect 548668 2728 548674 2740
rect 532384 2672 534028 2700
rect 532384 2660 532390 2672
rect 549806 2660 549812 2712
rect 549864 2700 549870 2712
rect 551940 2700 551968 2808
rect 552658 2796 552664 2808
rect 552716 2796 552722 2848
rect 554958 2836 554964 2848
rect 554700 2808 554964 2836
rect 552106 2728 552112 2780
rect 552164 2768 552170 2780
rect 554700 2768 554728 2808
rect 554958 2796 554964 2808
rect 555016 2796 555022 2848
rect 557350 2836 557356 2848
rect 555528 2808 557356 2836
rect 552164 2740 554728 2768
rect 552164 2728 552170 2740
rect 549864 2672 551968 2700
rect 549864 2660 549870 2672
rect 554498 2660 554504 2712
rect 554556 2700 554562 2712
rect 555528 2700 555556 2808
rect 557350 2796 557356 2808
rect 557408 2796 557414 2848
rect 558546 2836 558552 2848
rect 557506 2808 558552 2836
rect 555602 2728 555608 2780
rect 555660 2768 555666 2780
rect 557506 2768 557534 2808
rect 558546 2796 558552 2808
rect 558604 2796 558610 2848
rect 560846 2836 560852 2848
rect 560220 2808 560852 2836
rect 555660 2740 557534 2768
rect 555660 2728 555666 2740
rect 557994 2728 558000 2780
rect 558052 2768 558058 2780
rect 560220 2768 560248 2808
rect 560846 2796 560852 2808
rect 560904 2796 560910 2848
rect 563238 2836 563244 2848
rect 562980 2808 563244 2836
rect 558052 2740 560248 2768
rect 558052 2728 558058 2740
rect 560294 2728 560300 2780
rect 560352 2768 560358 2780
rect 562980 2768 563008 2808
rect 563238 2796 563244 2808
rect 563296 2796 563302 2848
rect 565630 2836 565636 2848
rect 564360 2808 565636 2836
rect 560352 2740 563008 2768
rect 560352 2728 560358 2740
rect 554556 2672 555556 2700
rect 554556 2660 554562 2672
rect 562594 2660 562600 2712
rect 562652 2700 562658 2712
rect 564360 2700 564388 2808
rect 565630 2796 565636 2808
rect 565688 2796 565694 2848
rect 566826 2836 566832 2848
rect 565740 2808 566832 2836
rect 565740 2768 565768 2808
rect 566826 2796 566832 2808
rect 566884 2796 566890 2848
rect 569126 2836 569132 2848
rect 567166 2808 569132 2836
rect 562652 2672 564388 2700
rect 565648 2740 565768 2768
rect 562652 2660 562658 2672
rect 563790 2592 563796 2644
rect 563848 2632 563854 2644
rect 565648 2632 565676 2740
rect 566090 2728 566096 2780
rect 566148 2768 566154 2780
rect 567166 2768 567194 2808
rect 569126 2796 569132 2808
rect 569184 2796 569190 2848
rect 570322 2836 570328 2848
rect 569880 2808 570328 2836
rect 566148 2740 567194 2768
rect 566148 2728 566154 2740
rect 567286 2728 567292 2780
rect 567344 2768 567350 2780
rect 569880 2768 569908 2808
rect 570322 2796 570328 2808
rect 570380 2796 570386 2848
rect 572714 2836 572720 2848
rect 571168 2808 572720 2836
rect 567344 2740 569908 2768
rect 567344 2728 567350 2740
rect 569586 2660 569592 2712
rect 569644 2700 569650 2712
rect 571168 2700 571196 2808
rect 572714 2796 572720 2808
rect 572772 2796 572778 2848
rect 575106 2836 575112 2848
rect 574020 2808 575112 2836
rect 571978 2728 571984 2780
rect 572036 2768 572042 2780
rect 574020 2768 574048 2808
rect 575106 2796 575112 2808
rect 575164 2796 575170 2848
rect 577406 2836 577412 2848
rect 576826 2808 577412 2836
rect 572036 2740 574048 2768
rect 572036 2728 572042 2740
rect 574278 2728 574284 2780
rect 574336 2768 574342 2780
rect 576826 2768 576854 2808
rect 577406 2796 577412 2808
rect 577464 2796 577470 2848
rect 582190 2836 582196 2848
rect 579540 2808 582196 2836
rect 574336 2740 576854 2768
rect 574336 2728 574342 2740
rect 577774 2728 577780 2780
rect 577832 2768 577838 2780
rect 579540 2768 579568 2808
rect 582190 2796 582196 2808
rect 582248 2796 582254 2848
rect 577832 2740 579568 2768
rect 577832 2728 577838 2740
rect 569644 2672 571196 2700
rect 569644 2660 569650 2672
rect 563848 2604 565676 2632
rect 563848 2592 563854 2604
rect 424962 2524 424968 2576
rect 425020 2564 425026 2576
rect 426066 2564 426072 2576
rect 425020 2536 426072 2564
rect 425020 2524 425026 2536
rect 426066 2524 426072 2536
rect 426124 2524 426130 2576
rect 428458 2456 428464 2508
rect 428516 2496 428522 2508
rect 429562 2496 429568 2508
rect 428516 2468 429568 2496
rect 428516 2456 428522 2468
rect 429562 2456 429568 2468
rect 429620 2456 429626 2508
rect 423766 2388 423772 2440
rect 423824 2428 423830 2440
rect 424962 2428 424968 2440
rect 423824 2400 424968 2428
rect 423824 2388 423830 2400
rect 424962 2388 424968 2400
rect 425020 2388 425026 2440
rect 427262 2320 427268 2372
rect 427320 2360 427326 2372
rect 428458 2360 428464 2372
rect 427320 2332 428464 2360
rect 427320 2320 427326 2332
rect 428458 2320 428464 2332
rect 428516 2320 428522 2372
rect 511258 2320 511264 2372
rect 511316 2360 511322 2372
rect 513558 2360 513564 2372
rect 511316 2332 513564 2360
rect 511316 2320 511322 2332
rect 513558 2320 513564 2332
rect 513616 2320 513622 2372
rect 514754 2320 514760 2372
rect 514812 2360 514818 2372
rect 517146 2360 517152 2372
rect 514812 2332 517152 2360
rect 514812 2320 514818 2332
rect 517146 2320 517152 2332
rect 517204 2320 517210 2372
rect 304350 2252 304356 2304
rect 304408 2292 304414 2304
rect 304810 2292 304816 2304
rect 304408 2264 304816 2292
rect 304408 2252 304414 2264
rect 304810 2252 304816 2264
rect 304868 2252 304874 2304
rect 380618 2252 380624 2304
rect 380676 2292 380682 2304
rect 381170 2292 381176 2304
rect 380676 2264 381176 2292
rect 380676 2252 380682 2264
rect 381170 2252 381176 2264
rect 381228 2252 381234 2304
rect 398098 2252 398104 2304
rect 398156 2292 398162 2304
rect 398926 2292 398932 2304
rect 398156 2264 398932 2292
rect 398156 2252 398162 2264
rect 398926 2252 398932 2264
rect 398984 2252 398990 2304
rect 402790 2252 402796 2304
rect 402848 2292 402854 2304
rect 403618 2292 403624 2304
rect 402848 2264 403624 2292
rect 402848 2252 402854 2264
rect 403618 2252 403624 2264
rect 403676 2252 403682 2304
rect 409782 2252 409788 2304
rect 409840 2292 409846 2304
rect 410794 2292 410800 2304
rect 409840 2264 410800 2292
rect 409840 2252 409846 2264
rect 410794 2252 410800 2264
rect 410852 2252 410858 2304
rect 412082 2252 412088 2304
rect 412140 2292 412146 2304
rect 413094 2292 413100 2304
rect 412140 2264 413100 2292
rect 412140 2252 412146 2264
rect 413094 2252 413100 2264
rect 413152 2252 413158 2304
rect 414474 2252 414480 2304
rect 414532 2292 414538 2304
rect 415486 2292 415492 2304
rect 414532 2264 415492 2292
rect 414532 2252 414538 2264
rect 415486 2252 415492 2264
rect 415544 2252 415550 2304
rect 422570 2252 422576 2304
rect 422628 2292 422634 2304
rect 423766 2292 423772 2304
rect 422628 2264 423772 2292
rect 422628 2252 422634 2264
rect 423766 2252 423772 2264
rect 423824 2252 423830 2304
rect 429654 2252 429660 2304
rect 429712 2292 429718 2304
rect 430850 2292 430856 2304
rect 429712 2264 430856 2292
rect 429712 2252 429718 2264
rect 430850 2252 430856 2264
rect 430908 2252 430914 2304
rect 435450 2252 435456 2304
rect 435508 2292 435514 2304
rect 436738 2292 436744 2304
rect 435508 2264 436744 2292
rect 435508 2252 435514 2264
rect 436738 2252 436744 2264
rect 436796 2252 436802 2304
rect 438946 2252 438952 2304
rect 439004 2292 439010 2304
rect 440326 2292 440332 2304
rect 439004 2264 440332 2292
rect 439004 2252 439010 2264
rect 440326 2252 440332 2264
rect 440384 2252 440390 2304
rect 441246 2252 441252 2304
rect 441304 2292 441310 2304
rect 442626 2292 442632 2304
rect 441304 2264 442632 2292
rect 441304 2252 441310 2264
rect 442626 2252 442632 2264
rect 442684 2252 442690 2304
rect 450630 2252 450636 2304
rect 450688 2292 450694 2304
rect 452102 2292 452108 2304
rect 450688 2264 452108 2292
rect 450688 2252 450694 2264
rect 452102 2252 452108 2264
rect 452160 2252 452166 2304
rect 452930 2252 452936 2304
rect 452988 2292 452994 2304
rect 454494 2292 454500 2304
rect 452988 2264 454500 2292
rect 452988 2252 452994 2264
rect 454494 2252 454500 2264
rect 454552 2252 454558 2304
rect 486786 2252 486792 2304
rect 486844 2292 486850 2304
rect 488810 2292 488816 2304
rect 486844 2264 488816 2292
rect 486844 2252 486850 2264
rect 488810 2252 488816 2264
rect 488868 2252 488874 2304
rect 494974 2252 494980 2304
rect 495032 2292 495038 2304
rect 497090 2292 497096 2304
rect 495032 2264 497096 2292
rect 495032 2252 495038 2264
rect 497090 2252 497096 2264
rect 497148 2252 497154 2304
rect 497274 2252 497280 2304
rect 497332 2292 497338 2304
rect 499390 2292 499396 2304
rect 497332 2264 499396 2292
rect 497332 2252 497338 2264
rect 499390 2252 499396 2264
rect 499448 2252 499454 2304
rect 520642 2252 520648 2304
rect 520700 2292 520706 2304
rect 523034 2292 523040 2304
rect 520700 2264 523040 2292
rect 520700 2252 520706 2264
rect 523034 2252 523040 2264
rect 523092 2252 523098 2304
rect 526438 2252 526444 2304
rect 526496 2292 526502 2304
rect 529014 2292 529020 2304
rect 526496 2264 529020 2292
rect 526496 2252 526502 2264
rect 529014 2252 529020 2264
rect 529072 2252 529078 2304
rect 535822 2252 535828 2304
rect 535880 2292 535886 2304
rect 535880 2264 536880 2292
rect 535880 2252 535886 2264
rect 566 2184 572 2236
rect 624 2224 630 2236
rect 4982 2224 4988 2236
rect 624 2196 4988 2224
rect 624 2184 630 2196
rect 4982 2184 4988 2196
rect 5040 2184 5046 2236
rect 251174 2184 251180 2236
rect 251232 2224 251238 2236
rect 252278 2224 252284 2236
rect 251232 2196 252284 2224
rect 251232 2184 251238 2196
rect 252278 2184 252284 2196
rect 252336 2184 252342 2236
rect 258258 2184 258264 2236
rect 258316 2224 258322 2236
rect 259270 2224 259276 2236
rect 258316 2196 259276 2224
rect 258316 2184 258322 2196
rect 259270 2184 259276 2196
rect 259328 2184 259334 2236
rect 290182 2184 290188 2236
rect 290240 2224 290246 2236
rect 290734 2224 290740 2236
rect 290240 2196 290740 2224
rect 290240 2184 290246 2196
rect 290734 2184 290740 2196
rect 290792 2184 290798 2236
rect 297266 2184 297272 2236
rect 297324 2224 297330 2236
rect 297818 2224 297824 2236
rect 297324 2196 297824 2224
rect 297324 2184 297330 2196
rect 297818 2184 297824 2196
rect 297876 2184 297882 2236
rect 367738 2184 367744 2236
rect 367796 2224 367802 2236
rect 368198 2224 368204 2236
rect 367796 2196 368204 2224
rect 367796 2184 367802 2196
rect 368198 2184 368204 2196
rect 368256 2184 368262 2236
rect 373626 2184 373632 2236
rect 373684 2224 373690 2236
rect 374086 2224 374092 2236
rect 373684 2196 374092 2224
rect 373684 2184 373690 2196
rect 374086 2184 374092 2196
rect 374144 2184 374150 2236
rect 374822 2184 374828 2236
rect 374880 2224 374886 2236
rect 375282 2224 375288 2236
rect 374880 2196 375288 2224
rect 374880 2184 374886 2196
rect 375282 2184 375288 2196
rect 375340 2184 375346 2236
rect 378318 2184 378324 2236
rect 378376 2224 378382 2236
rect 378870 2224 378876 2236
rect 378376 2196 378876 2224
rect 378376 2184 378382 2196
rect 378870 2184 378876 2196
rect 378928 2184 378934 2236
rect 379422 2184 379428 2236
rect 379480 2224 379486 2236
rect 379974 2224 379980 2236
rect 379480 2196 379980 2224
rect 379480 2184 379486 2196
rect 379974 2184 379980 2196
rect 380032 2184 380038 2236
rect 385310 2184 385316 2236
rect 385368 2224 385374 2236
rect 385954 2224 385960 2236
rect 385368 2196 385960 2224
rect 385368 2184 385374 2196
rect 385954 2184 385960 2196
rect 386012 2184 386018 2236
rect 387610 2184 387616 2236
rect 387668 2224 387674 2236
rect 388254 2224 388260 2236
rect 387668 2196 388260 2224
rect 387668 2184 387674 2196
rect 388254 2184 388260 2196
rect 388312 2184 388318 2236
rect 388806 2184 388812 2236
rect 388864 2224 388870 2236
rect 389450 2224 389456 2236
rect 388864 2196 389456 2224
rect 388864 2184 388870 2196
rect 389450 2184 389456 2196
rect 389508 2184 389514 2236
rect 389910 2184 389916 2236
rect 389968 2224 389974 2236
rect 390646 2224 390652 2236
rect 389968 2196 390652 2224
rect 389968 2184 389974 2196
rect 390646 2184 390652 2196
rect 390704 2184 390710 2236
rect 392302 2184 392308 2236
rect 392360 2224 392366 2236
rect 393038 2224 393044 2236
rect 392360 2196 393044 2224
rect 392360 2184 392366 2196
rect 393038 2184 393044 2196
rect 393096 2184 393102 2236
rect 394602 2184 394608 2236
rect 394660 2224 394666 2236
rect 395338 2224 395344 2236
rect 394660 2196 395344 2224
rect 394660 2184 394666 2196
rect 395338 2184 395344 2196
rect 395396 2184 395402 2236
rect 395798 2184 395804 2236
rect 395856 2224 395862 2236
rect 396534 2224 396540 2236
rect 395856 2196 396540 2224
rect 395856 2184 395862 2196
rect 396534 2184 396540 2196
rect 396592 2184 396598 2236
rect 399294 2184 399300 2236
rect 399352 2224 399358 2236
rect 400122 2224 400128 2236
rect 399352 2196 400128 2224
rect 399352 2184 399358 2196
rect 400122 2184 400128 2196
rect 400180 2184 400186 2236
rect 410978 2184 410984 2236
rect 411036 2224 411042 2236
rect 411898 2224 411904 2236
rect 411036 2196 411904 2224
rect 411036 2184 411042 2196
rect 411898 2184 411904 2196
rect 411956 2184 411962 2236
rect 417970 2184 417976 2236
rect 418028 2224 418034 2236
rect 418982 2224 418988 2236
rect 418028 2196 418988 2224
rect 418028 2184 418034 2196
rect 418982 2184 418988 2196
rect 419040 2184 419046 2236
rect 426158 2184 426164 2236
rect 426216 2224 426222 2236
rect 427262 2224 427268 2236
rect 426216 2196 427268 2224
rect 426216 2184 426222 2196
rect 427262 2184 427268 2196
rect 427320 2184 427326 2236
rect 437750 2184 437756 2236
rect 437808 2224 437814 2236
rect 439130 2224 439136 2236
rect 437808 2196 439136 2224
rect 437808 2184 437814 2196
rect 439130 2184 439136 2196
rect 439188 2184 439194 2236
rect 443638 2184 443644 2236
rect 443696 2224 443702 2236
rect 445018 2224 445024 2236
rect 443696 2196 445024 2224
rect 443696 2184 443702 2196
rect 445018 2184 445024 2196
rect 445076 2184 445082 2236
rect 451826 2184 451832 2236
rect 451884 2224 451890 2236
rect 453298 2224 453304 2236
rect 451884 2196 453304 2224
rect 451884 2184 451890 2196
rect 453298 2184 453304 2196
rect 453356 2184 453362 2236
rect 458818 2184 458824 2236
rect 458876 2224 458882 2236
rect 460382 2224 460388 2236
rect 458876 2196 460388 2224
rect 458876 2184 458882 2196
rect 460382 2184 460388 2196
rect 460440 2184 460446 2236
rect 463418 2184 463424 2236
rect 463476 2224 463482 2236
rect 465166 2224 465172 2236
rect 463476 2196 465172 2224
rect 463476 2184 463482 2196
rect 465166 2184 465172 2196
rect 465224 2184 465230 2236
rect 466914 2184 466920 2236
rect 466972 2224 466978 2236
rect 468662 2224 468668 2236
rect 466972 2196 468668 2224
rect 466972 2184 466978 2196
rect 468662 2184 468668 2196
rect 468720 2184 468726 2236
rect 471606 2184 471612 2236
rect 471664 2224 471670 2236
rect 473446 2224 473452 2236
rect 471664 2196 473452 2224
rect 471664 2184 471670 2196
rect 473446 2184 473452 2196
rect 473504 2184 473510 2236
rect 473906 2184 473912 2236
rect 473964 2224 473970 2236
rect 475746 2224 475752 2236
rect 473964 2196 475752 2224
rect 473964 2184 473970 2196
rect 475746 2184 475752 2196
rect 475804 2184 475810 2236
rect 476298 2184 476304 2236
rect 476356 2224 476362 2236
rect 478138 2224 478144 2236
rect 476356 2196 478144 2224
rect 476356 2184 476362 2196
rect 478138 2184 478144 2196
rect 478196 2184 478202 2236
rect 479794 2184 479800 2236
rect 479852 2224 479858 2236
rect 481726 2224 481732 2236
rect 479852 2196 481732 2224
rect 479852 2184 479858 2196
rect 481726 2184 481732 2196
rect 481784 2184 481790 2236
rect 483290 2184 483296 2236
rect 483348 2224 483354 2236
rect 485222 2224 485228 2236
rect 483348 2196 485228 2224
rect 483348 2184 483354 2196
rect 485222 2184 485228 2196
rect 485280 2184 485286 2236
rect 487982 2184 487988 2236
rect 488040 2224 488046 2236
rect 489914 2224 489920 2236
rect 488040 2196 489920 2224
rect 488040 2184 488046 2196
rect 489914 2184 489920 2196
rect 489972 2184 489978 2236
rect 496078 2184 496084 2236
rect 496136 2224 496142 2236
rect 498194 2224 498200 2236
rect 496136 2196 498200 2224
rect 496136 2184 496142 2196
rect 498194 2184 498200 2196
rect 498252 2184 498258 2236
rect 501966 2184 501972 2236
rect 502024 2224 502030 2236
rect 504174 2224 504180 2236
rect 502024 2196 504180 2224
rect 502024 2184 502030 2196
rect 504174 2184 504180 2196
rect 504232 2184 504238 2236
rect 504266 2184 504272 2236
rect 504324 2224 504330 2236
rect 506474 2224 506480 2236
rect 504324 2196 506480 2224
rect 504324 2184 504330 2196
rect 506474 2184 506480 2196
rect 506532 2184 506538 2236
rect 506658 2184 506664 2236
rect 506716 2224 506722 2236
rect 508866 2224 508872 2236
rect 506716 2196 508872 2224
rect 506716 2184 506722 2196
rect 508866 2184 508872 2196
rect 508924 2184 508930 2236
rect 508958 2184 508964 2236
rect 509016 2224 509022 2236
rect 511258 2224 511264 2236
rect 509016 2196 511264 2224
rect 509016 2184 509022 2196
rect 511258 2184 511264 2196
rect 511316 2184 511322 2236
rect 512546 2184 512552 2236
rect 512604 2224 512610 2236
rect 514754 2224 514760 2236
rect 512604 2196 514760 2224
rect 512604 2184 512610 2196
rect 514754 2184 514760 2196
rect 514812 2184 514818 2236
rect 518250 2184 518256 2236
rect 518308 2224 518314 2236
rect 520734 2224 520740 2236
rect 518308 2196 520740 2224
rect 518308 2184 518314 2196
rect 520734 2184 520740 2196
rect 520792 2184 520798 2236
rect 521746 2184 521752 2236
rect 521804 2224 521810 2236
rect 524230 2224 524236 2236
rect 521804 2196 524236 2224
rect 521804 2184 521810 2196
rect 524230 2184 524236 2196
rect 524288 2184 524294 2236
rect 527634 2184 527640 2236
rect 527692 2224 527698 2236
rect 530118 2224 530124 2236
rect 527692 2196 530124 2224
rect 527692 2184 527698 2196
rect 530118 2184 530124 2196
rect 530176 2184 530182 2236
rect 533430 2184 533436 2236
rect 533488 2224 533494 2236
rect 536098 2224 536104 2236
rect 533488 2196 536104 2224
rect 533488 2184 533494 2196
rect 536098 2184 536104 2196
rect 536156 2184 536162 2236
rect 536852 2224 536880 2264
rect 536926 2252 536932 2304
rect 536984 2292 536990 2304
rect 539594 2292 539600 2304
rect 536984 2264 539600 2292
rect 536984 2252 536990 2264
rect 539594 2252 539600 2264
rect 539652 2252 539658 2304
rect 545114 2252 545120 2304
rect 545172 2292 545178 2304
rect 547874 2292 547880 2304
rect 545172 2264 547880 2292
rect 545172 2252 545178 2264
rect 547874 2252 547880 2264
rect 547932 2252 547938 2304
rect 559098 2252 559104 2304
rect 559156 2292 559162 2304
rect 562042 2292 562048 2304
rect 559156 2264 562048 2292
rect 559156 2252 559162 2264
rect 562042 2252 562048 2264
rect 562100 2252 562106 2304
rect 538398 2224 538404 2236
rect 536852 2196 538404 2224
rect 538398 2184 538404 2196
rect 538456 2184 538462 2236
rect 543918 2184 543924 2236
rect 543976 2224 543982 2236
rect 546678 2224 546684 2236
rect 543976 2196 546684 2224
rect 543976 2184 543982 2196
rect 546678 2184 546684 2196
rect 546736 2184 546742 2236
rect 550910 2184 550916 2236
rect 550968 2224 550974 2236
rect 553762 2224 553768 2236
rect 550968 2196 553768 2224
rect 550968 2184 550974 2196
rect 553762 2184 553768 2196
rect 553820 2184 553826 2236
rect 556798 2184 556804 2236
rect 556856 2224 556862 2236
rect 559742 2224 559748 2236
rect 556856 2196 559748 2224
rect 556856 2184 556862 2196
rect 559742 2184 559748 2196
rect 559800 2184 559806 2236
rect 564986 2184 564992 2236
rect 565044 2224 565050 2236
rect 568022 2224 568028 2236
rect 565044 2196 568028 2224
rect 565044 2184 565050 2196
rect 568022 2184 568028 2196
rect 568080 2184 568086 2236
rect 575474 2184 575480 2236
rect 575532 2224 575538 2236
rect 578602 2224 578608 2236
rect 575532 2196 578608 2224
rect 575532 2184 575538 2196
rect 578602 2184 578608 2196
rect 578660 2184 578666 2236
rect 578970 2184 578976 2236
rect 579028 2224 579034 2236
rect 583386 2224 583392 2236
rect 579028 2196 583392 2224
rect 579028 2184 579034 2196
rect 583386 2184 583392 2196
rect 583444 2184 583450 2236
rect 372430 2116 372436 2168
rect 372488 2156 372494 2168
rect 372890 2156 372896 2168
rect 372488 2128 372896 2156
rect 372488 2116 372494 2128
rect 372890 2116 372896 2128
rect 372948 2116 372954 2168
rect 416774 2116 416780 2168
rect 416832 2156 416838 2168
rect 417878 2156 417884 2168
rect 416832 2128 417884 2156
rect 416832 2116 416838 2128
rect 417878 2116 417884 2128
rect 417936 2116 417942 2168
rect 420270 2116 420276 2168
rect 420328 2156 420334 2168
rect 421374 2156 421380 2168
rect 420328 2128 421380 2156
rect 420328 2116 420334 2128
rect 421374 2116 421380 2128
rect 421432 2116 421438 2168
rect 430758 2116 430764 2168
rect 430816 2156 430822 2168
rect 432046 2156 432052 2168
rect 430816 2128 432052 2156
rect 430816 2116 430822 2128
rect 432046 2116 432052 2128
rect 432104 2116 432110 2168
rect 434254 2116 434260 2168
rect 434312 2156 434318 2168
rect 435542 2156 435548 2168
rect 434312 2128 435548 2156
rect 434312 2116 434318 2128
rect 435542 2116 435548 2128
rect 435600 2116 435606 2168
rect 436646 2116 436652 2168
rect 436704 2156 436710 2168
rect 437934 2156 437940 2168
rect 436704 2128 437940 2156
rect 436704 2116 436710 2128
rect 437934 2116 437940 2128
rect 437992 2116 437998 2168
rect 444742 2116 444748 2168
rect 444800 2156 444806 2168
rect 446214 2156 446220 2168
rect 444800 2128 446220 2156
rect 444800 2116 444806 2128
rect 446214 2116 446220 2128
rect 446272 2116 446278 2168
rect 447134 2116 447140 2168
rect 447192 2156 447198 2168
rect 448606 2156 448612 2168
rect 447192 2128 448612 2156
rect 447192 2116 447198 2128
rect 448606 2116 448612 2128
rect 448664 2116 448670 2168
rect 454126 2116 454132 2168
rect 454184 2156 454190 2168
rect 455690 2156 455696 2168
rect 454184 2128 455696 2156
rect 454184 2116 454190 2128
rect 455690 2116 455696 2128
rect 455748 2116 455754 2168
rect 573082 2116 573088 2168
rect 573140 2156 573146 2168
rect 576302 2156 576308 2168
rect 573140 2128 576308 2156
rect 573140 2116 573146 2128
rect 576302 2116 576308 2128
rect 576360 2116 576366 2168
rect 406286 2048 406292 2100
rect 406344 2088 406350 2100
rect 407206 2088 407212 2100
rect 406344 2060 407212 2088
rect 406344 2048 406350 2060
rect 407206 2048 407212 2060
rect 407264 2048 407270 2100
rect 449434 2048 449440 2100
rect 449492 2088 449498 2100
rect 450906 2088 450912 2100
rect 449492 2060 450912 2088
rect 449492 2048 449498 2060
rect 450906 2048 450912 2060
rect 450964 2048 450970 2100
rect 455322 2048 455328 2100
rect 455380 2088 455386 2100
rect 456886 2088 456892 2100
rect 455380 2060 456892 2088
rect 455380 2048 455386 2060
rect 456886 2048 456892 2060
rect 456944 2048 456950 2100
rect 576578 2048 576584 2100
rect 576636 2088 576642 2100
rect 580994 2088 581000 2100
rect 576636 2060 581000 2088
rect 576636 2048 576642 2060
rect 580994 2048 581000 2060
rect 581052 2048 581058 2100
rect 265342 1980 265348 2032
rect 265400 2020 265406 2032
rect 266262 2020 266268 2032
rect 265400 1992 266268 2020
rect 265400 1980 265406 1992
rect 266262 1980 266268 1992
rect 266320 1980 266326 2032
rect 381814 1980 381820 2032
rect 381872 2020 381878 2032
rect 382366 2020 382372 2032
rect 381872 1992 382372 2020
rect 381872 1980 381878 1992
rect 382366 1980 382372 1992
rect 382424 1980 382430 2032
rect 440142 1980 440148 2032
rect 440200 2020 440206 2032
rect 441522 2020 441528 2032
rect 440200 1992 441528 2020
rect 440200 1980 440206 1992
rect 441522 1980 441528 1992
rect 441580 1980 441586 2032
rect 276014 1912 276020 1964
rect 276072 1952 276078 1964
rect 276750 1952 276756 1964
rect 276072 1924 276756 1952
rect 276072 1912 276078 1924
rect 276750 1912 276756 1924
rect 276808 1912 276814 1964
rect 442442 1912 442448 1964
rect 442500 1952 442506 1964
rect 443822 1952 443828 1964
rect 442500 1924 443828 1952
rect 442500 1912 442506 1924
rect 443822 1912 443828 1924
rect 443880 1912 443886 1964
rect 489086 1912 489092 1964
rect 489144 1952 489150 1964
rect 491110 1952 491116 1964
rect 489144 1924 491116 1952
rect 489144 1912 489150 1924
rect 491110 1912 491116 1924
rect 491168 1912 491174 1964
rect 513650 1912 513656 1964
rect 513708 1952 513714 1964
rect 515950 1952 515956 1964
rect 513708 1924 515956 1952
rect 513708 1912 513714 1924
rect 515950 1912 515956 1924
rect 516008 1912 516014 1964
rect 528830 1912 528836 1964
rect 528888 1952 528894 1964
rect 531314 1952 531320 1964
rect 528888 1924 531320 1952
rect 528888 1912 528894 1924
rect 531314 1912 531320 1924
rect 531372 1912 531378 1964
rect 419074 1844 419080 1896
rect 419132 1884 419138 1896
rect 420178 1884 420184 1896
rect 419132 1856 420184 1884
rect 419132 1844 419138 1856
rect 420178 1844 420184 1856
rect 420236 1844 420242 1896
rect 459922 1844 459928 1896
rect 459980 1884 459986 1896
rect 461578 1884 461584 1896
rect 459980 1856 461584 1884
rect 459980 1844 459986 1856
rect 461578 1844 461584 1856
rect 461636 1844 461642 1896
rect 396902 1776 396908 1828
rect 396960 1816 396966 1828
rect 397730 1816 397736 1828
rect 396960 1788 397736 1816
rect 396960 1776 396966 1788
rect 397730 1776 397736 1788
rect 397788 1776 397794 1828
rect 490282 1776 490288 1828
rect 490340 1816 490346 1828
rect 492306 1816 492312 1828
rect 490340 1788 492312 1816
rect 490340 1776 490346 1788
rect 492306 1776 492312 1788
rect 492364 1776 492370 1828
rect 498470 1776 498476 1828
rect 498528 1816 498534 1828
rect 500586 1816 500592 1828
rect 498528 1788 500592 1816
rect 498528 1776 498534 1788
rect 500586 1776 500592 1788
rect 500644 1776 500650 1828
rect 505462 1776 505468 1828
rect 505520 1816 505526 1828
rect 507670 1816 507676 1828
rect 505520 1788 507676 1816
rect 505520 1776 505526 1788
rect 507670 1776 507676 1788
rect 507728 1776 507734 1828
rect 529934 1776 529940 1828
rect 529992 1816 529998 1828
rect 532510 1816 532516 1828
rect 529992 1788 532516 1816
rect 529992 1776 529998 1788
rect 532510 1776 532516 1788
rect 532568 1776 532574 1828
rect 462314 1708 462320 1760
rect 462372 1748 462378 1760
rect 463970 1748 463976 1760
rect 462372 1720 463976 1748
rect 462372 1708 462378 1720
rect 463970 1708 463976 1720
rect 464028 1708 464034 1760
rect 482094 1708 482100 1760
rect 482152 1748 482158 1760
rect 484026 1748 484032 1760
rect 482152 1720 484032 1748
rect 482152 1708 482158 1720
rect 484026 1708 484032 1720
rect 484084 1708 484090 1760
rect 491478 1708 491484 1760
rect 491536 1748 491542 1760
rect 493502 1748 493508 1760
rect 491536 1720 493508 1748
rect 491536 1708 491542 1720
rect 493502 1708 493508 1720
rect 493560 1708 493566 1760
rect 499574 1708 499580 1760
rect 499632 1748 499638 1760
rect 501782 1748 501788 1760
rect 499632 1720 501788 1748
rect 499632 1708 499638 1720
rect 501782 1708 501788 1720
rect 501840 1708 501846 1760
rect 283098 1640 283104 1692
rect 283156 1680 283162 1692
rect 283742 1680 283748 1692
rect 283156 1652 283748 1680
rect 283156 1640 283162 1652
rect 283742 1640 283748 1652
rect 283800 1640 283806 1692
rect 421466 1640 421472 1692
rect 421524 1680 421530 1692
rect 422570 1680 422576 1692
rect 421524 1652 422576 1680
rect 421524 1640 421530 1652
rect 422570 1640 422576 1652
rect 422628 1640 422634 1692
rect 445938 1640 445944 1692
rect 445996 1680 446002 1692
rect 447410 1680 447416 1692
rect 445996 1652 447416 1680
rect 445996 1640 446002 1652
rect 447410 1640 447416 1652
rect 447468 1640 447474 1692
rect 448238 1640 448244 1692
rect 448296 1680 448302 1692
rect 449802 1680 449808 1692
rect 448296 1652 449808 1680
rect 448296 1640 448302 1652
rect 449802 1640 449808 1652
rect 449860 1640 449866 1692
rect 472802 1640 472808 1692
rect 472860 1680 472866 1692
rect 474550 1680 474556 1692
rect 472860 1652 474556 1680
rect 472860 1640 472866 1652
rect 474550 1640 474556 1652
rect 474608 1640 474614 1692
rect 475102 1640 475108 1692
rect 475160 1680 475166 1692
rect 476942 1680 476948 1692
rect 475160 1652 476948 1680
rect 475160 1640 475166 1652
rect 476942 1640 476948 1652
rect 477000 1640 477006 1692
rect 468110 1572 468116 1624
rect 468168 1612 468174 1624
rect 469858 1612 469864 1624
rect 468168 1584 469864 1612
rect 468168 1572 468174 1584
rect 469858 1572 469864 1584
rect 469916 1572 469922 1624
rect 480990 1572 480996 1624
rect 481048 1612 481054 1624
rect 482830 1612 482836 1624
rect 481048 1584 482836 1612
rect 481048 1572 481054 1584
rect 482830 1572 482836 1584
rect 482888 1572 482894 1624
rect 484486 1572 484492 1624
rect 484544 1612 484550 1624
rect 486418 1612 486424 1624
rect 484544 1584 486424 1612
rect 484544 1572 484550 1584
rect 486418 1572 486424 1584
rect 486476 1572 486482 1624
rect 405090 1504 405096 1556
rect 405148 1544 405154 1556
rect 406010 1544 406016 1556
rect 405148 1516 406016 1544
rect 405148 1504 405154 1516
rect 406010 1504 406016 1516
rect 406068 1504 406074 1556
rect 413278 1504 413284 1556
rect 413336 1544 413342 1556
rect 414290 1544 414296 1556
rect 413336 1516 414296 1544
rect 413336 1504 413342 1516
rect 414290 1504 414296 1516
rect 414348 1504 414354 1556
rect 433150 1504 433156 1556
rect 433208 1544 433214 1556
rect 434438 1544 434444 1556
rect 433208 1516 434444 1544
rect 433208 1504 433214 1516
rect 434438 1504 434444 1516
rect 434496 1504 434502 1556
rect 456426 1504 456432 1556
rect 456484 1544 456490 1556
rect 458082 1544 458088 1556
rect 456484 1516 458088 1544
rect 456484 1504 456490 1516
rect 458082 1504 458088 1516
rect 458140 1504 458146 1556
rect 465810 1504 465816 1556
rect 465868 1544 465874 1556
rect 467466 1544 467472 1556
rect 465868 1516 467472 1544
rect 465868 1504 465874 1516
rect 467466 1504 467472 1516
rect 467524 1504 467530 1556
rect 469306 1504 469312 1556
rect 469364 1544 469370 1556
rect 471054 1544 471060 1556
rect 469364 1516 471060 1544
rect 469364 1504 469370 1516
rect 471054 1504 471060 1516
rect 471112 1504 471118 1556
rect 477494 1504 477500 1556
rect 477552 1544 477558 1556
rect 479334 1544 479340 1556
rect 477552 1516 479340 1544
rect 477552 1504 477558 1516
rect 479334 1504 479340 1516
rect 479392 1504 479398 1556
rect 457622 1436 457628 1488
rect 457680 1476 457686 1488
rect 459186 1476 459192 1488
rect 457680 1448 459192 1476
rect 457680 1436 457686 1448
rect 459186 1436 459192 1448
rect 459244 1436 459250 1488
rect 461118 1436 461124 1488
rect 461176 1476 461182 1488
rect 462774 1476 462780 1488
rect 461176 1448 462780 1476
rect 461176 1436 461182 1448
rect 462774 1436 462780 1448
rect 462832 1436 462838 1488
rect 464614 1436 464620 1488
rect 464672 1476 464678 1488
rect 466270 1476 466276 1488
rect 464672 1448 466276 1476
rect 464672 1436 464678 1448
rect 466270 1436 466276 1448
rect 466328 1436 466334 1488
rect 403986 1368 403992 1420
rect 404044 1408 404050 1420
rect 404814 1408 404820 1420
rect 404044 1380 404820 1408
rect 404044 1368 404050 1380
rect 404814 1368 404820 1380
rect 404872 1368 404878 1420
<< via1 >>
rect 6920 703808 6972 703860
rect 581644 703808 581696 703860
rect 279332 703740 279384 703792
rect 356060 703740 356112 703792
rect 238944 703672 238996 703724
rect 316040 703672 316092 703724
rect 264152 703604 264204 703656
rect 364248 703604 364300 703656
rect 249064 703536 249116 703588
rect 410432 703536 410484 703588
rect 233884 703468 233936 703520
rect 430028 703468 430080 703520
rect 218796 703400 218848 703452
rect 581552 703400 581604 703452
rect 1492 703332 1544 703384
rect 370136 703332 370188 703384
rect 203616 703264 203668 703316
rect 582288 703264 582340 703316
rect 1676 703196 1728 703248
rect 385316 703196 385368 703248
rect 188528 703128 188580 703180
rect 582196 703128 582248 703180
rect 1768 703060 1820 703112
rect 400404 703060 400456 703112
rect 178408 702992 178460 703044
rect 173348 702924 173400 702976
rect 582104 702924 582156 702976
rect 1860 702856 1912 702908
rect 415584 702856 415636 702908
rect 158260 702788 158312 702840
rect 582012 702788 582064 702840
rect 2412 702720 2464 702772
rect 445852 702720 445904 702772
rect 127992 702652 128044 702704
rect 22008 702584 22060 702636
rect 581736 702584 581788 702636
rect 11888 702516 11940 702568
rect 270684 702448 270736 702500
rect 314660 702448 314712 702500
rect 57336 702312 57388 702364
rect 244004 702244 244056 702296
rect 320824 702244 320876 702296
rect 286968 702176 287020 702228
rect 410524 702176 410576 702228
rect 168288 702108 168340 702160
rect 336556 702108 336608 702160
rect 133052 702040 133104 702092
rect 329840 702040 329892 702092
rect 332600 702040 332652 702092
rect 380256 702040 380308 702092
rect 138020 701972 138072 702024
rect 342076 701972 342128 702024
rect 266360 701904 266412 701956
rect 481180 701904 481232 701956
rect 47216 701836 47268 701888
rect 144368 701836 144420 701888
rect 153200 701836 153252 701888
rect 4712 701768 4764 701820
rect 440792 701768 440844 701820
rect 32128 701700 32180 701752
rect 132684 701700 132736 701752
rect 148140 701700 148192 701752
rect 122932 701632 122984 701684
rect 572 701564 624 701616
rect 466000 701564 466052 701616
rect 4896 701496 4948 701548
rect 471060 701496 471112 701548
rect 117872 701428 117924 701480
rect 4804 701360 4856 701412
rect 486240 701360 486292 701412
rect 92664 701292 92716 701344
rect 581920 701292 581972 701344
rect 87604 701224 87656 701276
rect 4620 701156 4672 701208
rect 501328 701156 501380 701208
rect 571984 701156 572036 701208
rect 582564 701156 582616 701208
rect 77484 701088 77536 701140
rect 259184 701020 259236 701072
rect 303528 701020 303580 701072
rect 554780 701020 554832 701072
rect 577044 701020 577096 701072
rect 218980 700952 219032 701004
rect 319720 700952 319772 701004
rect 356060 700952 356112 701004
rect 364984 700952 365036 701004
rect 235172 700884 235224 700936
rect 309600 700884 309652 700936
rect 316040 700884 316092 700936
rect 527180 700884 527232 700936
rect 3792 700816 3844 700868
rect 218060 700816 218112 700868
rect 254124 700816 254176 700868
rect 462320 700816 462372 700868
rect 105452 700748 105504 700800
rect 339868 700748 339920 700800
rect 342076 700748 342128 700800
rect 580540 700748 580592 700800
rect 89168 700680 89220 700732
rect 349988 700680 350040 700732
rect 364248 700680 364300 700732
rect 429844 700680 429896 700732
rect 430028 700680 430080 700732
rect 559656 700680 559708 700732
rect 4068 700612 4120 700664
rect 266360 700612 266412 700664
rect 284392 700612 284444 700664
rect 332508 700612 332560 700664
rect 336556 700612 336608 700664
rect 580816 700612 580868 700664
rect 72976 700544 73028 700596
rect 344928 700544 344980 700596
rect 410432 700544 410484 700596
rect 494796 700544 494848 700596
rect 3240 700476 3292 700528
rect 286968 700476 287020 700528
rect 294512 700476 294564 700528
rect 300124 700476 300176 700528
rect 303528 700476 303580 700528
rect 329840 700476 329892 700528
rect 580724 700476 580776 700528
rect 40500 700408 40552 700460
rect 355048 700408 355100 700460
rect 24308 700340 24360 700392
rect 365076 700340 365128 700392
rect 8116 700272 8168 700324
rect 360016 700272 360068 700324
rect 137836 700204 137888 700256
rect 329748 700204 329800 700256
rect 154120 700136 154172 700188
rect 334808 700136 334860 700188
rect 202788 700068 202840 700120
rect 270684 700068 270736 700120
rect 283840 700068 283892 700120
rect 304540 700068 304592 700120
rect 478512 700068 478564 700120
rect 170312 700000 170364 700052
rect 324780 700000 324832 700052
rect 274272 699932 274324 699984
rect 413652 699932 413704 699984
rect 269212 699864 269264 699916
rect 397460 699864 397512 699916
rect 289452 699796 289504 699848
rect 348792 699796 348844 699848
rect 267648 699728 267700 699780
rect 299480 699728 299532 699780
rect 320824 699728 320876 699780
rect 543464 699728 543516 699780
rect 664 699660 716 699712
rect 435732 699660 435784 699712
rect 3700 699592 3752 699644
rect 332600 699592 332652 699644
rect 229008 699524 229060 699576
rect 579988 699524 580040 699576
rect 213828 699456 213880 699508
rect 580080 699456 580132 699508
rect 144368 699388 144420 699440
rect 580356 699388 580408 699440
rect 208952 699320 209004 699372
rect 579068 699320 579120 699372
rect 1584 699252 1636 699304
rect 374828 699252 374880 699304
rect 198740 699184 198792 699236
rect 580172 699184 580224 699236
rect 3056 699116 3108 699168
rect 395068 699116 395120 699168
rect 37280 699091 37332 699100
rect 37280 699057 37289 699091
rect 37289 699057 37323 699091
rect 37323 699057 37332 699091
rect 37280 699048 37332 699057
rect 42432 699091 42484 699100
rect 42432 699057 42441 699091
rect 42441 699057 42475 699091
rect 42475 699057 42484 699091
rect 42432 699048 42484 699057
rect 52368 699091 52420 699100
rect 52368 699057 52377 699091
rect 52377 699057 52411 699091
rect 52411 699057 52420 699091
rect 52368 699048 52420 699057
rect 67548 699091 67600 699100
rect 67548 699057 67557 699091
rect 67557 699057 67591 699091
rect 67591 699057 67600 699091
rect 67548 699048 67600 699057
rect 72792 699091 72844 699100
rect 72792 699057 72801 699091
rect 72801 699057 72835 699091
rect 72835 699057 72844 699091
rect 72792 699048 72844 699057
rect 82728 699091 82780 699100
rect 82728 699057 82737 699091
rect 82737 699057 82771 699091
rect 82771 699057 82780 699091
rect 82728 699048 82780 699057
rect 97908 699091 97960 699100
rect 97908 699057 97917 699091
rect 97917 699057 97951 699091
rect 97951 699057 97960 699091
rect 97908 699048 97960 699057
rect 103152 699091 103204 699100
rect 103152 699057 103161 699091
rect 103161 699057 103195 699091
rect 103195 699057 103204 699091
rect 103152 699048 103204 699057
rect 183560 699048 183612 699100
rect 580908 699048 580960 699100
rect 756 698980 808 699032
rect 405188 698980 405240 699032
rect 2596 698912 2648 698964
rect 420276 698980 420328 699032
rect 3148 698844 3200 698896
rect 425244 698980 425296 699032
rect 3332 698776 3384 698828
rect 455604 698980 455656 699032
rect 490932 699023 490984 699032
rect 490932 698989 490941 699023
rect 490941 698989 490975 699023
rect 490975 698989 490984 699023
rect 490932 698980 490984 698989
rect 495900 699023 495952 699032
rect 495900 698989 495909 699023
rect 495909 698989 495943 699023
rect 495943 698989 495952 699023
rect 495900 698980 495952 698989
rect 506020 699023 506072 699032
rect 506020 698989 506029 699023
rect 506029 698989 506063 699023
rect 506063 698989 506072 699023
rect 506020 698980 506072 698989
rect 511172 699023 511224 699032
rect 511172 698989 511181 699023
rect 511181 698989 511215 699023
rect 511215 698989 511224 699023
rect 511172 698980 511224 698989
rect 516140 699023 516192 699032
rect 516140 698989 516149 699023
rect 516149 698989 516183 699023
rect 516183 698989 516192 699023
rect 516140 698980 516192 698989
rect 521108 699023 521160 699032
rect 521108 698989 521117 699023
rect 521117 698989 521151 699023
rect 521151 698989 521160 699023
rect 521108 698980 521160 698989
rect 536380 699023 536432 699032
rect 536380 698989 536389 699023
rect 536389 698989 536423 699023
rect 536423 698989 536432 699023
rect 536380 698980 536432 698989
rect 546500 699023 546552 699032
rect 546500 698989 546509 699023
rect 546509 698989 546543 699023
rect 546543 698989 546552 699023
rect 546500 698980 546552 698989
rect 551468 699023 551520 699032
rect 551468 698989 551477 699023
rect 551477 698989 551511 699023
rect 551511 698989 551520 699023
rect 551468 698980 551520 698989
rect 566556 699023 566608 699032
rect 566556 698989 566565 699023
rect 566565 698989 566599 699023
rect 566599 698989 566608 699023
rect 566556 698980 566608 698989
rect 2228 698640 2280 698692
rect 3884 698572 3936 698624
rect 3976 698436 4028 698488
rect 3608 698300 3660 698352
rect 480 698164 532 698216
rect 388 698028 440 698080
rect 2136 697892 2188 697944
rect 204 697756 256 697808
rect 581828 697688 581880 697740
rect 112 697620 164 697672
rect 20 697552 72 697604
rect 3700 619556 3752 619608
rect 4528 619556 4580 619608
rect 583392 537820 583444 537872
rect 3240 516128 3292 516180
rect 4620 516128 4672 516180
rect 2780 462748 2832 462800
rect 4712 462748 4764 462800
rect 583392 431604 583444 431656
rect 583392 418276 583444 418328
rect 583392 351908 583444 351960
rect 583392 325252 583444 325304
rect 583392 312103 583444 312112
rect 583392 312069 583401 312103
rect 583401 312069 583435 312103
rect 583435 312069 583444 312103
rect 583392 312060 583444 312069
rect 2780 306212 2832 306264
rect 4804 306212 4856 306264
rect 583300 272255 583352 272264
rect 583300 272221 583309 272255
rect 583309 272221 583343 272255
rect 583343 272221 583352 272255
rect 583300 272212 583352 272221
rect 583208 245599 583260 245608
rect 583208 245565 583217 245599
rect 583217 245565 583251 245599
rect 583251 245565 583260 245599
rect 583208 245556 583260 245565
rect 583116 232407 583168 232416
rect 583116 232373 583125 232407
rect 583125 232373 583159 232407
rect 583159 232373 583168 232407
rect 583116 232364 583168 232373
rect 583024 205751 583076 205760
rect 583024 205717 583033 205751
rect 583033 205717 583067 205751
rect 583067 205717 583076 205751
rect 583024 205708 583076 205717
rect 582932 192559 582984 192568
rect 582932 192525 582941 192559
rect 582941 192525 582975 192559
rect 582975 192525 582984 192559
rect 582932 192516 582984 192525
rect 582840 179231 582892 179240
rect 582840 179197 582849 179231
rect 582849 179197 582883 179231
rect 582883 179197 582892 179231
rect 582840 179188 582892 179197
rect 582748 165903 582800 165912
rect 582748 165869 582757 165903
rect 582757 165869 582791 165903
rect 582791 165869 582800 165903
rect 582748 165860 582800 165869
rect 582656 152711 582708 152720
rect 582656 152677 582665 152711
rect 582665 152677 582699 152711
rect 582699 152677 582708 152711
rect 582656 152668 582708 152677
rect 582656 126012 582708 126064
rect 582656 112820 582708 112872
rect 582472 33056 582524 33108
rect 3424 4088 3476 4140
rect 582564 4088 582616 4140
rect 153016 4020 153068 4072
rect 155408 4020 155460 4072
rect 155408 3884 155460 3936
rect 157800 3884 157852 3936
rect 157800 3748 157852 3800
rect 160100 3748 160152 3800
rect 66720 3680 66772 3732
rect 70308 3680 70360 3732
rect 160100 3612 160152 3664
rect 162492 3612 162544 3664
rect 6460 3544 6512 3596
rect 10784 3544 10836 3596
rect 34796 3544 34848 3596
rect 38752 3544 38804 3596
rect 54944 3544 54996 3596
rect 58624 3544 58676 3596
rect 70308 3544 70360 3596
rect 73804 3544 73856 3596
rect 25320 3476 25372 3528
rect 29460 3476 29512 3528
rect 15936 3408 15988 3460
rect 20076 3408 20128 3460
rect 45468 3408 45520 3460
rect 49240 3408 49292 3460
rect 64328 3408 64380 3460
rect 67916 3408 67968 3460
rect 73804 3408 73856 3460
rect 77300 3408 77352 3460
rect 103336 3408 103388 3460
rect 106464 3408 106516 3460
rect 46664 3136 46716 3188
rect 50436 3136 50488 3188
rect 65524 3136 65576 3188
rect 69112 3136 69164 3188
rect 11152 3068 11204 3120
rect 15476 3068 15528 3120
rect 17040 3068 17092 3120
rect 21272 3068 21324 3120
rect 28908 3068 28960 3120
rect 32956 3068 33008 3120
rect 35992 3068 36044 3120
rect 39948 3068 40000 3120
rect 40684 3068 40736 3120
rect 44640 3068 44692 3120
rect 50160 3068 50212 3120
rect 53932 3068 53984 3120
rect 135260 3068 135312 3120
rect 137928 3068 137980 3120
rect 144736 3068 144788 3120
rect 147312 3068 147364 3120
rect 9956 3000 10008 3052
rect 14280 3000 14332 3052
rect 20628 3000 20680 3052
rect 24768 3000 24820 3052
rect 27712 3000 27764 3052
rect 31760 3000 31812 3052
rect 32404 3000 32456 3052
rect 36452 3000 36504 3052
rect 39580 3000 39632 3052
rect 43444 3000 43496 3052
rect 48964 3000 49016 3052
rect 52736 3000 52788 3052
rect 59636 3000 59688 3052
rect 63316 3000 63368 3052
rect 69112 3000 69164 3052
rect 72608 3000 72660 3052
rect 82084 3000 82136 3052
rect 85488 3000 85540 3052
rect 106924 3000 106976 3052
rect 109960 3000 110012 3052
rect 114008 3000 114060 3052
rect 116952 3000 117004 3052
rect 128176 3000 128228 3052
rect 130936 3000 130988 3052
rect 134156 3000 134208 3052
rect 136824 3000 136876 3052
rect 143540 3000 143592 3052
rect 146116 3000 146168 3052
rect 151820 3000 151872 3052
rect 154304 3000 154356 3052
rect 4068 2932 4120 2984
rect 8484 2932 8536 2984
rect 8760 2932 8812 2984
rect 13084 2932 13136 2984
rect 14740 2932 14792 2984
rect 18972 2932 19024 2984
rect 21824 2932 21876 2984
rect 25964 2932 26016 2984
rect 26516 2932 26568 2984
rect 30564 2932 30616 2984
rect 33600 2932 33652 2984
rect 37648 2932 37700 2984
rect 43076 2932 43128 2984
rect 46940 2932 46992 2984
rect 51356 2932 51408 2984
rect 55128 2932 55180 2984
rect 56048 2932 56100 2984
rect 59820 2932 59872 2984
rect 60832 2932 60884 2984
rect 64420 2932 64472 2984
rect 77392 2932 77444 2984
rect 80796 2932 80848 2984
rect 80888 2932 80940 2984
rect 84292 2932 84344 2984
rect 85672 2932 85724 2984
rect 88984 2932 89036 2984
rect 89168 2932 89220 2984
rect 92480 2932 92532 2984
rect 92756 2932 92808 2984
rect 95976 2932 96028 2984
rect 96252 2932 96304 2984
rect 99472 2932 99524 2984
rect 99840 2932 99892 2984
rect 102968 2932 103020 2984
rect 108120 2932 108172 2984
rect 111156 2932 111208 2984
rect 111616 2932 111668 2984
rect 114652 2932 114704 2984
rect 117596 2932 117648 2984
rect 120448 2932 120500 2984
rect 121092 2932 121144 2984
rect 123944 2932 123996 2984
rect 124680 2932 124732 2984
rect 127440 2932 127492 2984
rect 129372 2932 129424 2984
rect 132132 2932 132184 2984
rect 132960 2932 133012 2984
rect 135628 2932 135680 2984
rect 138848 2932 138900 2984
rect 141424 2932 141476 2984
rect 142436 2932 142488 2984
rect 144920 2932 144972 2984
rect 148324 2932 148376 2984
rect 150808 2932 150860 2984
rect 154212 2932 154264 2984
rect 156604 2932 156656 2984
rect 158996 2932 159048 2984
rect 161296 2932 161348 2984
rect 162492 2932 162544 2984
rect 164792 2932 164844 2984
rect 167184 2932 167236 2984
rect 169484 2932 169536 2984
rect 174268 2932 174320 2984
rect 176476 2932 176528 2984
rect 177856 2932 177908 2984
rect 179972 2932 180024 2984
rect 181444 2932 181496 2984
rect 183468 2932 183520 2984
rect 192024 2932 192076 2984
rect 193956 2932 194008 2984
rect 199108 2932 199160 2984
rect 200948 2932 201000 2984
rect 202696 2932 202748 2984
rect 204444 2932 204496 2984
rect 206192 2932 206244 2984
rect 207940 2932 207992 2984
rect 209780 2932 209832 2984
rect 211436 2932 211488 2984
rect 215668 2932 215720 2984
rect 217324 2932 217376 2984
rect 226340 2932 226392 2984
rect 227812 2932 227864 2984
rect 229836 2932 229888 2984
rect 231308 2932 231360 2984
rect 233424 2932 233476 2984
rect 234804 2932 234856 2984
rect 238116 2932 238168 2984
rect 239404 2932 239456 2984
rect 241704 2932 241756 2984
rect 242992 2932 243044 2984
rect 246396 2932 246448 2984
rect 247592 2932 247644 2984
rect 248880 2932 248932 2984
rect 249984 2932 250036 2984
rect 252376 2932 252428 2984
rect 253480 2932 253532 2984
rect 570788 2932 570840 2984
rect 573916 2932 573968 2984
rect 2872 2864 2924 2916
rect 7288 2864 7340 2916
rect 12348 2864 12400 2916
rect 16488 2864 16540 2916
rect 19432 2864 19484 2916
rect 23572 2864 23624 2916
rect 24216 2864 24268 2916
rect 28264 2864 28316 2916
rect 30104 2864 30156 2916
rect 34152 2864 34204 2916
rect 37188 2864 37240 2916
rect 41144 2864 41196 2916
rect 41880 2864 41932 2916
rect 45744 2864 45796 2916
rect 47860 2864 47912 2916
rect 51632 2864 51684 2916
rect 53748 2864 53800 2916
rect 57428 2864 57480 2916
rect 58440 2864 58492 2916
rect 62120 2864 62172 2916
rect 63224 2864 63276 2916
rect 66812 2864 66864 2916
rect 72608 2864 72660 2916
rect 76104 2864 76156 2916
rect 76196 2864 76248 2916
rect 79600 2864 79652 2916
rect 79692 2864 79744 2916
rect 83096 2864 83148 2916
rect 84476 2864 84528 2916
rect 87788 2864 87840 2916
rect 87972 2864 88024 2916
rect 91284 2864 91336 2916
rect 91560 2864 91612 2916
rect 94780 2864 94832 2916
rect 95148 2864 95200 2916
rect 98276 2864 98328 2916
rect 98644 2864 98696 2916
rect 101772 2864 101824 2916
rect 102232 2864 102284 2916
rect 105268 2864 105320 2916
rect 105728 2864 105780 2916
rect 108764 2864 108816 2916
rect 110512 2864 110564 2916
rect 113456 2864 113508 2916
rect 1676 2796 1728 2848
rect 5264 2796 5316 2848
rect 6092 2728 6144 2780
rect 7656 2796 7708 2848
rect 11980 2796 12032 2848
rect 13544 2796 13596 2848
rect 17776 2796 17828 2848
rect 18236 2796 18288 2848
rect 22468 2796 22520 2848
rect 23020 2796 23072 2848
rect 27068 2796 27120 2848
rect 31300 2796 31352 2848
rect 35256 2796 35308 2848
rect 38384 2796 38436 2848
rect 42248 2796 42300 2848
rect 44272 2796 44324 2848
rect 48136 2796 48188 2848
rect 52552 2796 52604 2848
rect 56232 2796 56284 2848
rect 57244 2796 57296 2848
rect 60924 2796 60976 2848
rect 62028 2796 62080 2848
rect 65616 2796 65668 2848
rect 67916 2796 67968 2848
rect 71412 2796 71464 2848
rect 71504 2796 71556 2848
rect 74908 2796 74960 2848
rect 75000 2796 75052 2848
rect 78404 2796 78456 2848
rect 78588 2796 78640 2848
rect 81900 2796 81952 2848
rect 83280 2796 83332 2848
rect 86592 2796 86644 2848
rect 86868 2796 86920 2848
rect 90088 2796 90140 2848
rect 90364 2796 90416 2848
rect 93584 2796 93636 2848
rect 93952 2796 94004 2848
rect 97080 2796 97132 2848
rect 97448 2796 97500 2848
rect 100576 2796 100628 2848
rect 101036 2796 101088 2848
rect 104072 2796 104124 2848
rect 104532 2796 104584 2848
rect 107568 2796 107620 2848
rect 109316 2796 109368 2848
rect 112260 2796 112312 2848
rect 112812 2796 112864 2848
rect 115756 2864 115808 2916
rect 116400 2864 116452 2916
rect 119252 2864 119304 2916
rect 119896 2864 119948 2916
rect 122748 2864 122800 2916
rect 123484 2864 123536 2916
rect 126244 2864 126296 2916
rect 126980 2864 127032 2916
rect 129740 2864 129792 2916
rect 131764 2864 131816 2916
rect 134432 2864 134484 2916
rect 137652 2864 137704 2916
rect 140320 2864 140372 2916
rect 141240 2864 141292 2916
rect 143816 2864 143868 2916
rect 147128 2864 147180 2916
rect 149612 2864 149664 2916
rect 150624 2864 150676 2916
rect 153108 2864 153160 2916
rect 163688 2864 163740 2916
rect 165988 2864 166040 2916
rect 166080 2864 166132 2916
rect 168288 2864 168340 2916
rect 169576 2864 169628 2916
rect 171784 2864 171836 2916
rect 115204 2796 115256 2848
rect 118148 2796 118200 2848
rect 118792 2796 118844 2848
rect 121644 2796 121696 2848
rect 122288 2796 122340 2848
rect 125140 2796 125192 2848
rect 125876 2796 125928 2848
rect 128636 2796 128688 2848
rect 130568 2796 130620 2848
rect 133236 2796 133288 2848
rect 136456 2796 136508 2848
rect 139124 2796 139176 2848
rect 140044 2796 140096 2848
rect 142620 2796 142672 2848
rect 145932 2796 145984 2848
rect 148416 2796 148468 2848
rect 149520 2796 149572 2848
rect 151912 2796 151964 2848
rect 156604 2796 156656 2848
rect 158904 2796 158956 2848
rect 161296 2796 161348 2848
rect 163596 2796 163648 2848
rect 164884 2796 164936 2848
rect 167092 2796 167144 2848
rect 168380 2796 168432 2848
rect 170588 2796 170640 2848
rect 170772 2796 170824 2848
rect 172980 2864 173032 2916
rect 173164 2864 173216 2916
rect 175280 2864 175332 2916
rect 176660 2864 176712 2916
rect 178776 2864 178828 2916
rect 180248 2864 180300 2916
rect 182272 2864 182324 2916
rect 183744 2864 183796 2916
rect 185768 2864 185820 2916
rect 186136 2864 186188 2916
rect 188160 2864 188212 2916
rect 188528 2864 188580 2916
rect 190460 2864 190512 2916
rect 171968 2796 172020 2848
rect 174084 2796 174136 2848
rect 175464 2796 175516 2848
rect 177580 2796 177632 2848
rect 179052 2796 179104 2848
rect 181076 2796 181128 2848
rect 182548 2796 182600 2848
rect 184572 2796 184624 2848
rect 184940 2796 184992 2848
rect 186964 2796 187016 2848
rect 187332 2796 187384 2848
rect 189264 2796 189316 2848
rect 189724 2796 189776 2848
rect 191656 2864 191708 2916
rect 193220 2864 193272 2916
rect 195152 2864 195204 2916
rect 195612 2864 195664 2916
rect 197452 2864 197504 2916
rect 197912 2864 197964 2916
rect 199752 2864 199804 2916
rect 200304 2864 200356 2916
rect 202144 2864 202196 2916
rect 203892 2864 203944 2916
rect 205640 2864 205692 2916
rect 207388 2864 207440 2916
rect 209136 2864 209188 2916
rect 210976 2864 211028 2916
rect 212632 2864 212684 2916
rect 213368 2864 213420 2916
rect 214932 2864 214984 2916
rect 216864 2864 216916 2916
rect 218428 2864 218480 2916
rect 219256 2864 219308 2916
rect 220820 2864 220872 2916
rect 221556 2864 221608 2916
rect 223120 2864 223172 2916
rect 223948 2864 224000 2916
rect 225420 2864 225472 2916
rect 227536 2864 227588 2916
rect 228916 2864 228968 2916
rect 231032 2864 231084 2916
rect 232412 2864 232464 2916
rect 234620 2864 234672 2916
rect 235908 2864 235960 2916
rect 237012 2864 237064 2916
rect 238300 2864 238352 2916
rect 240508 2864 240560 2916
rect 241796 2864 241848 2916
rect 245200 2864 245252 2916
rect 246488 2864 246540 2916
rect 540428 2864 540480 2916
rect 543188 2864 543240 2916
rect 547420 2864 547472 2916
rect 550272 2864 550324 2916
rect 553400 2864 553452 2916
rect 556160 2864 556212 2916
rect 561680 2864 561732 2916
rect 564440 2864 564492 2916
rect 568580 2864 568632 2916
rect 571524 2864 571576 2916
rect 190828 2796 190880 2848
rect 192760 2796 192812 2848
rect 194416 2796 194468 2848
rect 196256 2796 196308 2848
rect 196808 2796 196860 2848
rect 198648 2796 198700 2848
rect 201500 2796 201552 2848
rect 203248 2796 203300 2848
rect 205088 2796 205140 2848
rect 206744 2796 206796 2848
rect 208584 2796 208636 2848
rect 210240 2796 210292 2848
rect 212172 2796 212224 2848
rect 213736 2796 213788 2848
rect 214472 2796 214524 2848
rect 216128 2796 216180 2848
rect 218060 2796 218112 2848
rect 219624 2796 219676 2848
rect 220452 2796 220504 2848
rect 221924 2796 221976 2848
rect 222752 2796 222804 2848
rect 224316 2796 224368 2848
rect 225144 2796 225196 2848
rect 226616 2796 226668 2848
rect 228732 2796 228784 2848
rect 230112 2796 230164 2848
rect 232228 2796 232280 2848
rect 233608 2796 233660 2848
rect 235816 2796 235868 2848
rect 237104 2796 237156 2848
rect 239312 2796 239364 2848
rect 240600 2796 240652 2848
rect 242900 2796 242952 2848
rect 244096 2796 244148 2848
rect 244188 2796 244240 2848
rect 245292 2796 245344 2848
rect 247592 2796 247644 2848
rect 248788 2796 248840 2848
rect 249984 2796 250036 2848
rect 251088 2796 251140 2848
rect 253480 2796 253532 2848
rect 254584 2796 254636 2848
rect 254676 2796 254728 2848
rect 255780 2796 255832 2848
rect 255872 2796 255924 2848
rect 256976 2796 257028 2848
rect 257068 2796 257120 2848
rect 258080 2796 258132 2848
rect 259460 2796 259512 2848
rect 260472 2796 260524 2848
rect 260656 2796 260708 2848
rect 261576 2796 261628 2848
rect 261760 2796 261812 2848
rect 262772 2796 262824 2848
rect 262956 2796 263008 2848
rect 263968 2796 264020 2848
rect 264152 2796 264204 2848
rect 265072 2796 265124 2848
rect 266544 2796 266596 2848
rect 267464 2796 267516 2848
rect 267740 2796 267792 2848
rect 268660 2796 268712 2848
rect 268844 2796 268896 2848
rect 269764 2796 269816 2848
rect 270040 2796 270092 2848
rect 270960 2796 271012 2848
rect 271236 2796 271288 2848
rect 272156 2796 272208 2848
rect 272432 2796 272484 2848
rect 273260 2796 273312 2848
rect 273628 2796 273680 2848
rect 274456 2796 274508 2848
rect 274824 2796 274876 2848
rect 275652 2796 275704 2848
rect 277124 2796 277176 2848
rect 277952 2796 278004 2848
rect 278320 2796 278372 2848
rect 279148 2796 279200 2848
rect 279516 2796 279568 2848
rect 280252 2796 280304 2848
rect 280712 2796 280764 2848
rect 281448 2796 281500 2848
rect 281908 2796 281960 2848
rect 282644 2796 282696 2848
rect 284300 2796 284352 2848
rect 284944 2796 284996 2848
rect 285404 2796 285456 2848
rect 286140 2796 286192 2848
rect 286600 2796 286652 2848
rect 287244 2796 287296 2848
rect 287796 2796 287848 2848
rect 288440 2796 288492 2848
rect 288992 2796 289044 2848
rect 289636 2796 289688 2848
rect 291384 2796 291436 2848
rect 291936 2796 291988 2848
rect 292580 2796 292632 2848
rect 293132 2796 293184 2848
rect 293684 2796 293736 2848
rect 294328 2796 294380 2848
rect 294880 2796 294932 2848
rect 295432 2796 295484 2848
rect 296076 2796 296128 2848
rect 296628 2796 296680 2848
rect 298468 2796 298520 2848
rect 298928 2796 298980 2848
rect 299664 2796 299716 2848
rect 300124 2796 300176 2848
rect 300768 2796 300820 2848
rect 301320 2796 301372 2848
rect 301964 2796 302016 2848
rect 302424 2796 302476 2848
rect 303160 2796 303212 2848
rect 303620 2796 303672 2848
rect 368940 2796 368992 2848
rect 369400 2796 369452 2848
rect 370136 2796 370188 2848
rect 370596 2796 370648 2848
rect 375932 2796 375984 2848
rect 376484 2796 376536 2848
rect 377128 2796 377180 2848
rect 377680 2796 377732 2848
rect 382924 2796 382976 2848
rect 383568 2796 383620 2848
rect 384120 2796 384172 2848
rect 384764 2796 384816 2848
rect 386420 2796 386472 2848
rect 387156 2796 387208 2848
rect 391112 2796 391164 2848
rect 391848 2796 391900 2848
rect 393412 2796 393464 2848
rect 394240 2796 394292 2848
rect 400496 2796 400548 2848
rect 401324 2796 401376 2848
rect 401600 2796 401652 2848
rect 402520 2796 402572 2848
rect 407488 2796 407540 2848
rect 408408 2796 408460 2848
rect 408592 2796 408644 2848
rect 409604 2796 409656 2848
rect 415584 2796 415636 2848
rect 416688 2796 416740 2848
rect 431960 2796 432012 2848
rect 433248 2796 433300 2848
rect 9588 2728 9640 2780
rect 470416 2728 470468 2780
rect 472256 2796 472308 2848
rect 478604 2728 478656 2780
rect 480536 2796 480588 2848
rect 485596 2728 485648 2780
rect 487620 2796 487672 2848
rect 492680 2796 492732 2848
rect 494704 2796 494756 2848
rect 493784 2728 493836 2780
rect 495900 2796 495952 2848
rect 500776 2728 500828 2780
rect 502984 2796 503036 2848
rect 503168 2728 503220 2780
rect 505376 2796 505428 2848
rect 507860 2796 507912 2848
rect 510068 2796 510120 2848
rect 510160 2728 510212 2780
rect 512460 2796 512512 2848
rect 515956 2728 516008 2780
rect 518348 2796 518400 2848
rect 517152 2728 517204 2780
rect 519544 2796 519596 2848
rect 519452 2728 519504 2780
rect 521844 2796 521896 2848
rect 523040 2796 523092 2848
rect 525432 2796 525484 2848
rect 524144 2728 524196 2780
rect 526628 2796 526680 2848
rect 525248 2660 525300 2712
rect 527824 2796 527876 2848
rect 531136 2728 531188 2780
rect 533712 2796 533764 2848
rect 532332 2660 532384 2712
rect 534908 2796 534960 2848
rect 534632 2728 534684 2780
rect 537208 2796 537260 2848
rect 538220 2796 538272 2848
rect 540796 2796 540848 2848
rect 539324 2728 539376 2780
rect 541992 2796 542044 2848
rect 541624 2728 541676 2780
rect 544384 2796 544436 2848
rect 542820 2728 542872 2780
rect 545488 2796 545540 2848
rect 546316 2728 546368 2780
rect 549076 2796 549128 2848
rect 548616 2728 548668 2780
rect 551468 2796 551520 2848
rect 549812 2660 549864 2712
rect 552664 2796 552716 2848
rect 552112 2728 552164 2780
rect 554964 2796 555016 2848
rect 554504 2660 554556 2712
rect 557356 2796 557408 2848
rect 555608 2728 555660 2780
rect 558552 2796 558604 2848
rect 558000 2728 558052 2780
rect 560852 2796 560904 2848
rect 560300 2728 560352 2780
rect 563244 2796 563296 2848
rect 562600 2660 562652 2712
rect 565636 2796 565688 2848
rect 566832 2796 566884 2848
rect 563796 2592 563848 2644
rect 566096 2728 566148 2780
rect 569132 2796 569184 2848
rect 567292 2728 567344 2780
rect 570328 2796 570380 2848
rect 569592 2660 569644 2712
rect 572720 2796 572772 2848
rect 571984 2728 572036 2780
rect 575112 2796 575164 2848
rect 574284 2728 574336 2780
rect 577412 2796 577464 2848
rect 577780 2728 577832 2780
rect 582196 2796 582248 2848
rect 424968 2524 425020 2576
rect 426072 2524 426124 2576
rect 428464 2456 428516 2508
rect 429568 2456 429620 2508
rect 423772 2388 423824 2440
rect 424968 2388 425020 2440
rect 427268 2320 427320 2372
rect 428464 2320 428516 2372
rect 511264 2320 511316 2372
rect 513564 2320 513616 2372
rect 514760 2320 514812 2372
rect 517152 2320 517204 2372
rect 304356 2252 304408 2304
rect 304816 2252 304868 2304
rect 380624 2252 380676 2304
rect 381176 2252 381228 2304
rect 398104 2252 398156 2304
rect 398932 2252 398984 2304
rect 402796 2252 402848 2304
rect 403624 2252 403676 2304
rect 409788 2252 409840 2304
rect 410800 2252 410852 2304
rect 412088 2252 412140 2304
rect 413100 2252 413152 2304
rect 414480 2252 414532 2304
rect 415492 2252 415544 2304
rect 422576 2252 422628 2304
rect 423772 2252 423824 2304
rect 429660 2252 429712 2304
rect 430856 2252 430908 2304
rect 435456 2252 435508 2304
rect 436744 2252 436796 2304
rect 438952 2252 439004 2304
rect 440332 2252 440384 2304
rect 441252 2252 441304 2304
rect 442632 2252 442684 2304
rect 450636 2252 450688 2304
rect 452108 2252 452160 2304
rect 452936 2252 452988 2304
rect 454500 2252 454552 2304
rect 486792 2252 486844 2304
rect 488816 2252 488868 2304
rect 494980 2252 495032 2304
rect 497096 2252 497148 2304
rect 497280 2252 497332 2304
rect 499396 2252 499448 2304
rect 520648 2252 520700 2304
rect 523040 2252 523092 2304
rect 526444 2252 526496 2304
rect 529020 2252 529072 2304
rect 535828 2252 535880 2304
rect 572 2184 624 2236
rect 4988 2184 5040 2236
rect 251180 2184 251232 2236
rect 252284 2184 252336 2236
rect 258264 2184 258316 2236
rect 259276 2184 259328 2236
rect 290188 2184 290240 2236
rect 290740 2184 290792 2236
rect 297272 2184 297324 2236
rect 297824 2184 297876 2236
rect 367744 2184 367796 2236
rect 368204 2184 368256 2236
rect 373632 2184 373684 2236
rect 374092 2184 374144 2236
rect 374828 2184 374880 2236
rect 375288 2184 375340 2236
rect 378324 2184 378376 2236
rect 378876 2184 378928 2236
rect 379428 2184 379480 2236
rect 379980 2184 380032 2236
rect 385316 2184 385368 2236
rect 385960 2184 386012 2236
rect 387616 2184 387668 2236
rect 388260 2184 388312 2236
rect 388812 2184 388864 2236
rect 389456 2184 389508 2236
rect 389916 2184 389968 2236
rect 390652 2184 390704 2236
rect 392308 2184 392360 2236
rect 393044 2184 393096 2236
rect 394608 2184 394660 2236
rect 395344 2184 395396 2236
rect 395804 2184 395856 2236
rect 396540 2184 396592 2236
rect 399300 2184 399352 2236
rect 400128 2184 400180 2236
rect 410984 2184 411036 2236
rect 411904 2184 411956 2236
rect 417976 2184 418028 2236
rect 418988 2184 419040 2236
rect 426164 2184 426216 2236
rect 427268 2184 427320 2236
rect 437756 2184 437808 2236
rect 439136 2184 439188 2236
rect 443644 2184 443696 2236
rect 445024 2184 445076 2236
rect 451832 2184 451884 2236
rect 453304 2184 453356 2236
rect 458824 2184 458876 2236
rect 460388 2184 460440 2236
rect 463424 2184 463476 2236
rect 465172 2184 465224 2236
rect 466920 2184 466972 2236
rect 468668 2184 468720 2236
rect 471612 2184 471664 2236
rect 473452 2184 473504 2236
rect 473912 2184 473964 2236
rect 475752 2184 475804 2236
rect 476304 2184 476356 2236
rect 478144 2184 478196 2236
rect 479800 2184 479852 2236
rect 481732 2184 481784 2236
rect 483296 2184 483348 2236
rect 485228 2184 485280 2236
rect 487988 2184 488040 2236
rect 489920 2184 489972 2236
rect 496084 2184 496136 2236
rect 498200 2184 498252 2236
rect 501972 2184 502024 2236
rect 504180 2184 504232 2236
rect 504272 2184 504324 2236
rect 506480 2184 506532 2236
rect 506664 2184 506716 2236
rect 508872 2184 508924 2236
rect 508964 2184 509016 2236
rect 511264 2184 511316 2236
rect 512552 2184 512604 2236
rect 514760 2184 514812 2236
rect 518256 2184 518308 2236
rect 520740 2184 520792 2236
rect 521752 2184 521804 2236
rect 524236 2184 524288 2236
rect 527640 2184 527692 2236
rect 530124 2184 530176 2236
rect 533436 2184 533488 2236
rect 536104 2184 536156 2236
rect 536932 2252 536984 2304
rect 539600 2252 539652 2304
rect 545120 2252 545172 2304
rect 547880 2252 547932 2304
rect 559104 2252 559156 2304
rect 562048 2252 562100 2304
rect 538404 2184 538456 2236
rect 543924 2184 543976 2236
rect 546684 2184 546736 2236
rect 550916 2184 550968 2236
rect 553768 2184 553820 2236
rect 556804 2184 556856 2236
rect 559748 2184 559800 2236
rect 564992 2184 565044 2236
rect 568028 2184 568080 2236
rect 575480 2184 575532 2236
rect 578608 2184 578660 2236
rect 578976 2184 579028 2236
rect 583392 2184 583444 2236
rect 372436 2116 372488 2168
rect 372896 2116 372948 2168
rect 416780 2116 416832 2168
rect 417884 2116 417936 2168
rect 420276 2116 420328 2168
rect 421380 2116 421432 2168
rect 430764 2116 430816 2168
rect 432052 2116 432104 2168
rect 434260 2116 434312 2168
rect 435548 2116 435600 2168
rect 436652 2116 436704 2168
rect 437940 2116 437992 2168
rect 444748 2116 444800 2168
rect 446220 2116 446272 2168
rect 447140 2116 447192 2168
rect 448612 2116 448664 2168
rect 454132 2116 454184 2168
rect 455696 2116 455748 2168
rect 573088 2116 573140 2168
rect 576308 2116 576360 2168
rect 406292 2048 406344 2100
rect 407212 2048 407264 2100
rect 449440 2048 449492 2100
rect 450912 2048 450964 2100
rect 455328 2048 455380 2100
rect 456892 2048 456944 2100
rect 576584 2048 576636 2100
rect 581000 2048 581052 2100
rect 265348 1980 265400 2032
rect 266268 1980 266320 2032
rect 381820 1980 381872 2032
rect 382372 1980 382424 2032
rect 440148 1980 440200 2032
rect 441528 1980 441580 2032
rect 276020 1912 276072 1964
rect 276756 1912 276808 1964
rect 442448 1912 442500 1964
rect 443828 1912 443880 1964
rect 489092 1912 489144 1964
rect 491116 1912 491168 1964
rect 513656 1912 513708 1964
rect 515956 1912 516008 1964
rect 528836 1912 528888 1964
rect 531320 1912 531372 1964
rect 419080 1844 419132 1896
rect 420184 1844 420236 1896
rect 459928 1844 459980 1896
rect 461584 1844 461636 1896
rect 396908 1776 396960 1828
rect 397736 1776 397788 1828
rect 490288 1776 490340 1828
rect 492312 1776 492364 1828
rect 498476 1776 498528 1828
rect 500592 1776 500644 1828
rect 505468 1776 505520 1828
rect 507676 1776 507728 1828
rect 529940 1776 529992 1828
rect 532516 1776 532568 1828
rect 462320 1708 462372 1760
rect 463976 1708 464028 1760
rect 482100 1708 482152 1760
rect 484032 1708 484084 1760
rect 491484 1708 491536 1760
rect 493508 1708 493560 1760
rect 499580 1708 499632 1760
rect 501788 1708 501840 1760
rect 283104 1640 283156 1692
rect 283748 1640 283800 1692
rect 421472 1640 421524 1692
rect 422576 1640 422628 1692
rect 445944 1640 445996 1692
rect 447416 1640 447468 1692
rect 448244 1640 448296 1692
rect 449808 1640 449860 1692
rect 472808 1640 472860 1692
rect 474556 1640 474608 1692
rect 475108 1640 475160 1692
rect 476948 1640 477000 1692
rect 468116 1572 468168 1624
rect 469864 1572 469916 1624
rect 480996 1572 481048 1624
rect 482836 1572 482888 1624
rect 484492 1572 484544 1624
rect 486424 1572 486476 1624
rect 405096 1504 405148 1556
rect 406016 1504 406068 1556
rect 413284 1504 413336 1556
rect 414296 1504 414348 1556
rect 433156 1504 433208 1556
rect 434444 1504 434496 1556
rect 456432 1504 456484 1556
rect 458088 1504 458140 1556
rect 465816 1504 465868 1556
rect 467472 1504 467524 1556
rect 469312 1504 469364 1556
rect 471060 1504 471112 1556
rect 477500 1504 477552 1556
rect 479340 1504 479392 1556
rect 457628 1436 457680 1488
rect 459192 1436 459244 1488
rect 461124 1436 461176 1488
rect 462780 1436 462832 1488
rect 464620 1436 464672 1488
rect 466276 1436 466328 1488
rect 403992 1368 404044 1420
rect 404820 1368 404872 1420
<< metal2 >>
rect 6920 703860 6972 703866
rect 6920 703802 6972 703808
rect 1492 703384 1544 703390
rect 1492 703326 1544 703332
rect 572 701616 624 701622
rect 572 701558 624 701564
rect 294 701448 350 701457
rect 294 701383 350 701392
rect 204 697808 256 697814
rect 204 697750 256 697756
rect 112 697672 164 697678
rect 112 697614 164 697620
rect 20 697604 72 697610
rect 20 697546 72 697552
rect 32 33017 60 697546
rect 124 71913 152 697614
rect 216 111217 244 697750
rect 308 151814 336 701383
rect 480 698216 532 698222
rect 480 698158 532 698164
rect 388 698080 440 698086
rect 388 698022 440 698028
rect 400 229094 428 698022
rect 492 267186 520 698158
rect 584 345409 612 701558
rect 664 699712 716 699718
rect 664 699654 716 699660
rect 676 449585 704 699654
rect 756 699032 808 699038
rect 756 698974 808 698980
rect 768 553897 796 698974
rect 846 697096 902 697105
rect 846 697031 902 697040
rect 860 606121 888 697031
rect 1504 684321 1532 703326
rect 1676 703248 1728 703254
rect 1676 703190 1728 703196
rect 1584 699304 1636 699310
rect 1584 699246 1636 699252
rect 1490 684312 1546 684321
rect 1490 684247 1546 684256
rect 1596 658209 1624 699246
rect 1582 658200 1638 658209
rect 1582 658135 1638 658144
rect 1688 632097 1716 703190
rect 1768 703112 1820 703118
rect 1768 703054 1820 703060
rect 1674 632088 1730 632097
rect 1674 632023 1730 632032
rect 846 606112 902 606121
rect 846 606047 902 606056
rect 1780 580009 1808 703054
rect 1860 702908 1912 702914
rect 1860 702850 1912 702856
rect 1766 580000 1822 580009
rect 1766 579935 1822 579944
rect 754 553888 810 553897
rect 754 553823 810 553832
rect 1872 527921 1900 702850
rect 2412 702772 2464 702778
rect 2412 702714 2464 702720
rect 2042 701720 2098 701729
rect 2042 701655 2098 701664
rect 1950 698184 2006 698193
rect 1950 698119 2006 698128
rect 1858 527912 1914 527921
rect 1858 527847 1914 527856
rect 1964 475697 1992 698119
rect 1950 475688 2006 475697
rect 1950 475623 2006 475632
rect 662 449576 718 449585
rect 662 449511 718 449520
rect 570 345400 626 345409
rect 570 345335 626 345344
rect 570 267200 626 267209
rect 492 267158 570 267186
rect 570 267135 626 267144
rect 400 229066 612 229094
rect 584 214985 612 229066
rect 570 214976 626 214985
rect 570 214911 626 214920
rect 308 151786 612 151814
rect 584 136785 612 151786
rect 570 136776 626 136785
rect 570 136711 626 136720
rect 202 111208 258 111217
rect 202 111143 258 111152
rect 110 71904 166 71913
rect 110 71839 166 71848
rect 2056 58585 2084 701655
rect 2228 698692 2280 698698
rect 2228 698634 2280 698640
rect 2136 697944 2188 697950
rect 2136 697886 2188 697892
rect 2148 162897 2176 697886
rect 2240 241097 2268 698634
rect 2318 697504 2374 697513
rect 2318 697439 2374 697448
rect 2332 319297 2360 697439
rect 2424 423609 2452 702714
rect 4712 701820 4764 701826
rect 4712 701762 4764 701768
rect 4526 701312 4582 701321
rect 4526 701247 4582 701256
rect 3792 700868 3844 700874
rect 3792 700810 3844 700816
rect 3240 700528 3292 700534
rect 3240 700470 3292 700476
rect 3056 699168 3108 699174
rect 3056 699110 3108 699116
rect 2596 698964 2648 698970
rect 2596 698906 2648 698912
rect 2502 697776 2558 697785
rect 2502 697711 2558 697720
rect 2410 423600 2466 423609
rect 2410 423535 2466 423544
rect 2516 371385 2544 697711
rect 2608 501809 2636 698906
rect 2686 697912 2742 697921
rect 2686 697847 2742 697856
rect 2594 501800 2650 501809
rect 2594 501735 2650 501744
rect 2700 397497 2728 697847
rect 3068 619177 3096 699110
rect 3148 698896 3200 698902
rect 3148 698838 3200 698844
rect 3054 619168 3110 619177
rect 3054 619103 3110 619112
rect 3160 514865 3188 698838
rect 3252 566953 3280 700470
rect 3422 700360 3478 700369
rect 3422 700295 3478 700304
rect 3332 698828 3384 698834
rect 3332 698770 3384 698776
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3240 516180 3292 516186
rect 3240 516122 3292 516128
rect 3146 514856 3202 514865
rect 3146 514791 3202 514800
rect 2780 462800 2832 462806
rect 2780 462742 2832 462748
rect 2792 462641 2820 462742
rect 2778 462632 2834 462641
rect 2778 462567 2834 462576
rect 2686 397488 2742 397497
rect 2686 397423 2742 397432
rect 2502 371376 2558 371385
rect 2502 371311 2558 371320
rect 2318 319288 2374 319297
rect 2318 319223 2374 319232
rect 2780 306264 2832 306270
rect 2778 306232 2780 306241
rect 2832 306232 2834 306241
rect 2778 306167 2834 306176
rect 3252 254153 3280 516122
rect 3344 410553 3372 698770
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3238 254144 3294 254153
rect 3238 254079 3294 254088
rect 2226 241088 2282 241097
rect 2226 241023 2282 241032
rect 2134 162888 2190 162897
rect 2134 162823 2190 162832
rect 2042 58576 2098 58585
rect 2042 58511 2098 58520
rect 18 33008 74 33017
rect 18 32943 74 32952
rect 3436 19417 3464 700295
rect 3700 699644 3752 699650
rect 3700 699586 3752 699592
rect 3514 698456 3570 698465
rect 3514 698391 3570 698400
rect 3528 84697 3556 698391
rect 3608 698352 3660 698358
rect 3608 698294 3660 698300
rect 3620 97617 3648 698294
rect 3712 671265 3740 699586
rect 3698 671256 3754 671265
rect 3698 671191 3754 671200
rect 3700 619608 3752 619614
rect 3700 619550 3752 619556
rect 3606 97608 3662 97617
rect 3606 97543 3662 97552
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3712 45529 3740 619550
rect 3804 149841 3832 700810
rect 4068 700664 4120 700670
rect 4068 700606 4120 700612
rect 3884 698624 3936 698630
rect 3884 698566 3936 698572
rect 3896 188873 3924 698566
rect 3976 698488 4028 698494
rect 3976 698430 4028 698436
rect 3988 201929 4016 698430
rect 4080 293185 4108 700606
rect 4540 619614 4568 701247
rect 4620 701208 4672 701214
rect 4620 701150 4672 701156
rect 4528 619608 4580 619614
rect 4528 619550 4580 619556
rect 4632 516186 4660 701150
rect 4620 516180 4672 516186
rect 4620 516122 4672 516128
rect 4724 462806 4752 701762
rect 4896 701548 4948 701554
rect 4896 701490 4948 701496
rect 4804 701412 4856 701418
rect 4804 701354 4856 701360
rect 4712 462800 4764 462806
rect 4712 462742 4764 462748
rect 4816 367094 4844 701354
rect 4632 367066 4844 367094
rect 4632 357434 4660 367066
rect 4802 358456 4858 358465
rect 4908 358442 4936 701490
rect 6932 699516 6960 703802
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 233884 703520 233936 703526
rect 235142 703520 235254 704960
rect 238944 703724 238996 703730
rect 238944 703666 238996 703672
rect 8128 700330 8156 703520
rect 22008 702636 22060 702642
rect 22008 702578 22060 702584
rect 11888 702568 11940 702574
rect 11888 702510 11940 702516
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 11900 699516 11928 702510
rect 22020 699516 22048 702578
rect 24320 700398 24348 703520
rect 32128 701752 32180 701758
rect 32128 701694 32180 701700
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 27066 699816 27122 699825
rect 27066 699751 27122 699760
rect 27080 699516 27108 699751
rect 32140 699516 32168 701694
rect 40512 700466 40540 703520
rect 57336 702364 57388 702370
rect 57336 702306 57388 702312
rect 47216 701888 47268 701894
rect 47216 701830 47268 701836
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 47228 699516 47256 701830
rect 57348 699516 57376 702306
rect 72988 700602 73016 703520
rect 87604 701276 87656 701282
rect 87604 701218 87656 701224
rect 77484 701140 77536 701146
rect 77484 701082 77536 701088
rect 72976 700596 73028 700602
rect 72976 700538 73028 700544
rect 62394 699952 62450 699961
rect 62394 699887 62450 699896
rect 62408 699516 62436 699887
rect 77496 699516 77524 701082
rect 87616 699516 87644 701218
rect 89180 700738 89208 703520
rect 92664 701344 92716 701350
rect 92664 701286 92716 701292
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 92676 699516 92704 701286
rect 105464 700806 105492 703520
rect 127992 702704 128044 702710
rect 127992 702646 128044 702652
rect 122932 701684 122984 701690
rect 122932 701626 122984 701632
rect 117872 701480 117924 701486
rect 117872 701422 117924 701428
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 107750 700088 107806 700097
rect 107750 700023 107806 700032
rect 107764 699516 107792 700023
rect 117884 699516 117912 701422
rect 122944 699516 122972 701626
rect 128004 699516 128032 702646
rect 133052 702092 133104 702098
rect 133052 702034 133104 702040
rect 132684 701752 132736 701758
rect 132684 701694 132736 701700
rect 37214 699106 37320 699122
rect 42182 699106 42472 699122
rect 52302 699106 52408 699122
rect 67482 699106 67588 699122
rect 72450 699106 72832 699122
rect 82570 699106 82768 699122
rect 97750 699106 97948 699122
rect 102810 699106 103192 699122
rect 37214 699100 37332 699106
rect 37214 699094 37280 699100
rect 42182 699100 42484 699106
rect 42182 699094 42432 699100
rect 37280 699042 37332 699048
rect 52302 699100 52420 699106
rect 52302 699094 52368 699100
rect 42432 699042 42484 699048
rect 67482 699100 67600 699106
rect 67482 699094 67548 699100
rect 52368 699042 52420 699048
rect 72450 699100 72844 699106
rect 72450 699094 72792 699100
rect 67548 699042 67600 699048
rect 82570 699100 82780 699106
rect 82570 699094 82728 699100
rect 72792 699042 72844 699048
rect 97750 699100 97960 699106
rect 97750 699094 97908 699100
rect 82728 699042 82780 699048
rect 102810 699100 103204 699106
rect 102810 699094 103152 699100
rect 97908 699042 97960 699048
rect 103152 699042 103204 699048
rect 132696 699009 132724 701694
rect 133064 699516 133092 702034
rect 137848 700262 137876 703520
rect 138020 702024 138072 702030
rect 138020 701966 138072 701972
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 138032 699516 138060 701966
rect 144368 701888 144420 701894
rect 144368 701830 144420 701836
rect 153200 701888 153252 701894
rect 153200 701830 153252 701836
rect 144380 699446 144408 701830
rect 148140 701752 148192 701758
rect 148140 701694 148192 701700
rect 148152 699516 148180 701694
rect 153212 699516 153240 701830
rect 154132 700194 154160 703520
rect 158260 702840 158312 702846
rect 158260 702782 158312 702788
rect 154120 700188 154172 700194
rect 154120 700130 154172 700136
rect 158272 699516 158300 702782
rect 168288 702160 168340 702166
rect 168288 702102 168340 702108
rect 168300 699516 168328 702102
rect 170324 700058 170352 703520
rect 188528 703180 188580 703186
rect 188528 703122 188580 703128
rect 178408 703044 178460 703050
rect 178408 702986 178460 702992
rect 173348 702976 173400 702982
rect 173348 702918 173400 702924
rect 170312 700052 170364 700058
rect 170312 699994 170364 700000
rect 173360 699516 173388 702918
rect 178420 699516 178448 702986
rect 188540 699516 188568 703122
rect 202800 700126 202828 703520
rect 218796 703452 218848 703458
rect 218796 703394 218848 703400
rect 203616 703316 203668 703322
rect 203616 703258 203668 703264
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 203628 699516 203656 703258
rect 218058 701584 218114 701593
rect 218058 701519 218114 701528
rect 218072 700874 218100 701519
rect 218060 700868 218112 700874
rect 218060 700810 218112 700816
rect 213762 699514 213868 699530
rect 218808 699516 218836 703394
rect 218992 701010 219020 703520
rect 233884 703462 233936 703468
rect 218980 701004 219032 701010
rect 218980 700946 219032 700952
rect 223854 700224 223910 700233
rect 223854 700159 223910 700168
rect 223868 699516 223896 700159
rect 229008 699576 229060 699582
rect 228942 699524 229008 699530
rect 228942 699518 229060 699524
rect 213762 699508 213880 699514
rect 213762 699502 213828 699508
rect 228942 699502 229048 699518
rect 233896 699516 233924 703462
rect 235184 700942 235212 703520
rect 235172 700936 235224 700942
rect 235172 700878 235224 700884
rect 238956 699516 238984 703666
rect 249064 703588 249116 703594
rect 249064 703530 249116 703536
rect 244004 702296 244056 702302
rect 244004 702238 244056 702244
rect 244016 699516 244044 702238
rect 249076 699516 249104 703530
rect 251426 703520 251538 704960
rect 264152 703656 264204 703662
rect 264152 703598 264204 703604
rect 259184 701072 259236 701078
rect 259184 701014 259236 701020
rect 254124 700868 254176 700874
rect 254124 700810 254176 700816
rect 254136 699516 254164 700810
rect 259196 699516 259224 701014
rect 264164 699516 264192 703598
rect 267618 703520 267730 704960
rect 279332 703792 279384 703798
rect 279332 703734 279384 703740
rect 266360 701956 266412 701962
rect 266360 701898 266412 701904
rect 266372 700670 266400 701898
rect 266360 700664 266412 700670
rect 266360 700606 266412 700612
rect 267660 699786 267688 703520
rect 270684 702500 270736 702506
rect 270684 702442 270736 702448
rect 270696 700126 270724 702442
rect 270684 700120 270736 700126
rect 270684 700062 270736 700068
rect 274272 699984 274324 699990
rect 274272 699926 274324 699932
rect 269212 699916 269264 699922
rect 269212 699858 269264 699864
rect 267648 699780 267700 699786
rect 267648 699722 267700 699728
rect 269224 699516 269252 699858
rect 274284 699516 274312 699926
rect 279344 699516 279372 703734
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316040 703724 316092 703730
rect 316040 703666 316092 703672
rect 283852 700126 283880 703520
rect 286968 702228 287020 702234
rect 286968 702170 287020 702176
rect 284392 700664 284444 700670
rect 284392 700606 284444 700612
rect 283840 700120 283892 700126
rect 283840 700062 283892 700068
rect 284404 699516 284432 700606
rect 286980 700534 287008 702170
rect 300136 700534 300164 703520
rect 314660 702500 314712 702506
rect 314660 702442 314712 702448
rect 303528 701072 303580 701078
rect 303528 701014 303580 701020
rect 303540 700534 303568 701014
rect 309600 700936 309652 700942
rect 309600 700878 309652 700884
rect 286968 700528 287020 700534
rect 286968 700470 287020 700476
rect 294512 700528 294564 700534
rect 294512 700470 294564 700476
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 303528 700528 303580 700534
rect 303528 700470 303580 700476
rect 289452 699848 289504 699854
rect 289452 699790 289504 699796
rect 289464 699516 289492 699790
rect 294524 699516 294552 700470
rect 304540 700120 304592 700126
rect 304540 700062 304592 700068
rect 299480 699780 299532 699786
rect 299480 699722 299532 699728
rect 299492 699516 299520 699722
rect 304552 699516 304580 700062
rect 309612 699516 309640 700878
rect 314672 699516 314700 702442
rect 316052 700942 316080 703666
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 356060 703792 356112 703798
rect 356060 703734 356112 703740
rect 320824 702296 320876 702302
rect 320824 702238 320876 702244
rect 319720 701004 319772 701010
rect 319720 700946 319772 700952
rect 316040 700936 316092 700942
rect 316040 700878 316092 700884
rect 319732 699516 319760 700946
rect 320836 699786 320864 702238
rect 329840 702092 329892 702098
rect 329840 702034 329892 702040
rect 329852 700534 329880 702034
rect 332520 700670 332548 703520
rect 336556 702160 336608 702166
rect 336556 702102 336608 702108
rect 332600 702092 332652 702098
rect 332600 702034 332652 702040
rect 332508 700664 332560 700670
rect 332508 700606 332560 700612
rect 329840 700528 329892 700534
rect 329840 700470 329892 700476
rect 329748 700256 329800 700262
rect 329748 700198 329800 700204
rect 324780 700052 324832 700058
rect 324780 699994 324832 700000
rect 320824 699780 320876 699786
rect 320824 699722 320876 699728
rect 324792 699516 324820 699994
rect 329760 699516 329788 700198
rect 332612 699650 332640 702034
rect 336568 700670 336596 702102
rect 342076 702024 342128 702030
rect 342076 701966 342128 701972
rect 342088 700806 342116 701966
rect 339868 700800 339920 700806
rect 339868 700742 339920 700748
rect 342076 700800 342128 700806
rect 342076 700742 342128 700748
rect 336556 700664 336608 700670
rect 336556 700606 336608 700612
rect 334808 700188 334860 700194
rect 334808 700130 334860 700136
rect 332600 699644 332652 699650
rect 332600 699586 332652 699592
rect 334820 699516 334848 700130
rect 339880 699516 339908 700742
rect 344928 700596 344980 700602
rect 344928 700538 344980 700544
rect 344940 699516 344968 700538
rect 348804 699854 348832 703520
rect 356072 701010 356100 703734
rect 364248 703656 364300 703662
rect 364248 703598 364300 703604
rect 356060 701004 356112 701010
rect 356060 700946 356112 700952
rect 364260 700738 364288 703598
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 410432 703588 410484 703594
rect 410432 703530 410484 703536
rect 364996 701010 365024 703520
rect 370136 703384 370188 703390
rect 370136 703326 370188 703332
rect 364984 701004 365036 701010
rect 364984 700946 365036 700952
rect 349988 700732 350040 700738
rect 349988 700674 350040 700680
rect 364248 700732 364300 700738
rect 364248 700674 364300 700680
rect 348792 699848 348844 699854
rect 348792 699790 348844 699796
rect 350000 699516 350028 700674
rect 355048 700460 355100 700466
rect 355048 700402 355100 700408
rect 355060 699516 355088 700402
rect 365076 700392 365128 700398
rect 365076 700334 365128 700340
rect 360016 700324 360068 700330
rect 360016 700266 360068 700272
rect 360028 699516 360056 700266
rect 365088 699516 365116 700334
rect 370148 699516 370176 703326
rect 385316 703248 385368 703254
rect 385316 703190 385368 703196
rect 380256 702092 380308 702098
rect 380256 702034 380308 702040
rect 380268 699516 380296 702034
rect 385328 699516 385356 703190
rect 397472 699922 397500 703520
rect 400404 703112 400456 703118
rect 400404 703054 400456 703060
rect 397460 699916 397512 699922
rect 397460 699858 397512 699864
rect 400416 699516 400444 703054
rect 410444 700602 410472 703530
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 430028 703520 430080 703526
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 581644 703860 581696 703866
rect 581644 703802 581696 703808
rect 410524 702228 410576 702234
rect 410524 702170 410576 702176
rect 410432 700596 410484 700602
rect 410432 700538 410484 700544
rect 410536 699516 410564 702170
rect 413664 699990 413692 703520
rect 415584 702908 415636 702914
rect 415584 702850 415636 702856
rect 413652 699984 413704 699990
rect 413652 699926 413704 699932
rect 415596 699516 415624 702850
rect 429856 700738 429884 703520
rect 430028 703462 430080 703468
rect 430040 700738 430068 703462
rect 445852 702772 445904 702778
rect 445852 702714 445904 702720
rect 440792 701820 440844 701826
rect 440792 701762 440844 701768
rect 429844 700732 429896 700738
rect 429844 700674 429896 700680
rect 430028 700732 430080 700738
rect 430028 700674 430080 700680
rect 435732 699712 435784 699718
rect 435732 699654 435784 699660
rect 435744 699516 435772 699654
rect 440804 699516 440832 701762
rect 445864 699516 445892 702714
rect 462332 700874 462360 703520
rect 466000 701616 466052 701622
rect 466000 701558 466052 701564
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 466012 699516 466040 701558
rect 471060 701548 471112 701554
rect 471060 701490 471112 701496
rect 471072 699516 471100 701490
rect 478524 700126 478552 703520
rect 481180 701956 481232 701962
rect 481180 701898 481232 701904
rect 478512 700120 478564 700126
rect 478512 700062 478564 700068
rect 481192 699516 481220 701898
rect 486240 701412 486292 701418
rect 486240 701354 486292 701360
rect 486252 699516 486280 701354
rect 494808 700602 494836 703520
rect 526534 701448 526590 701457
rect 526534 701383 526590 701392
rect 501328 701208 501380 701214
rect 501328 701150 501380 701156
rect 494796 700596 494848 700602
rect 494796 700538 494848 700544
rect 501340 699516 501368 701150
rect 526548 699516 526576 701383
rect 527192 700942 527220 703520
rect 531594 701584 531650 701593
rect 531594 701519 531650 701528
rect 527180 700936 527232 700942
rect 527180 700878 527232 700884
rect 531608 699516 531636 701519
rect 543476 699786 543504 703520
rect 556802 701312 556858 701321
rect 556802 701247 556858 701256
rect 554780 701072 554832 701078
rect 554780 701014 554832 701020
rect 554792 700369 554820 701014
rect 554778 700360 554834 700369
rect 554778 700295 554834 700304
rect 543464 699780 543516 699786
rect 543464 699722 543516 699728
rect 556816 699516 556844 701247
rect 559668 700738 559696 703520
rect 581552 703452 581604 703458
rect 581552 703394 581604 703400
rect 561862 701720 561918 701729
rect 561862 701655 561918 701664
rect 559656 700732 559708 700738
rect 559656 700674 559708 700680
rect 561876 699516 561904 701655
rect 571984 701208 572036 701214
rect 571984 701150 572036 701156
rect 571996 699516 572024 701150
rect 577044 701072 577096 701078
rect 577044 701014 577096 701020
rect 577056 699516 577084 701014
rect 580540 700800 580592 700806
rect 580540 700742 580592 700748
rect 580446 699952 580502 699961
rect 580446 699887 580502 699896
rect 579988 699576 580040 699582
rect 579988 699518 580040 699524
rect 213828 699450 213880 699456
rect 144368 699440 144420 699446
rect 144368 699382 144420 699388
rect 208702 699378 208992 699394
rect 208702 699372 209004 699378
rect 208702 699366 208952 699372
rect 208952 699314 209004 699320
rect 579068 699372 579120 699378
rect 579068 699314 579120 699320
rect 374828 699304 374880 699310
rect 198674 699242 198780 699258
rect 374880 699252 375222 699258
rect 374828 699246 375222 699252
rect 198674 699236 198792 699242
rect 198674 699230 198740 699236
rect 374840 699230 375222 699246
rect 198740 699178 198792 699184
rect 395068 699168 395120 699174
rect 143354 699136 143410 699145
rect 143106 699094 143354 699122
rect 163594 699136 163650 699145
rect 163346 699094 163594 699122
rect 143354 699071 143410 699080
rect 193770 699136 193826 699145
rect 183494 699106 183600 699122
rect 183494 699100 183612 699106
rect 183494 699094 183560 699100
rect 163594 699071 163650 699080
rect 193614 699094 193770 699122
rect 193770 699071 193826 699080
rect 390098 699136 390154 699145
rect 390154 699094 390402 699122
rect 430762 699136 430818 699145
rect 395120 699116 395370 699122
rect 395068 699110 395370 699116
rect 395080 699094 395370 699110
rect 430698 699094 430762 699122
rect 390098 699071 390154 699080
rect 430762 699071 430818 699080
rect 450726 699136 450782 699145
rect 461030 699136 461086 699145
rect 450782 699094 450938 699122
rect 460966 699094 461030 699122
rect 450726 699071 450782 699080
rect 476210 699136 476266 699145
rect 476146 699094 476210 699122
rect 461030 699071 461086 699080
rect 476210 699071 476266 699080
rect 541346 699136 541402 699145
rect 541402 699094 541742 699122
rect 541346 699071 541402 699080
rect 183560 699042 183612 699048
rect 405188 699032 405240 699038
rect 17222 699000 17278 699009
rect 16974 698958 17222 698986
rect 112994 699000 113050 699009
rect 112838 698958 112994 698986
rect 17222 698935 17278 698944
rect 112994 698935 113050 698944
rect 132682 699000 132738 699009
rect 420276 699032 420328 699038
rect 405240 698980 405490 698986
rect 405188 698974 405490 698980
rect 425244 699032 425296 699038
rect 420328 698980 420670 698986
rect 420276 698974 420670 698980
rect 455604 699032 455656 699038
rect 425296 698980 425638 698986
rect 425244 698974 425638 698980
rect 490932 699032 490984 699038
rect 455656 698980 455906 698986
rect 455604 698974 455906 698980
rect 495900 699032 495952 699038
rect 490984 698980 491234 698986
rect 490932 698974 491234 698980
rect 506020 699032 506072 699038
rect 495952 698980 496294 698986
rect 495900 698974 496294 698980
rect 511172 699032 511224 699038
rect 506072 698980 506414 698986
rect 506020 698974 506414 698980
rect 516140 699032 516192 699038
rect 511224 698980 511474 698986
rect 511172 698974 511474 698980
rect 521108 699032 521160 699038
rect 516192 698980 516534 698986
rect 516140 698974 516534 698980
rect 536380 699032 536432 699038
rect 521160 698980 521502 698986
rect 521108 698974 521502 698980
rect 546500 699032 546552 699038
rect 536432 698980 536682 698986
rect 536380 698974 536682 698980
rect 551468 699032 551520 699038
rect 546552 698980 546802 698986
rect 546500 698974 546802 698980
rect 566556 699032 566608 699038
rect 551520 698980 551770 698986
rect 551468 698974 551770 698980
rect 566608 698980 566950 698986
rect 566556 698974 566950 698980
rect 405200 698958 405490 698974
rect 420288 698958 420670 698974
rect 425256 698958 425638 698974
rect 455616 698958 455906 698974
rect 490944 698958 491234 698974
rect 495912 698958 496294 698974
rect 506032 698958 506414 698974
rect 511184 698958 511474 698974
rect 516152 698958 516534 698974
rect 521120 698958 521502 698974
rect 536392 698958 536682 698974
rect 546512 698958 546802 698974
rect 551480 698958 551770 698974
rect 566568 698958 566950 698974
rect 132682 698935 132738 698944
rect 579080 654134 579108 699314
rect 579894 697232 579950 697241
rect 579894 697167 579950 697176
rect 579908 696969 579936 697167
rect 579894 696960 579950 696969
rect 579894 696895 579950 696904
rect 580000 683913 580028 699518
rect 580080 699508 580132 699514
rect 580080 699450 580132 699456
rect 579986 683904 580042 683913
rect 579986 683839 580042 683848
rect 579080 654106 579200 654134
rect 579172 644065 579200 654106
rect 579158 644056 579214 644065
rect 579158 643991 579214 644000
rect 580092 630873 580120 699450
rect 580356 699440 580408 699446
rect 580356 699382 580408 699388
rect 580172 699236 580224 699242
rect 580172 699178 580224 699184
rect 580078 630864 580134 630873
rect 580078 630799 580134 630808
rect 580184 577697 580212 699178
rect 580262 699000 580318 699009
rect 580262 698935 580318 698944
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 4858 358414 4936 358442
rect 4802 358391 4858 358400
rect 4632 357406 4844 357434
rect 4816 306270 4844 357406
rect 4804 306264 4856 306270
rect 4804 306206 4856 306212
rect 4066 293176 4122 293185
rect 4066 293111 4122 293120
rect 3974 201920 4030 201929
rect 3974 201855 4030 201864
rect 3882 188864 3938 188873
rect 3882 188799 3938 188808
rect 3790 149832 3846 149841
rect 3790 149767 3846 149776
rect 580276 59673 580304 698935
rect 580368 99521 580396 699382
rect 580460 139369 580488 699887
rect 580552 365129 580580 700742
rect 580816 700664 580868 700670
rect 580816 700606 580868 700612
rect 580724 700528 580776 700534
rect 580724 700470 580776 700476
rect 580630 700088 580686 700097
rect 580630 700023 580686 700032
rect 580538 365120 580594 365129
rect 580538 365055 580594 365064
rect 580644 258913 580672 700023
rect 580736 378457 580764 700470
rect 580828 471481 580856 700606
rect 580908 699100 580960 699106
rect 580908 699042 580960 699048
rect 580920 524521 580948 699042
rect 581564 670721 581592 703394
rect 581550 670712 581606 670721
rect 581550 670647 581606 670656
rect 580906 524512 580962 524521
rect 580906 524447 580962 524456
rect 580814 471472 580870 471481
rect 580814 471407 580870 471416
rect 580722 378448 580778 378457
rect 580722 378383 580778 378392
rect 580630 258904 580686 258913
rect 580630 258839 580686 258848
rect 580446 139360 580502 139369
rect 580446 139295 580502 139304
rect 580354 99512 580410 99521
rect 580354 99447 580410 99456
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 3698 45520 3754 45529
rect 3698 45455 3754 45464
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 581656 6633 581684 703802
rect 582288 703316 582340 703322
rect 582288 703258 582340 703264
rect 582196 703180 582248 703186
rect 582196 703122 582248 703128
rect 582104 702976 582156 702982
rect 582104 702918 582156 702924
rect 582012 702840 582064 702846
rect 582012 702782 582064 702788
rect 581736 702636 581788 702642
rect 581736 702578 581788 702584
rect 581748 46345 581776 702578
rect 581920 701344 581972 701350
rect 581920 701286 581972 701292
rect 581828 697740 581880 697746
rect 581828 697682 581880 697688
rect 581840 86193 581868 697682
rect 581932 219065 581960 701286
rect 582024 458153 582052 702782
rect 582116 511329 582144 702918
rect 582208 564369 582236 703122
rect 582300 617545 582328 703258
rect 582564 701208 582616 701214
rect 582564 701150 582616 701156
rect 582470 699816 582526 699825
rect 582470 699751 582526 699760
rect 582378 698320 582434 698329
rect 582378 698255 582434 698264
rect 582286 617536 582342 617545
rect 582286 617471 582342 617480
rect 582194 564360 582250 564369
rect 582194 564295 582250 564304
rect 582102 511320 582158 511329
rect 582102 511255 582158 511264
rect 582010 458144 582066 458153
rect 582010 458079 582066 458088
rect 581918 219056 581974 219065
rect 581918 218991 581974 219000
rect 581826 86184 581882 86193
rect 581826 86119 581882 86128
rect 581734 46336 581790 46345
rect 581734 46271 581790 46280
rect 582392 19825 582420 698255
rect 582484 73001 582512 699751
rect 582470 72992 582526 73001
rect 582470 72927 582526 72936
rect 582470 33144 582526 33153
rect 582470 33079 582472 33088
rect 582524 33079 582526 33088
rect 582472 33050 582524 33056
rect 582378 19816 582434 19825
rect 582378 19751 582434 19760
rect 581642 6624 581698 6633
rect 581642 6559 581698 6568
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3436 4146 3464 6423
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 572 2236 624 2242
rect 572 2178 624 2184
rect 584 480 612 2178
rect 1688 480 1716 2790
rect 2884 480 2912 2858
rect 4080 480 4108 2926
rect 5000 2242 5028 4420
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 4988 2236 5040 2242
rect 4988 2178 5040 2184
rect 5276 480 5304 2790
rect 6104 2786 6132 4420
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6092 2780 6144 2786
rect 6092 2722 6144 2728
rect 6472 480 6500 3538
rect 7300 2922 7328 4420
rect 8496 2990 8524 4420
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7668 480 7696 2790
rect 8772 480 8800 2926
rect 9600 2786 9628 4420
rect 10796 3602 10824 4420
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9588 2780 9640 2786
rect 9588 2722 9640 2728
rect 9968 480 9996 2994
rect 11164 480 11192 3062
rect 11992 2854 12020 4420
rect 13096 2990 13124 4420
rect 14292 3058 14320 4420
rect 15488 3126 15516 4420
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 12360 480 12388 2858
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13556 480 13584 2790
rect 14752 480 14780 2926
rect 15948 480 15976 3402
rect 16488 2916 16540 2922
rect 16592 2904 16620 4420
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 16540 2876 16620 2904
rect 16488 2858 16540 2864
rect 17052 480 17080 3062
rect 17788 2854 17816 4420
rect 18984 2990 19012 4420
rect 20088 3466 20116 4420
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 21284 3126 21312 4420
rect 21272 3120 21324 3126
rect 21272 3062 21324 3068
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18248 480 18276 2790
rect 19444 480 19472 2858
rect 20640 480 20668 2994
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21836 480 21864 2926
rect 22480 2854 22508 4420
rect 23584 2922 23612 4420
rect 24780 3058 24808 4420
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 24216 2916 24268 2922
rect 24216 2858 24268 2864
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 23032 480 23060 2790
rect 24228 480 24256 2858
rect 25332 480 25360 3470
rect 25976 2990 26004 4420
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 26516 2984 26568 2990
rect 26516 2926 26568 2932
rect 26528 480 26556 2926
rect 27080 2854 27108 4420
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 27724 480 27752 2994
rect 28276 2922 28304 4420
rect 29472 3534 29500 4420
rect 29460 3528 29512 3534
rect 29460 3470 29512 3476
rect 28908 3120 28960 3126
rect 28908 3062 28960 3068
rect 28264 2916 28316 2922
rect 28264 2858 28316 2864
rect 28920 480 28948 3062
rect 30576 2990 30604 4420
rect 31772 3058 31800 4420
rect 32968 3126 32996 4420
rect 32956 3120 33008 3126
rect 32956 3062 33008 3068
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 30564 2984 30616 2990
rect 30564 2926 30616 2932
rect 30104 2916 30156 2922
rect 30104 2858 30156 2864
rect 30116 480 30144 2858
rect 31300 2848 31352 2854
rect 31300 2790 31352 2796
rect 31312 480 31340 2790
rect 32416 480 32444 2994
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 33612 480 33640 2926
rect 34164 2922 34192 4420
rect 34796 3596 34848 3602
rect 34796 3538 34848 3544
rect 34152 2916 34204 2922
rect 34152 2858 34204 2864
rect 34808 480 34836 3538
rect 35268 2854 35296 4420
rect 35992 3120 36044 3126
rect 35992 3062 36044 3068
rect 35256 2848 35308 2854
rect 35256 2790 35308 2796
rect 36004 480 36032 3062
rect 36464 3058 36492 4420
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 37660 2990 37688 4420
rect 38764 3602 38792 4420
rect 38752 3596 38804 3602
rect 38752 3538 38804 3544
rect 39960 3126 39988 4420
rect 39948 3120 40000 3126
rect 39948 3062 40000 3068
rect 40684 3120 40736 3126
rect 40684 3062 40736 3068
rect 39580 3052 39632 3058
rect 39580 2994 39632 3000
rect 37648 2984 37700 2990
rect 37648 2926 37700 2932
rect 37188 2916 37240 2922
rect 37188 2858 37240 2864
rect 37200 480 37228 2858
rect 38384 2848 38436 2854
rect 38384 2790 38436 2796
rect 38396 480 38424 2790
rect 39592 480 39620 2994
rect 40696 480 40724 3062
rect 41156 2922 41184 4420
rect 41144 2916 41196 2922
rect 41144 2858 41196 2864
rect 41880 2916 41932 2922
rect 41880 2858 41932 2864
rect 41892 480 41920 2858
rect 42260 2854 42288 4420
rect 43456 3058 43484 4420
rect 44652 3126 44680 4420
rect 45468 3460 45520 3466
rect 45468 3402 45520 3408
rect 44640 3120 44692 3126
rect 44640 3062 44692 3068
rect 43444 3052 43496 3058
rect 43444 2994 43496 3000
rect 43076 2984 43128 2990
rect 43076 2926 43128 2932
rect 42248 2848 42300 2854
rect 42248 2790 42300 2796
rect 43088 480 43116 2926
rect 44272 2848 44324 2854
rect 44272 2790 44324 2796
rect 44284 480 44312 2790
rect 45480 480 45508 3402
rect 45756 2922 45784 4420
rect 46664 3188 46716 3194
rect 46664 3130 46716 3136
rect 45744 2916 45796 2922
rect 45744 2858 45796 2864
rect 46676 480 46704 3130
rect 46952 2990 46980 4420
rect 46940 2984 46992 2990
rect 46940 2926 46992 2932
rect 47860 2916 47912 2922
rect 47860 2858 47912 2864
rect 47872 480 47900 2858
rect 48148 2854 48176 4420
rect 49252 3466 49280 4420
rect 49240 3460 49292 3466
rect 49240 3402 49292 3408
rect 50448 3194 50476 4420
rect 50436 3188 50488 3194
rect 50436 3130 50488 3136
rect 50160 3120 50212 3126
rect 50160 3062 50212 3068
rect 48964 3052 49016 3058
rect 48964 2994 49016 3000
rect 48136 2848 48188 2854
rect 48136 2790 48188 2796
rect 48976 480 49004 2994
rect 50172 480 50200 3062
rect 51356 2984 51408 2990
rect 51356 2926 51408 2932
rect 51368 480 51396 2926
rect 51644 2922 51672 4420
rect 52748 3058 52776 4420
rect 53944 3126 53972 4420
rect 54944 3596 54996 3602
rect 54944 3538 54996 3544
rect 53932 3120 53984 3126
rect 53932 3062 53984 3068
rect 52736 3052 52788 3058
rect 52736 2994 52788 3000
rect 51632 2916 51684 2922
rect 51632 2858 51684 2864
rect 53748 2916 53800 2922
rect 53748 2858 53800 2864
rect 52552 2848 52604 2854
rect 52552 2790 52604 2796
rect 52564 480 52592 2790
rect 53760 480 53788 2858
rect 54956 480 54984 3538
rect 55140 2990 55168 4420
rect 55128 2984 55180 2990
rect 55128 2926 55180 2932
rect 56048 2984 56100 2990
rect 56048 2926 56100 2932
rect 56060 480 56088 2926
rect 56244 2854 56272 4420
rect 57440 2922 57468 4420
rect 58636 3602 58664 4420
rect 58624 3596 58676 3602
rect 58624 3538 58676 3544
rect 59636 3052 59688 3058
rect 59636 2994 59688 3000
rect 57428 2916 57480 2922
rect 57428 2858 57480 2864
rect 58440 2916 58492 2922
rect 58440 2858 58492 2864
rect 56232 2848 56284 2854
rect 56232 2790 56284 2796
rect 57244 2848 57296 2854
rect 57244 2790 57296 2796
rect 57256 480 57284 2790
rect 58452 480 58480 2858
rect 59648 480 59676 2994
rect 59832 2990 59860 4420
rect 59820 2984 59872 2990
rect 59820 2926 59872 2932
rect 60832 2984 60884 2990
rect 60832 2926 60884 2932
rect 60844 480 60872 2926
rect 60936 2854 60964 4420
rect 62132 2922 62160 4420
rect 63328 3058 63356 4420
rect 64328 3460 64380 3466
rect 64328 3402 64380 3408
rect 63316 3052 63368 3058
rect 63316 2994 63368 3000
rect 62120 2916 62172 2922
rect 62120 2858 62172 2864
rect 63224 2916 63276 2922
rect 63224 2858 63276 2864
rect 60924 2848 60976 2854
rect 60924 2790 60976 2796
rect 62028 2848 62080 2854
rect 62028 2790 62080 2796
rect 62040 480 62068 2790
rect 63236 480 63264 2858
rect 64340 480 64368 3402
rect 64432 2990 64460 4420
rect 65524 3188 65576 3194
rect 65524 3130 65576 3136
rect 64420 2984 64472 2990
rect 64420 2926 64472 2932
rect 65536 480 65564 3130
rect 65628 2854 65656 4420
rect 66720 3732 66772 3738
rect 66720 3674 66772 3680
rect 65616 2848 65668 2854
rect 65616 2790 65668 2796
rect 66732 480 66760 3674
rect 66824 2922 66852 4420
rect 67928 3466 67956 4420
rect 67916 3460 67968 3466
rect 67916 3402 67968 3408
rect 69124 3194 69152 4420
rect 70320 3738 70348 4420
rect 70308 3732 70360 3738
rect 70308 3674 70360 3680
rect 70308 3596 70360 3602
rect 70308 3538 70360 3544
rect 69112 3188 69164 3194
rect 69112 3130 69164 3136
rect 69112 3052 69164 3058
rect 69112 2994 69164 3000
rect 66812 2916 66864 2922
rect 66812 2858 66864 2864
rect 67916 2848 67968 2854
rect 67916 2790 67968 2796
rect 67928 480 67956 2790
rect 69124 480 69152 2994
rect 70320 480 70348 3538
rect 71424 2854 71452 4420
rect 72620 3058 72648 4420
rect 73816 3602 73844 4420
rect 73804 3596 73856 3602
rect 73804 3538 73856 3544
rect 73804 3460 73856 3466
rect 73804 3402 73856 3408
rect 72608 3052 72660 3058
rect 72608 2994 72660 3000
rect 72608 2916 72660 2922
rect 72608 2858 72660 2864
rect 71412 2848 71464 2854
rect 71412 2790 71464 2796
rect 71504 2848 71556 2854
rect 71504 2790 71556 2796
rect 71516 480 71544 2790
rect 72620 480 72648 2858
rect 73816 480 73844 3402
rect 74920 2854 74948 4420
rect 76116 2922 76144 4420
rect 77312 3466 77340 4420
rect 77300 3460 77352 3466
rect 77300 3402 77352 3408
rect 77392 2984 77444 2990
rect 77392 2926 77444 2932
rect 76104 2916 76156 2922
rect 76104 2858 76156 2864
rect 76196 2916 76248 2922
rect 76196 2858 76248 2864
rect 74908 2848 74960 2854
rect 74908 2790 74960 2796
rect 75000 2848 75052 2854
rect 75000 2790 75052 2796
rect 75012 480 75040 2790
rect 76208 480 76236 2858
rect 77404 480 77432 2926
rect 78416 2854 78444 4420
rect 79612 2922 79640 4420
rect 80808 2990 80836 4420
rect 80796 2984 80848 2990
rect 80796 2926 80848 2932
rect 80888 2984 80940 2990
rect 80888 2926 80940 2932
rect 79600 2916 79652 2922
rect 79600 2858 79652 2864
rect 79692 2916 79744 2922
rect 79692 2858 79744 2864
rect 78404 2848 78456 2854
rect 78404 2790 78456 2796
rect 78588 2848 78640 2854
rect 78588 2790 78640 2796
rect 78600 480 78628 2790
rect 79704 480 79732 2858
rect 80900 480 80928 2926
rect 81912 2854 81940 4420
rect 82084 3052 82136 3058
rect 82084 2994 82136 3000
rect 81900 2848 81952 2854
rect 81900 2790 81952 2796
rect 82096 480 82124 2994
rect 83108 2922 83136 4420
rect 84304 2990 84332 4420
rect 85500 3058 85528 4420
rect 85488 3052 85540 3058
rect 85488 2994 85540 3000
rect 84292 2984 84344 2990
rect 84292 2926 84344 2932
rect 85672 2984 85724 2990
rect 85672 2926 85724 2932
rect 83096 2916 83148 2922
rect 83096 2858 83148 2864
rect 84476 2916 84528 2922
rect 84476 2858 84528 2864
rect 83280 2848 83332 2854
rect 83280 2790 83332 2796
rect 83292 480 83320 2790
rect 84488 480 84516 2858
rect 85684 480 85712 2926
rect 86604 2854 86632 4420
rect 87800 2922 87828 4420
rect 88996 2990 89024 4420
rect 88984 2984 89036 2990
rect 88984 2926 89036 2932
rect 89168 2984 89220 2990
rect 89168 2926 89220 2932
rect 87788 2916 87840 2922
rect 87788 2858 87840 2864
rect 87972 2916 88024 2922
rect 87972 2858 88024 2864
rect 86592 2848 86644 2854
rect 86592 2790 86644 2796
rect 86868 2848 86920 2854
rect 86868 2790 86920 2796
rect 86880 480 86908 2790
rect 87984 480 88012 2858
rect 89180 480 89208 2926
rect 90100 2854 90128 4420
rect 91296 2922 91324 4420
rect 92492 2990 92520 4420
rect 92480 2984 92532 2990
rect 92480 2926 92532 2932
rect 92756 2984 92808 2990
rect 92756 2926 92808 2932
rect 91284 2916 91336 2922
rect 91284 2858 91336 2864
rect 91560 2916 91612 2922
rect 91560 2858 91612 2864
rect 90088 2848 90140 2854
rect 90088 2790 90140 2796
rect 90364 2848 90416 2854
rect 90364 2790 90416 2796
rect 90376 480 90404 2790
rect 91572 480 91600 2858
rect 92768 480 92796 2926
rect 93596 2854 93624 4420
rect 94792 2922 94820 4420
rect 95988 2990 96016 4420
rect 95976 2984 96028 2990
rect 95976 2926 96028 2932
rect 96252 2984 96304 2990
rect 96252 2926 96304 2932
rect 94780 2916 94832 2922
rect 94780 2858 94832 2864
rect 95148 2916 95200 2922
rect 95148 2858 95200 2864
rect 93584 2848 93636 2854
rect 93584 2790 93636 2796
rect 93952 2848 94004 2854
rect 93952 2790 94004 2796
rect 93964 480 93992 2790
rect 95160 480 95188 2858
rect 96264 480 96292 2926
rect 97092 2854 97120 4420
rect 98288 2922 98316 4420
rect 99484 2990 99512 4420
rect 99472 2984 99524 2990
rect 99472 2926 99524 2932
rect 99840 2984 99892 2990
rect 99840 2926 99892 2932
rect 98276 2916 98328 2922
rect 98276 2858 98328 2864
rect 98644 2916 98696 2922
rect 98644 2858 98696 2864
rect 97080 2848 97132 2854
rect 97080 2790 97132 2796
rect 97448 2848 97500 2854
rect 97448 2790 97500 2796
rect 97460 480 97488 2790
rect 98656 480 98684 2858
rect 99852 480 99880 2926
rect 100588 2854 100616 4420
rect 101784 2922 101812 4420
rect 102980 2990 103008 4420
rect 103336 3460 103388 3466
rect 103336 3402 103388 3408
rect 102968 2984 103020 2990
rect 102968 2926 103020 2932
rect 101772 2916 101824 2922
rect 101772 2858 101824 2864
rect 102232 2916 102284 2922
rect 102232 2858 102284 2864
rect 100576 2848 100628 2854
rect 100576 2790 100628 2796
rect 101036 2848 101088 2854
rect 101036 2790 101088 2796
rect 101048 480 101076 2790
rect 102244 480 102272 2858
rect 103348 480 103376 3402
rect 104084 2854 104112 4420
rect 105280 2922 105308 4420
rect 106476 3466 106504 4420
rect 106464 3460 106516 3466
rect 106464 3402 106516 3408
rect 106924 3052 106976 3058
rect 106924 2994 106976 3000
rect 105268 2916 105320 2922
rect 105268 2858 105320 2864
rect 105728 2916 105780 2922
rect 105728 2858 105780 2864
rect 104072 2848 104124 2854
rect 104072 2790 104124 2796
rect 104532 2848 104584 2854
rect 104532 2790 104584 2796
rect 104544 480 104572 2790
rect 105740 480 105768 2858
rect 106936 480 106964 2994
rect 107580 2854 107608 4420
rect 108120 2984 108172 2990
rect 108120 2926 108172 2932
rect 107568 2848 107620 2854
rect 107568 2790 107620 2796
rect 108132 480 108160 2926
rect 108776 2922 108804 4420
rect 109972 3058 110000 4420
rect 109960 3052 110012 3058
rect 109960 2994 110012 3000
rect 111168 2990 111196 4420
rect 111156 2984 111208 2990
rect 111156 2926 111208 2932
rect 111616 2984 111668 2990
rect 111616 2926 111668 2932
rect 108764 2916 108816 2922
rect 108764 2858 108816 2864
rect 110512 2916 110564 2922
rect 110512 2858 110564 2864
rect 109316 2848 109368 2854
rect 109316 2790 109368 2796
rect 109328 480 109356 2790
rect 110524 480 110552 2858
rect 111628 480 111656 2926
rect 112272 2854 112300 4420
rect 113468 2922 113496 4420
rect 114008 3052 114060 3058
rect 114008 2994 114060 3000
rect 113456 2916 113508 2922
rect 113456 2858 113508 2864
rect 112260 2848 112312 2854
rect 112260 2790 112312 2796
rect 112812 2848 112864 2854
rect 112812 2790 112864 2796
rect 112824 480 112852 2790
rect 114020 480 114048 2994
rect 114664 2990 114692 4420
rect 114652 2984 114704 2990
rect 114652 2926 114704 2932
rect 115768 2922 115796 4420
rect 116964 3058 116992 4420
rect 116952 3052 117004 3058
rect 116952 2994 117004 3000
rect 117596 2984 117648 2990
rect 117596 2926 117648 2932
rect 115756 2916 115808 2922
rect 115756 2858 115808 2864
rect 116400 2916 116452 2922
rect 116400 2858 116452 2864
rect 115204 2848 115256 2854
rect 115204 2790 115256 2796
rect 115216 480 115244 2790
rect 116412 480 116440 2858
rect 117608 480 117636 2926
rect 118160 2854 118188 4420
rect 119264 2922 119292 4420
rect 120460 2990 120488 4420
rect 120448 2984 120500 2990
rect 120448 2926 120500 2932
rect 121092 2984 121144 2990
rect 121092 2926 121144 2932
rect 119252 2916 119304 2922
rect 119252 2858 119304 2864
rect 119896 2916 119948 2922
rect 119896 2858 119948 2864
rect 118148 2848 118200 2854
rect 118148 2790 118200 2796
rect 118792 2848 118844 2854
rect 118792 2790 118844 2796
rect 118804 480 118832 2790
rect 119908 480 119936 2858
rect 121104 480 121132 2926
rect 121656 2854 121684 4420
rect 122760 2922 122788 4420
rect 123956 2990 123984 4420
rect 123944 2984 123996 2990
rect 123944 2926 123996 2932
rect 124680 2984 124732 2990
rect 124680 2926 124732 2932
rect 122748 2916 122800 2922
rect 122748 2858 122800 2864
rect 123484 2916 123536 2922
rect 123484 2858 123536 2864
rect 121644 2848 121696 2854
rect 121644 2790 121696 2796
rect 122288 2848 122340 2854
rect 122288 2790 122340 2796
rect 122300 480 122328 2790
rect 123496 480 123524 2858
rect 124692 480 124720 2926
rect 125152 2854 125180 4420
rect 126256 2922 126284 4420
rect 127452 2990 127480 4420
rect 128176 3052 128228 3058
rect 128176 2994 128228 3000
rect 127440 2984 127492 2990
rect 127440 2926 127492 2932
rect 126244 2916 126296 2922
rect 126244 2858 126296 2864
rect 126980 2916 127032 2922
rect 126980 2858 127032 2864
rect 125140 2848 125192 2854
rect 125140 2790 125192 2796
rect 125876 2848 125928 2854
rect 125876 2790 125928 2796
rect 125888 480 125916 2790
rect 126992 480 127020 2858
rect 128188 480 128216 2994
rect 128648 2854 128676 4420
rect 129372 2984 129424 2990
rect 129372 2926 129424 2932
rect 128636 2848 128688 2854
rect 128636 2790 128688 2796
rect 129384 480 129412 2926
rect 129752 2922 129780 4420
rect 130948 3058 130976 4420
rect 130936 3052 130988 3058
rect 130936 2994 130988 3000
rect 132144 2990 132172 4420
rect 132132 2984 132184 2990
rect 132132 2926 132184 2932
rect 132960 2984 133012 2990
rect 132960 2926 133012 2932
rect 129740 2916 129792 2922
rect 129740 2858 129792 2864
rect 131764 2916 131816 2922
rect 131764 2858 131816 2864
rect 130568 2848 130620 2854
rect 130568 2790 130620 2796
rect 130580 480 130608 2790
rect 131776 480 131804 2858
rect 132972 480 133000 2926
rect 133248 2854 133276 4420
rect 134156 3052 134208 3058
rect 134156 2994 134208 3000
rect 133236 2848 133288 2854
rect 133236 2790 133288 2796
rect 134168 480 134196 2994
rect 134444 2922 134472 4420
rect 135260 3120 135312 3126
rect 135260 3062 135312 3068
rect 134432 2916 134484 2922
rect 134432 2858 134484 2864
rect 135272 480 135300 3062
rect 135640 2990 135668 4420
rect 136836 3058 136864 4420
rect 137940 3126 137968 4420
rect 137928 3120 137980 3126
rect 137928 3062 137980 3068
rect 136824 3052 136876 3058
rect 136824 2994 136876 3000
rect 135628 2984 135680 2990
rect 135628 2926 135680 2932
rect 138848 2984 138900 2990
rect 138848 2926 138900 2932
rect 137652 2916 137704 2922
rect 137652 2858 137704 2864
rect 136456 2848 136508 2854
rect 136456 2790 136508 2796
rect 136468 480 136496 2790
rect 137664 480 137692 2858
rect 138860 480 138888 2926
rect 139136 2854 139164 4420
rect 140332 2922 140360 4420
rect 141436 2990 141464 4420
rect 141424 2984 141476 2990
rect 141424 2926 141476 2932
rect 142436 2984 142488 2990
rect 142436 2926 142488 2932
rect 140320 2916 140372 2922
rect 140320 2858 140372 2864
rect 141240 2916 141292 2922
rect 141240 2858 141292 2864
rect 139124 2848 139176 2854
rect 139124 2790 139176 2796
rect 140044 2848 140096 2854
rect 140044 2790 140096 2796
rect 140056 480 140084 2790
rect 141252 480 141280 2858
rect 142448 480 142476 2926
rect 142632 2854 142660 4420
rect 143540 3052 143592 3058
rect 143540 2994 143592 3000
rect 142620 2848 142672 2854
rect 142620 2790 142672 2796
rect 143552 480 143580 2994
rect 143828 2922 143856 4420
rect 144736 3120 144788 3126
rect 144736 3062 144788 3068
rect 143816 2916 143868 2922
rect 143816 2858 143868 2864
rect 144748 480 144776 3062
rect 144932 2990 144960 4420
rect 146128 3058 146156 4420
rect 147324 3126 147352 4420
rect 147312 3120 147364 3126
rect 147312 3062 147364 3068
rect 146116 3052 146168 3058
rect 146116 2994 146168 3000
rect 144920 2984 144972 2990
rect 144920 2926 144972 2932
rect 148324 2984 148376 2990
rect 148324 2926 148376 2932
rect 147128 2916 147180 2922
rect 147128 2858 147180 2864
rect 145932 2848 145984 2854
rect 145932 2790 145984 2796
rect 145944 480 145972 2790
rect 147140 480 147168 2858
rect 148336 480 148364 2926
rect 148428 2854 148456 4420
rect 149624 2922 149652 4420
rect 150820 2990 150848 4420
rect 151820 3052 151872 3058
rect 151820 2994 151872 3000
rect 150808 2984 150860 2990
rect 150808 2926 150860 2932
rect 149612 2916 149664 2922
rect 149612 2858 149664 2864
rect 150624 2916 150676 2922
rect 150624 2858 150676 2864
rect 148416 2848 148468 2854
rect 148416 2790 148468 2796
rect 149520 2848 149572 2854
rect 149520 2790 149572 2796
rect 149532 480 149560 2790
rect 150636 480 150664 2858
rect 151832 480 151860 2994
rect 151924 2854 151952 4420
rect 153016 4072 153068 4078
rect 153016 4014 153068 4020
rect 151912 2848 151964 2854
rect 151912 2790 151964 2796
rect 153028 480 153056 4014
rect 153120 2922 153148 4420
rect 154316 3058 154344 4420
rect 155420 4078 155448 4420
rect 155408 4072 155460 4078
rect 155408 4014 155460 4020
rect 155408 3936 155460 3942
rect 155408 3878 155460 3884
rect 154304 3052 154356 3058
rect 154304 2994 154356 3000
rect 154212 2984 154264 2990
rect 154212 2926 154264 2932
rect 153108 2916 153160 2922
rect 153108 2858 153160 2864
rect 154224 480 154252 2926
rect 155420 480 155448 3878
rect 156616 2990 156644 4420
rect 157812 3942 157840 4420
rect 157800 3936 157852 3942
rect 157800 3878 157852 3884
rect 157800 3800 157852 3806
rect 157800 3742 157852 3748
rect 156604 2984 156656 2990
rect 156604 2926 156656 2932
rect 156604 2848 156656 2854
rect 156604 2790 156656 2796
rect 156616 480 156644 2790
rect 157812 480 157840 3742
rect 158916 2854 158944 4420
rect 160112 3806 160140 4420
rect 160100 3800 160152 3806
rect 160100 3742 160152 3748
rect 160100 3664 160152 3670
rect 160100 3606 160152 3612
rect 158996 2984 159048 2990
rect 158996 2926 159048 2932
rect 158904 2848 158956 2854
rect 158904 2790 158956 2796
rect 159008 2258 159036 2926
rect 158916 2230 159036 2258
rect 158916 480 158944 2230
rect 160112 480 160140 3606
rect 161308 2990 161336 4420
rect 162504 3670 162532 4420
rect 162492 3664 162544 3670
rect 162492 3606 162544 3612
rect 161296 2984 161348 2990
rect 161296 2926 161348 2932
rect 162492 2984 162544 2990
rect 162492 2926 162544 2932
rect 161296 2848 161348 2854
rect 161296 2790 161348 2796
rect 161308 480 161336 2790
rect 162504 480 162532 2926
rect 163608 2854 163636 4420
rect 164804 2990 164832 4420
rect 164792 2984 164844 2990
rect 164792 2926 164844 2932
rect 166000 2922 166028 4420
rect 163688 2916 163740 2922
rect 163688 2858 163740 2864
rect 165988 2916 166040 2922
rect 165988 2858 166040 2864
rect 166080 2916 166132 2922
rect 166080 2858 166132 2864
rect 163596 2848 163648 2854
rect 163596 2790 163648 2796
rect 163700 480 163728 2858
rect 164884 2848 164936 2854
rect 164884 2790 164936 2796
rect 164896 480 164924 2790
rect 166092 480 166120 2858
rect 167104 2854 167132 4420
rect 167184 2984 167236 2990
rect 167184 2926 167236 2932
rect 167092 2848 167144 2854
rect 167092 2790 167144 2796
rect 167196 480 167224 2926
rect 168300 2922 168328 4420
rect 169496 2990 169524 4420
rect 169484 2984 169536 2990
rect 169484 2926 169536 2932
rect 168288 2916 168340 2922
rect 168288 2858 168340 2864
rect 169576 2916 169628 2922
rect 169576 2858 169628 2864
rect 168380 2848 168432 2854
rect 168380 2790 168432 2796
rect 168392 480 168420 2790
rect 169588 480 169616 2858
rect 170600 2854 170628 4420
rect 171796 2922 171824 4420
rect 172992 2922 173020 4420
rect 171784 2916 171836 2922
rect 171784 2858 171836 2864
rect 172980 2916 173032 2922
rect 172980 2858 173032 2864
rect 173164 2916 173216 2922
rect 173164 2858 173216 2864
rect 170588 2848 170640 2854
rect 170588 2790 170640 2796
rect 170772 2848 170824 2854
rect 170772 2790 170824 2796
rect 171968 2848 172020 2854
rect 171968 2790 172020 2796
rect 170784 480 170812 2790
rect 171980 480 172008 2790
rect 173176 480 173204 2858
rect 174096 2854 174124 4420
rect 174268 2984 174320 2990
rect 174268 2926 174320 2932
rect 174084 2848 174136 2854
rect 174084 2790 174136 2796
rect 174280 480 174308 2926
rect 175292 2922 175320 4420
rect 176488 2990 176516 4420
rect 176476 2984 176528 2990
rect 176476 2926 176528 2932
rect 175280 2916 175332 2922
rect 175280 2858 175332 2864
rect 176660 2916 176712 2922
rect 176660 2858 176712 2864
rect 175464 2848 175516 2854
rect 175464 2790 175516 2796
rect 175476 480 175504 2790
rect 176672 480 176700 2858
rect 177592 2854 177620 4420
rect 177856 2984 177908 2990
rect 177856 2926 177908 2932
rect 177580 2848 177632 2854
rect 177580 2790 177632 2796
rect 177868 480 177896 2926
rect 178788 2922 178816 4420
rect 179984 2990 180012 4420
rect 179972 2984 180024 2990
rect 179972 2926 180024 2932
rect 178776 2916 178828 2922
rect 178776 2858 178828 2864
rect 180248 2916 180300 2922
rect 180248 2858 180300 2864
rect 179052 2848 179104 2854
rect 179052 2790 179104 2796
rect 179064 480 179092 2790
rect 180260 480 180288 2858
rect 181088 2854 181116 4420
rect 181444 2984 181496 2990
rect 181444 2926 181496 2932
rect 181076 2848 181128 2854
rect 181076 2790 181128 2796
rect 181456 480 181484 2926
rect 182284 2922 182312 4420
rect 183480 2990 183508 4420
rect 183468 2984 183520 2990
rect 183468 2926 183520 2932
rect 182272 2916 182324 2922
rect 182272 2858 182324 2864
rect 183744 2916 183796 2922
rect 183744 2858 183796 2864
rect 182548 2848 182600 2854
rect 182548 2790 182600 2796
rect 182560 480 182588 2790
rect 183756 480 183784 2858
rect 184584 2854 184612 4420
rect 185780 2922 185808 4420
rect 185768 2916 185820 2922
rect 185768 2858 185820 2864
rect 186136 2916 186188 2922
rect 186136 2858 186188 2864
rect 184572 2848 184624 2854
rect 184572 2790 184624 2796
rect 184940 2848 184992 2854
rect 184940 2790 184992 2796
rect 184952 480 184980 2790
rect 186148 480 186176 2858
rect 186976 2854 187004 4420
rect 188172 2922 188200 4420
rect 188160 2916 188212 2922
rect 188160 2858 188212 2864
rect 188528 2916 188580 2922
rect 188528 2858 188580 2864
rect 186964 2848 187016 2854
rect 186964 2790 187016 2796
rect 187332 2848 187384 2854
rect 187332 2790 187384 2796
rect 187344 480 187372 2790
rect 188540 480 188568 2858
rect 189276 2854 189304 4420
rect 190472 2922 190500 4420
rect 191668 2922 191696 4420
rect 192024 2984 192076 2990
rect 192024 2926 192076 2932
rect 190460 2916 190512 2922
rect 190460 2858 190512 2864
rect 191656 2916 191708 2922
rect 191656 2858 191708 2864
rect 189264 2848 189316 2854
rect 189264 2790 189316 2796
rect 189724 2848 189776 2854
rect 189724 2790 189776 2796
rect 190828 2848 190880 2854
rect 190828 2790 190880 2796
rect 189736 480 189764 2790
rect 190840 480 190868 2790
rect 192036 480 192064 2926
rect 192772 2854 192800 4420
rect 193968 2990 193996 4420
rect 193956 2984 194008 2990
rect 193956 2926 194008 2932
rect 195164 2922 195192 4420
rect 193220 2916 193272 2922
rect 193220 2858 193272 2864
rect 195152 2916 195204 2922
rect 195152 2858 195204 2864
rect 195612 2916 195664 2922
rect 195612 2858 195664 2864
rect 192760 2848 192812 2854
rect 192760 2790 192812 2796
rect 193232 480 193260 2858
rect 194416 2848 194468 2854
rect 194416 2790 194468 2796
rect 194428 480 194456 2790
rect 195624 480 195652 2858
rect 196268 2854 196296 4420
rect 197464 2922 197492 4420
rect 197452 2916 197504 2922
rect 197452 2858 197504 2864
rect 197912 2916 197964 2922
rect 197912 2858 197964 2864
rect 196256 2848 196308 2854
rect 196256 2790 196308 2796
rect 196808 2848 196860 2854
rect 196808 2790 196860 2796
rect 196820 480 196848 2790
rect 197924 480 197952 2858
rect 198660 2854 198688 4420
rect 199108 2984 199160 2990
rect 199108 2926 199160 2932
rect 198648 2848 198700 2854
rect 198648 2790 198700 2796
rect 199120 480 199148 2926
rect 199764 2922 199792 4420
rect 200960 2990 200988 4420
rect 200948 2984 201000 2990
rect 200948 2926 201000 2932
rect 202156 2922 202184 4420
rect 202696 2984 202748 2990
rect 202696 2926 202748 2932
rect 199752 2916 199804 2922
rect 199752 2858 199804 2864
rect 200304 2916 200356 2922
rect 200304 2858 200356 2864
rect 202144 2916 202196 2922
rect 202144 2858 202196 2864
rect 200316 480 200344 2858
rect 201500 2848 201552 2854
rect 201500 2790 201552 2796
rect 201512 480 201540 2790
rect 202708 480 202736 2926
rect 203260 2854 203288 4420
rect 204456 2990 204484 4420
rect 204444 2984 204496 2990
rect 204444 2926 204496 2932
rect 205652 2922 205680 4420
rect 206192 2984 206244 2990
rect 206192 2926 206244 2932
rect 203892 2916 203944 2922
rect 203892 2858 203944 2864
rect 205640 2916 205692 2922
rect 205640 2858 205692 2864
rect 203248 2848 203300 2854
rect 203248 2790 203300 2796
rect 203904 480 203932 2858
rect 205088 2848 205140 2854
rect 205088 2790 205140 2796
rect 205100 480 205128 2790
rect 206204 480 206232 2926
rect 206756 2854 206784 4420
rect 207952 2990 207980 4420
rect 207940 2984 207992 2990
rect 207940 2926 207992 2932
rect 209148 2922 209176 4420
rect 209780 2984 209832 2990
rect 209780 2926 209832 2932
rect 207388 2916 207440 2922
rect 207388 2858 207440 2864
rect 209136 2916 209188 2922
rect 209136 2858 209188 2864
rect 206744 2848 206796 2854
rect 206744 2790 206796 2796
rect 207400 480 207428 2858
rect 208584 2848 208636 2854
rect 208584 2790 208636 2796
rect 208596 480 208624 2790
rect 209792 480 209820 2926
rect 210252 2854 210280 4420
rect 211448 2990 211476 4420
rect 211436 2984 211488 2990
rect 211436 2926 211488 2932
rect 212644 2922 212672 4420
rect 210976 2916 211028 2922
rect 210976 2858 211028 2864
rect 212632 2916 212684 2922
rect 212632 2858 212684 2864
rect 213368 2916 213420 2922
rect 213368 2858 213420 2864
rect 210240 2848 210292 2854
rect 210240 2790 210292 2796
rect 210988 480 211016 2858
rect 212172 2848 212224 2854
rect 212172 2790 212224 2796
rect 212184 480 212212 2790
rect 213380 480 213408 2858
rect 213748 2854 213776 4420
rect 214944 2922 214972 4420
rect 215668 2984 215720 2990
rect 215668 2926 215720 2932
rect 214932 2916 214984 2922
rect 214932 2858 214984 2864
rect 213736 2848 213788 2854
rect 213736 2790 213788 2796
rect 214472 2848 214524 2854
rect 214472 2790 214524 2796
rect 214484 480 214512 2790
rect 215680 480 215708 2926
rect 216140 2854 216168 4420
rect 217336 2990 217364 4420
rect 217324 2984 217376 2990
rect 217324 2926 217376 2932
rect 218440 2922 218468 4420
rect 216864 2916 216916 2922
rect 216864 2858 216916 2864
rect 218428 2916 218480 2922
rect 218428 2858 218480 2864
rect 219256 2916 219308 2922
rect 219256 2858 219308 2864
rect 216128 2848 216180 2854
rect 216128 2790 216180 2796
rect 216876 480 216904 2858
rect 218060 2848 218112 2854
rect 218060 2790 218112 2796
rect 218072 480 218100 2790
rect 219268 480 219296 2858
rect 219636 2854 219664 4420
rect 220832 2922 220860 4420
rect 220820 2916 220872 2922
rect 220820 2858 220872 2864
rect 221556 2916 221608 2922
rect 221556 2858 221608 2864
rect 219624 2848 219676 2854
rect 219624 2790 219676 2796
rect 220452 2848 220504 2854
rect 220452 2790 220504 2796
rect 220464 480 220492 2790
rect 221568 480 221596 2858
rect 221936 2854 221964 4420
rect 223132 2922 223160 4420
rect 223120 2916 223172 2922
rect 223120 2858 223172 2864
rect 223948 2916 224000 2922
rect 223948 2858 224000 2864
rect 221924 2848 221976 2854
rect 221924 2790 221976 2796
rect 222752 2848 222804 2854
rect 222752 2790 222804 2796
rect 222764 480 222792 2790
rect 223960 480 223988 2858
rect 224328 2854 224356 4420
rect 225432 2922 225460 4420
rect 226340 2984 226392 2990
rect 226340 2926 226392 2932
rect 225420 2916 225472 2922
rect 225420 2858 225472 2864
rect 224316 2848 224368 2854
rect 224316 2790 224368 2796
rect 225144 2848 225196 2854
rect 225144 2790 225196 2796
rect 225156 480 225184 2790
rect 226352 480 226380 2926
rect 226628 2854 226656 4420
rect 227824 2990 227852 4420
rect 227812 2984 227864 2990
rect 227812 2926 227864 2932
rect 228928 2922 228956 4420
rect 229836 2984 229888 2990
rect 229836 2926 229888 2932
rect 227536 2916 227588 2922
rect 227536 2858 227588 2864
rect 228916 2916 228968 2922
rect 228916 2858 228968 2864
rect 226616 2848 226668 2854
rect 226616 2790 226668 2796
rect 227548 480 227576 2858
rect 228732 2848 228784 2854
rect 228732 2790 228784 2796
rect 228744 480 228772 2790
rect 229848 480 229876 2926
rect 230124 2854 230152 4420
rect 231320 2990 231348 4420
rect 231308 2984 231360 2990
rect 231308 2926 231360 2932
rect 232424 2922 232452 4420
rect 233424 2984 233476 2990
rect 233424 2926 233476 2932
rect 231032 2916 231084 2922
rect 231032 2858 231084 2864
rect 232412 2916 232464 2922
rect 232412 2858 232464 2864
rect 230112 2848 230164 2854
rect 230112 2790 230164 2796
rect 231044 480 231072 2858
rect 232228 2848 232280 2854
rect 232228 2790 232280 2796
rect 232240 480 232268 2790
rect 233436 480 233464 2926
rect 233620 2854 233648 4420
rect 234816 2990 234844 4420
rect 234804 2984 234856 2990
rect 234804 2926 234856 2932
rect 235920 2922 235948 4420
rect 234620 2916 234672 2922
rect 234620 2858 234672 2864
rect 235908 2916 235960 2922
rect 235908 2858 235960 2864
rect 237012 2916 237064 2922
rect 237012 2858 237064 2864
rect 233608 2848 233660 2854
rect 233608 2790 233660 2796
rect 234632 480 234660 2858
rect 235816 2848 235868 2854
rect 235816 2790 235868 2796
rect 235828 480 235856 2790
rect 237024 480 237052 2858
rect 237116 2854 237144 4420
rect 238116 2984 238168 2990
rect 238116 2926 238168 2932
rect 237104 2848 237156 2854
rect 237104 2790 237156 2796
rect 238128 480 238156 2926
rect 238312 2922 238340 4420
rect 239416 2990 239444 4420
rect 239404 2984 239456 2990
rect 239404 2926 239456 2932
rect 238300 2916 238352 2922
rect 238300 2858 238352 2864
rect 240508 2916 240560 2922
rect 240508 2858 240560 2864
rect 239312 2848 239364 2854
rect 239312 2790 239364 2796
rect 239324 480 239352 2790
rect 240520 480 240548 2858
rect 240612 2854 240640 4420
rect 241704 2984 241756 2990
rect 241704 2926 241756 2932
rect 240600 2848 240652 2854
rect 240600 2790 240652 2796
rect 241716 480 241744 2926
rect 241808 2922 241836 4420
rect 243004 2990 243032 4420
rect 242992 2984 243044 2990
rect 242992 2926 243044 2932
rect 241796 2916 241848 2922
rect 241796 2858 241848 2864
rect 244108 2854 244136 4420
rect 245200 2916 245252 2922
rect 245200 2858 245252 2864
rect 242900 2848 242952 2854
rect 242900 2790 242952 2796
rect 244096 2848 244148 2854
rect 244096 2790 244148 2796
rect 244188 2848 244240 2854
rect 244188 2790 244240 2796
rect 242912 480 242940 2790
rect 244200 2258 244228 2790
rect 244108 2230 244228 2258
rect 244108 480 244136 2230
rect 245212 480 245240 2858
rect 245304 2854 245332 4420
rect 246396 2984 246448 2990
rect 246396 2926 246448 2932
rect 245292 2848 245344 2854
rect 245292 2790 245344 2796
rect 246408 480 246436 2926
rect 246500 2922 246528 4420
rect 247604 2990 247632 4420
rect 247592 2984 247644 2990
rect 247592 2926 247644 2932
rect 246488 2916 246540 2922
rect 246488 2858 246540 2864
rect 248800 2854 248828 4420
rect 249996 2990 250024 4420
rect 248880 2984 248932 2990
rect 248880 2926 248932 2932
rect 249984 2984 250036 2990
rect 249984 2926 250036 2932
rect 247592 2848 247644 2854
rect 247592 2790 247644 2796
rect 248788 2848 248840 2854
rect 248788 2790 248840 2796
rect 247604 480 247632 2790
rect 248892 2258 248920 2926
rect 251100 2854 251128 4420
rect 249984 2848 250036 2854
rect 249984 2790 250036 2796
rect 251088 2848 251140 2854
rect 251088 2790 251140 2796
rect 248800 2230 248920 2258
rect 248800 480 248828 2230
rect 249996 480 250024 2790
rect 252296 2242 252324 4420
rect 253492 2990 253520 4420
rect 252376 2984 252428 2990
rect 252376 2926 252428 2932
rect 253480 2984 253532 2990
rect 253480 2926 253532 2932
rect 251180 2236 251232 2242
rect 251180 2178 251232 2184
rect 252284 2236 252336 2242
rect 252284 2178 252336 2184
rect 251192 480 251220 2178
rect 252388 480 252416 2926
rect 254596 2854 254624 4420
rect 255792 2854 255820 4420
rect 256988 2854 257016 4420
rect 258092 2854 258120 4420
rect 253480 2848 253532 2854
rect 253480 2790 253532 2796
rect 254584 2848 254636 2854
rect 254584 2790 254636 2796
rect 254676 2848 254728 2854
rect 254676 2790 254728 2796
rect 255780 2848 255832 2854
rect 255780 2790 255832 2796
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 256976 2848 257028 2854
rect 256976 2790 257028 2796
rect 257068 2848 257120 2854
rect 257068 2790 257120 2796
rect 258080 2848 258132 2854
rect 258080 2790 258132 2796
rect 253492 480 253520 2790
rect 254688 480 254716 2790
rect 255884 480 255912 2790
rect 257080 480 257108 2790
rect 259288 2242 259316 4420
rect 260484 2854 260512 4420
rect 261588 2854 261616 4420
rect 262784 2854 262812 4420
rect 263980 2854 264008 4420
rect 265084 2854 265112 4420
rect 259460 2848 259512 2854
rect 259460 2790 259512 2796
rect 260472 2848 260524 2854
rect 260472 2790 260524 2796
rect 260656 2848 260708 2854
rect 260656 2790 260708 2796
rect 261576 2848 261628 2854
rect 261576 2790 261628 2796
rect 261760 2848 261812 2854
rect 261760 2790 261812 2796
rect 262772 2848 262824 2854
rect 262772 2790 262824 2796
rect 262956 2848 263008 2854
rect 262956 2790 263008 2796
rect 263968 2848 264020 2854
rect 263968 2790 264020 2796
rect 264152 2848 264204 2854
rect 264152 2790 264204 2796
rect 265072 2848 265124 2854
rect 265072 2790 265124 2796
rect 258264 2236 258316 2242
rect 258264 2178 258316 2184
rect 259276 2236 259328 2242
rect 259276 2178 259328 2184
rect 258276 480 258304 2178
rect 259472 480 259500 2790
rect 260668 480 260696 2790
rect 261772 480 261800 2790
rect 262968 480 262996 2790
rect 264164 480 264192 2790
rect 266280 2038 266308 4420
rect 267476 2854 267504 4420
rect 268672 2854 268700 4420
rect 269776 2854 269804 4420
rect 270972 2854 271000 4420
rect 272168 2854 272196 4420
rect 273272 2854 273300 4420
rect 274468 2854 274496 4420
rect 275664 2854 275692 4420
rect 266544 2848 266596 2854
rect 266544 2790 266596 2796
rect 267464 2848 267516 2854
rect 267464 2790 267516 2796
rect 267740 2848 267792 2854
rect 267740 2790 267792 2796
rect 268660 2848 268712 2854
rect 268660 2790 268712 2796
rect 268844 2848 268896 2854
rect 268844 2790 268896 2796
rect 269764 2848 269816 2854
rect 269764 2790 269816 2796
rect 270040 2848 270092 2854
rect 270040 2790 270092 2796
rect 270960 2848 271012 2854
rect 270960 2790 271012 2796
rect 271236 2848 271288 2854
rect 271236 2790 271288 2796
rect 272156 2848 272208 2854
rect 272156 2790 272208 2796
rect 272432 2848 272484 2854
rect 272432 2790 272484 2796
rect 273260 2848 273312 2854
rect 273260 2790 273312 2796
rect 273628 2848 273680 2854
rect 273628 2790 273680 2796
rect 274456 2848 274508 2854
rect 274456 2790 274508 2796
rect 274824 2848 274876 2854
rect 274824 2790 274876 2796
rect 275652 2848 275704 2854
rect 275652 2790 275704 2796
rect 265348 2032 265400 2038
rect 265348 1974 265400 1980
rect 266268 2032 266320 2038
rect 266268 1974 266320 1980
rect 265360 480 265388 1974
rect 266556 480 266584 2790
rect 267752 480 267780 2790
rect 268856 480 268884 2790
rect 270052 480 270080 2790
rect 271248 480 271276 2790
rect 272444 480 272472 2790
rect 273640 480 273668 2790
rect 274836 480 274864 2790
rect 276768 1970 276796 4420
rect 277964 2854 277992 4420
rect 279160 2854 279188 4420
rect 280264 2854 280292 4420
rect 281460 2854 281488 4420
rect 282656 2854 282684 4420
rect 277124 2848 277176 2854
rect 277124 2790 277176 2796
rect 277952 2848 278004 2854
rect 277952 2790 278004 2796
rect 278320 2848 278372 2854
rect 278320 2790 278372 2796
rect 279148 2848 279200 2854
rect 279148 2790 279200 2796
rect 279516 2848 279568 2854
rect 279516 2790 279568 2796
rect 280252 2848 280304 2854
rect 280252 2790 280304 2796
rect 280712 2848 280764 2854
rect 280712 2790 280764 2796
rect 281448 2848 281500 2854
rect 281448 2790 281500 2796
rect 281908 2848 281960 2854
rect 281908 2790 281960 2796
rect 282644 2848 282696 2854
rect 282644 2790 282696 2796
rect 276020 1964 276072 1970
rect 276020 1906 276072 1912
rect 276756 1964 276808 1970
rect 276756 1906 276808 1912
rect 276032 480 276060 1906
rect 277136 480 277164 2790
rect 278332 480 278360 2790
rect 279528 480 279556 2790
rect 280724 480 280752 2790
rect 281920 480 281948 2790
rect 283760 1698 283788 4420
rect 284956 2854 284984 4420
rect 286152 2854 286180 4420
rect 287256 2854 287284 4420
rect 288452 2854 288480 4420
rect 289648 2854 289676 4420
rect 284300 2848 284352 2854
rect 284300 2790 284352 2796
rect 284944 2848 284996 2854
rect 284944 2790 284996 2796
rect 285404 2848 285456 2854
rect 285404 2790 285456 2796
rect 286140 2848 286192 2854
rect 286140 2790 286192 2796
rect 286600 2848 286652 2854
rect 286600 2790 286652 2796
rect 287244 2848 287296 2854
rect 287244 2790 287296 2796
rect 287796 2848 287848 2854
rect 287796 2790 287848 2796
rect 288440 2848 288492 2854
rect 288440 2790 288492 2796
rect 288992 2848 289044 2854
rect 288992 2790 289044 2796
rect 289636 2848 289688 2854
rect 289636 2790 289688 2796
rect 283104 1692 283156 1698
rect 283104 1634 283156 1640
rect 283748 1692 283800 1698
rect 283748 1634 283800 1640
rect 283116 480 283144 1634
rect 284312 480 284340 2790
rect 285416 480 285444 2790
rect 286612 480 286640 2790
rect 287808 480 287836 2790
rect 289004 480 289032 2790
rect 290752 2242 290780 4420
rect 291948 2854 291976 4420
rect 293144 2854 293172 4420
rect 294340 2854 294368 4420
rect 295444 2854 295472 4420
rect 296640 2854 296668 4420
rect 291384 2848 291436 2854
rect 291384 2790 291436 2796
rect 291936 2848 291988 2854
rect 291936 2790 291988 2796
rect 292580 2848 292632 2854
rect 292580 2790 292632 2796
rect 293132 2848 293184 2854
rect 293132 2790 293184 2796
rect 293684 2848 293736 2854
rect 293684 2790 293736 2796
rect 294328 2848 294380 2854
rect 294328 2790 294380 2796
rect 294880 2848 294932 2854
rect 294880 2790 294932 2796
rect 295432 2848 295484 2854
rect 295432 2790 295484 2796
rect 296076 2848 296128 2854
rect 296076 2790 296128 2796
rect 296628 2848 296680 2854
rect 296628 2790 296680 2796
rect 290188 2236 290240 2242
rect 290188 2178 290240 2184
rect 290740 2236 290792 2242
rect 290740 2178 290792 2184
rect 290200 480 290228 2178
rect 291396 480 291424 2790
rect 292592 480 292620 2790
rect 293696 480 293724 2790
rect 294892 480 294920 2790
rect 296088 480 296116 2790
rect 297836 2242 297864 4420
rect 298940 2854 298968 4420
rect 300136 2854 300164 4420
rect 301332 2854 301360 4420
rect 302436 2854 302464 4420
rect 303632 2854 303660 4420
rect 298468 2848 298520 2854
rect 298468 2790 298520 2796
rect 298928 2848 298980 2854
rect 298928 2790 298980 2796
rect 299664 2848 299716 2854
rect 299664 2790 299716 2796
rect 300124 2848 300176 2854
rect 300124 2790 300176 2796
rect 300768 2848 300820 2854
rect 300768 2790 300820 2796
rect 301320 2848 301372 2854
rect 301320 2790 301372 2796
rect 301964 2848 302016 2854
rect 301964 2790 302016 2796
rect 302424 2848 302476 2854
rect 302424 2790 302476 2796
rect 303160 2848 303212 2854
rect 303160 2790 303212 2796
rect 303620 2848 303672 2854
rect 303620 2790 303672 2796
rect 297272 2236 297324 2242
rect 297272 2178 297324 2184
rect 297824 2236 297876 2242
rect 297824 2178 297876 2184
rect 297284 480 297312 2178
rect 298480 480 298508 2790
rect 299676 480 299704 2790
rect 300780 480 300808 2790
rect 301976 480 302004 2790
rect 303172 480 303200 2790
rect 304828 2310 304856 4420
rect 304356 2304 304408 2310
rect 304356 2246 304408 2252
rect 304816 2304 304868 2310
rect 304816 2246 304868 2252
rect 304368 480 304396 2246
rect 305564 598 305776 626
rect 305564 480 305592 598
rect 305748 490 305776 598
rect 305932 490 305960 4420
rect 307128 2258 307156 4420
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 305748 462 305960 490
rect 306760 2230 307156 2258
rect 306760 480 306788 2230
rect 307956 598 308168 626
rect 307956 480 307984 598
rect 308140 490 308168 598
rect 308324 490 308352 4420
rect 309428 2258 309456 4420
rect 310624 2258 310652 4420
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 308140 462 308352 490
rect 309060 2230 309456 2258
rect 310256 2230 310652 2258
rect 309060 480 309088 2230
rect 310256 480 310284 2230
rect 311452 598 311664 626
rect 311452 480 311480 598
rect 311636 490 311664 598
rect 311820 490 311848 4420
rect 312924 2258 312952 4420
rect 314120 2258 314148 4420
rect 315316 2258 315344 4420
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 311636 462 311848 490
rect 312648 2230 312952 2258
rect 313844 2230 314148 2258
rect 315040 2230 315344 2258
rect 312648 480 312676 2230
rect 313844 480 313872 2230
rect 315040 480 315068 2230
rect 316420 626 316448 4420
rect 317616 2258 317644 4420
rect 318812 2258 318840 4420
rect 320008 2258 320036 4420
rect 321112 2258 321140 4420
rect 316236 598 316448 626
rect 317340 2230 317644 2258
rect 318536 2230 318840 2258
rect 319732 2230 320036 2258
rect 320928 2230 321140 2258
rect 316236 480 316264 598
rect 317340 480 317368 2230
rect 318536 480 318564 2230
rect 319732 480 319760 2230
rect 320928 480 320956 2230
rect 322308 626 322336 4420
rect 323504 2258 323532 4420
rect 324608 2258 324636 4420
rect 325804 2258 325832 4420
rect 327000 2258 327028 4420
rect 328104 2258 328132 4420
rect 329300 2258 329328 4420
rect 330496 2258 330524 4420
rect 322124 598 322336 626
rect 323320 2230 323532 2258
rect 324424 2230 324636 2258
rect 325620 2230 325832 2258
rect 326816 2230 327028 2258
rect 328012 2230 328132 2258
rect 329208 2230 329328 2258
rect 330404 2230 330524 2258
rect 322124 480 322152 598
rect 323320 480 323348 2230
rect 324424 480 324452 2230
rect 325620 480 325648 2230
rect 326816 480 326844 2230
rect 328012 480 328040 2230
rect 329208 480 329236 2230
rect 330404 480 330432 2230
rect 331600 480 331628 4420
rect 332796 2258 332824 4420
rect 333992 2258 334020 4420
rect 332704 2230 332824 2258
rect 333900 2230 334020 2258
rect 332704 480 332732 2230
rect 333900 480 333928 2230
rect 335096 480 335124 4420
rect 336292 480 336320 4420
rect 337488 480 337516 4420
rect 338592 2258 338620 4420
rect 339788 2258 339816 4420
rect 338592 2230 338712 2258
rect 339788 2230 339908 2258
rect 338684 480 338712 2230
rect 339880 480 339908 2230
rect 340984 480 341012 4420
rect 342088 2258 342116 4420
rect 343284 2258 343312 4420
rect 344480 2258 344508 4420
rect 345676 2258 345704 4420
rect 346780 2258 346808 4420
rect 347976 2258 348004 4420
rect 342088 2230 342208 2258
rect 343284 2230 343404 2258
rect 344480 2230 344600 2258
rect 345676 2230 345796 2258
rect 346780 2230 346992 2258
rect 347976 2230 348096 2258
rect 342180 480 342208 2230
rect 343376 480 343404 2230
rect 344572 480 344600 2230
rect 345768 480 345796 2230
rect 346964 480 346992 2230
rect 348068 480 348096 2230
rect 349172 1850 349200 4420
rect 350276 2258 350304 4420
rect 350276 2230 350488 2258
rect 349172 1822 349292 1850
rect 349264 480 349292 1822
rect 350460 480 350488 2230
rect 351472 1714 351500 4420
rect 352668 2258 352696 4420
rect 353772 2258 353800 4420
rect 354968 2258 354996 4420
rect 356164 2258 356192 4420
rect 357268 2258 357296 4420
rect 358464 2258 358492 4420
rect 359660 2258 359688 4420
rect 360764 2258 360792 4420
rect 352668 2230 352880 2258
rect 353772 2230 354076 2258
rect 354968 2230 355272 2258
rect 356164 2230 356376 2258
rect 357268 2230 357572 2258
rect 358464 2230 358768 2258
rect 359660 2230 359964 2258
rect 360764 2230 361160 2258
rect 351472 1686 351684 1714
rect 351656 480 351684 1686
rect 352852 480 352880 2230
rect 354048 480 354076 2230
rect 355244 480 355272 2230
rect 356348 480 356376 2230
rect 357544 480 357572 2230
rect 358740 480 358768 2230
rect 359936 480 359964 2230
rect 361132 480 361160 2230
rect 361960 490 361988 4420
rect 363156 2258 363184 4420
rect 363156 2230 363552 2258
rect 362144 598 362356 626
rect 362144 490 362172 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361960 462 362172 490
rect 362328 480 362356 598
rect 363524 480 363552 2230
rect 364260 1442 364288 4420
rect 365456 2258 365484 4420
rect 366652 2258 366680 4420
rect 365456 2230 365852 2258
rect 366652 2230 367048 2258
rect 367756 2242 367784 4420
rect 368952 2854 368980 4420
rect 370148 2854 370176 4420
rect 368940 2848 368992 2854
rect 368940 2790 368992 2796
rect 369400 2848 369452 2854
rect 369400 2790 369452 2796
rect 370136 2848 370188 2854
rect 370136 2790 370188 2796
rect 370596 2848 370648 2854
rect 370596 2790 370648 2796
rect 364260 1414 364656 1442
rect 364628 480 364656 1414
rect 365824 480 365852 2230
rect 367020 480 367048 2230
rect 367744 2236 367796 2242
rect 367744 2178 367796 2184
rect 368204 2236 368256 2242
rect 368204 2178 368256 2184
rect 368216 480 368244 2178
rect 369412 480 369440 2790
rect 370608 480 370636 2790
rect 371344 490 371372 4420
rect 372448 2174 372476 4420
rect 373644 2242 373672 4420
rect 374840 2242 374868 4420
rect 375944 2854 375972 4420
rect 377140 2854 377168 4420
rect 375932 2848 375984 2854
rect 375932 2790 375984 2796
rect 376484 2848 376536 2854
rect 376484 2790 376536 2796
rect 377128 2848 377180 2854
rect 377128 2790 377180 2796
rect 377680 2848 377732 2854
rect 377680 2790 377732 2796
rect 373632 2236 373684 2242
rect 373632 2178 373684 2184
rect 374092 2236 374144 2242
rect 374092 2178 374144 2184
rect 374828 2236 374880 2242
rect 374828 2178 374880 2184
rect 375288 2236 375340 2242
rect 375288 2178 375340 2184
rect 372436 2168 372488 2174
rect 372436 2110 372488 2116
rect 372896 2168 372948 2174
rect 372896 2110 372948 2116
rect 371528 598 371740 626
rect 371528 490 371556 598
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371344 462 371556 490
rect 371712 480 371740 598
rect 372908 480 372936 2110
rect 374104 480 374132 2178
rect 375300 480 375328 2178
rect 376496 480 376524 2790
rect 377692 480 377720 2790
rect 378336 2242 378364 4420
rect 379440 2242 379468 4420
rect 380636 2310 380664 4420
rect 380624 2304 380676 2310
rect 380624 2246 380676 2252
rect 381176 2304 381228 2310
rect 381176 2246 381228 2252
rect 378324 2236 378376 2242
rect 378324 2178 378376 2184
rect 378876 2236 378928 2242
rect 378876 2178 378928 2184
rect 379428 2236 379480 2242
rect 379428 2178 379480 2184
rect 379980 2236 380032 2242
rect 379980 2178 380032 2184
rect 378888 480 378916 2178
rect 379992 480 380020 2178
rect 381188 480 381216 2246
rect 381832 2038 381860 4420
rect 382936 2854 382964 4420
rect 384132 2854 384160 4420
rect 382924 2848 382976 2854
rect 382924 2790 382976 2796
rect 383568 2848 383620 2854
rect 383568 2790 383620 2796
rect 384120 2848 384172 2854
rect 384120 2790 384172 2796
rect 384764 2848 384816 2854
rect 384764 2790 384816 2796
rect 381820 2032 381872 2038
rect 381820 1974 381872 1980
rect 382372 2032 382424 2038
rect 382372 1974 382424 1980
rect 382384 480 382412 1974
rect 383580 480 383608 2790
rect 384776 480 384804 2790
rect 385328 2242 385356 4420
rect 386432 2854 386460 4420
rect 386420 2848 386472 2854
rect 386420 2790 386472 2796
rect 387156 2848 387208 2854
rect 387156 2790 387208 2796
rect 385316 2236 385368 2242
rect 385316 2178 385368 2184
rect 385960 2236 386012 2242
rect 385960 2178 386012 2184
rect 385972 480 386000 2178
rect 387168 480 387196 2790
rect 387628 2242 387656 4420
rect 388824 2242 388852 4420
rect 389928 2242 389956 4420
rect 391124 2854 391152 4420
rect 391112 2848 391164 2854
rect 391112 2790 391164 2796
rect 391848 2848 391900 2854
rect 391848 2790 391900 2796
rect 387616 2236 387668 2242
rect 387616 2178 387668 2184
rect 388260 2236 388312 2242
rect 388260 2178 388312 2184
rect 388812 2236 388864 2242
rect 388812 2178 388864 2184
rect 389456 2236 389508 2242
rect 389456 2178 389508 2184
rect 389916 2236 389968 2242
rect 389916 2178 389968 2184
rect 390652 2236 390704 2242
rect 390652 2178 390704 2184
rect 388272 480 388300 2178
rect 389468 480 389496 2178
rect 390664 480 390692 2178
rect 391860 480 391888 2790
rect 392320 2242 392348 4420
rect 393424 2854 393452 4420
rect 393412 2848 393464 2854
rect 393412 2790 393464 2796
rect 394240 2848 394292 2854
rect 394240 2790 394292 2796
rect 392308 2236 392360 2242
rect 392308 2178 392360 2184
rect 393044 2236 393096 2242
rect 393044 2178 393096 2184
rect 393056 480 393084 2178
rect 394252 480 394280 2790
rect 394620 2242 394648 4420
rect 395816 2242 395844 4420
rect 394608 2236 394660 2242
rect 394608 2178 394660 2184
rect 395344 2236 395396 2242
rect 395344 2178 395396 2184
rect 395804 2236 395856 2242
rect 395804 2178 395856 2184
rect 396540 2236 396592 2242
rect 396540 2178 396592 2184
rect 395356 480 395384 2178
rect 396552 480 396580 2178
rect 396920 1834 396948 4420
rect 398116 2310 398144 4420
rect 398104 2304 398156 2310
rect 398104 2246 398156 2252
rect 398932 2304 398984 2310
rect 398932 2246 398984 2252
rect 396908 1828 396960 1834
rect 396908 1770 396960 1776
rect 397736 1828 397788 1834
rect 397736 1770 397788 1776
rect 397748 480 397776 1770
rect 398944 480 398972 2246
rect 399312 2242 399340 4420
rect 400508 2854 400536 4420
rect 401612 2854 401640 4420
rect 400496 2848 400548 2854
rect 400496 2790 400548 2796
rect 401324 2848 401376 2854
rect 401324 2790 401376 2796
rect 401600 2848 401652 2854
rect 401600 2790 401652 2796
rect 402520 2848 402572 2854
rect 402520 2790 402572 2796
rect 399300 2236 399352 2242
rect 399300 2178 399352 2184
rect 400128 2236 400180 2242
rect 400128 2178 400180 2184
rect 400140 480 400168 2178
rect 401336 480 401364 2790
rect 402532 480 402560 2790
rect 402808 2310 402836 4420
rect 402796 2304 402848 2310
rect 402796 2246 402848 2252
rect 403624 2304 403676 2310
rect 403624 2246 403676 2252
rect 403636 480 403664 2246
rect 404004 1426 404032 4420
rect 405108 1562 405136 4420
rect 406304 2106 406332 4420
rect 407500 2854 407528 4420
rect 408604 2854 408632 4420
rect 407488 2848 407540 2854
rect 407488 2790 407540 2796
rect 408408 2848 408460 2854
rect 408408 2790 408460 2796
rect 408592 2848 408644 2854
rect 408592 2790 408644 2796
rect 409604 2848 409656 2854
rect 409604 2790 409656 2796
rect 406292 2100 406344 2106
rect 406292 2042 406344 2048
rect 407212 2100 407264 2106
rect 407212 2042 407264 2048
rect 405096 1556 405148 1562
rect 405096 1498 405148 1504
rect 406016 1556 406068 1562
rect 406016 1498 406068 1504
rect 403992 1420 404044 1426
rect 403992 1362 404044 1368
rect 404820 1420 404872 1426
rect 404820 1362 404872 1368
rect 404832 480 404860 1362
rect 406028 480 406056 1498
rect 407224 480 407252 2042
rect 408420 480 408448 2790
rect 409616 480 409644 2790
rect 409800 2310 409828 4420
rect 409788 2304 409840 2310
rect 409788 2246 409840 2252
rect 410800 2304 410852 2310
rect 410800 2246 410852 2252
rect 410812 480 410840 2246
rect 410996 2242 411024 4420
rect 412100 2310 412128 4420
rect 412088 2304 412140 2310
rect 412088 2246 412140 2252
rect 413100 2304 413152 2310
rect 413100 2246 413152 2252
rect 410984 2236 411036 2242
rect 410984 2178 411036 2184
rect 411904 2236 411956 2242
rect 411904 2178 411956 2184
rect 411916 480 411944 2178
rect 413112 480 413140 2246
rect 413296 1562 413324 4420
rect 414492 2310 414520 4420
rect 415596 2854 415624 4420
rect 415584 2848 415636 2854
rect 415584 2790 415636 2796
rect 416688 2848 416740 2854
rect 416688 2790 416740 2796
rect 414480 2304 414532 2310
rect 414480 2246 414532 2252
rect 415492 2304 415544 2310
rect 415492 2246 415544 2252
rect 413284 1556 413336 1562
rect 413284 1498 413336 1504
rect 414296 1556 414348 1562
rect 414296 1498 414348 1504
rect 414308 480 414336 1498
rect 415504 480 415532 2246
rect 416700 480 416728 2790
rect 416792 2174 416820 4420
rect 417988 2242 418016 4420
rect 417976 2236 418028 2242
rect 417976 2178 418028 2184
rect 418988 2236 419040 2242
rect 418988 2178 419040 2184
rect 416780 2168 416832 2174
rect 416780 2110 416832 2116
rect 417884 2168 417936 2174
rect 417884 2110 417936 2116
rect 417896 480 417924 2110
rect 419000 480 419028 2178
rect 419092 1902 419120 4420
rect 420288 2174 420316 4420
rect 420276 2168 420328 2174
rect 420276 2110 420328 2116
rect 421380 2168 421432 2174
rect 421380 2110 421432 2116
rect 419080 1896 419132 1902
rect 419080 1838 419132 1844
rect 420184 1896 420236 1902
rect 420184 1838 420236 1844
rect 420196 480 420224 1838
rect 421392 480 421420 2110
rect 421484 1698 421512 4420
rect 422588 2310 422616 4420
rect 423784 2446 423812 4420
rect 424980 2582 425008 4420
rect 424968 2576 425020 2582
rect 424968 2518 425020 2524
rect 426072 2576 426124 2582
rect 426072 2518 426124 2524
rect 423772 2440 423824 2446
rect 423772 2382 423824 2388
rect 424968 2440 425020 2446
rect 424968 2382 425020 2388
rect 422576 2304 422628 2310
rect 422576 2246 422628 2252
rect 423772 2304 423824 2310
rect 423772 2246 423824 2252
rect 421472 1692 421524 1698
rect 421472 1634 421524 1640
rect 422576 1692 422628 1698
rect 422576 1634 422628 1640
rect 422588 480 422616 1634
rect 423784 480 423812 2246
rect 424980 480 425008 2382
rect 426084 2122 426112 2518
rect 426176 2242 426204 4420
rect 427280 2378 427308 4420
rect 428476 2514 428504 4420
rect 428464 2508 428516 2514
rect 428464 2450 428516 2456
rect 429568 2508 429620 2514
rect 429568 2450 429620 2456
rect 427268 2372 427320 2378
rect 427268 2314 427320 2320
rect 428464 2372 428516 2378
rect 428464 2314 428516 2320
rect 426164 2236 426216 2242
rect 426164 2178 426216 2184
rect 427268 2236 427320 2242
rect 427268 2178 427320 2184
rect 426084 2094 426204 2122
rect 426176 480 426204 2094
rect 427280 480 427308 2178
rect 428476 480 428504 2314
rect 429580 1850 429608 2450
rect 429672 2310 429700 4420
rect 429660 2304 429712 2310
rect 429660 2246 429712 2252
rect 430776 2174 430804 4420
rect 431972 2854 432000 4420
rect 431960 2848 432012 2854
rect 431960 2790 432012 2796
rect 430856 2304 430908 2310
rect 430856 2246 430908 2252
rect 430764 2168 430816 2174
rect 430764 2110 430816 2116
rect 429580 1822 429700 1850
rect 429672 480 429700 1822
rect 430868 480 430896 2246
rect 432052 2168 432104 2174
rect 432052 2110 432104 2116
rect 432064 480 432092 2110
rect 433168 1562 433196 4420
rect 433248 2848 433300 2854
rect 433248 2790 433300 2796
rect 433156 1556 433208 1562
rect 433156 1498 433208 1504
rect 433260 480 433288 2790
rect 434272 2174 434300 4420
rect 435468 2310 435496 4420
rect 435456 2304 435508 2310
rect 435456 2246 435508 2252
rect 436664 2174 436692 4420
rect 436744 2304 436796 2310
rect 436744 2246 436796 2252
rect 434260 2168 434312 2174
rect 434260 2110 434312 2116
rect 435548 2168 435600 2174
rect 435548 2110 435600 2116
rect 436652 2168 436704 2174
rect 436652 2110 436704 2116
rect 434444 1556 434496 1562
rect 434444 1498 434496 1504
rect 434456 480 434484 1498
rect 435560 480 435588 2110
rect 436756 480 436784 2246
rect 437768 2242 437796 4420
rect 438964 2310 438992 4420
rect 438952 2304 439004 2310
rect 438952 2246 439004 2252
rect 437756 2236 437808 2242
rect 437756 2178 437808 2184
rect 439136 2236 439188 2242
rect 439136 2178 439188 2184
rect 437940 2168 437992 2174
rect 437940 2110 437992 2116
rect 437952 480 437980 2110
rect 439148 480 439176 2178
rect 440160 2038 440188 4420
rect 441264 2310 441292 4420
rect 440332 2304 440384 2310
rect 440332 2246 440384 2252
rect 441252 2304 441304 2310
rect 441252 2246 441304 2252
rect 440148 2032 440200 2038
rect 440148 1974 440200 1980
rect 440344 480 440372 2246
rect 441528 2032 441580 2038
rect 441528 1974 441580 1980
rect 441540 480 441568 1974
rect 442460 1970 442488 4420
rect 442632 2304 442684 2310
rect 442632 2246 442684 2252
rect 442448 1964 442500 1970
rect 442448 1906 442500 1912
rect 442644 480 442672 2246
rect 443656 2242 443684 4420
rect 443644 2236 443696 2242
rect 443644 2178 443696 2184
rect 444760 2174 444788 4420
rect 445024 2236 445076 2242
rect 445024 2178 445076 2184
rect 444748 2168 444800 2174
rect 444748 2110 444800 2116
rect 443828 1964 443880 1970
rect 443828 1906 443880 1912
rect 443840 480 443868 1906
rect 445036 480 445064 2178
rect 445956 1698 445984 4420
rect 447152 2174 447180 4420
rect 446220 2168 446272 2174
rect 446220 2110 446272 2116
rect 447140 2168 447192 2174
rect 447140 2110 447192 2116
rect 445944 1692 445996 1698
rect 445944 1634 445996 1640
rect 446232 480 446260 2110
rect 448256 1698 448284 4420
rect 448612 2168 448664 2174
rect 448612 2110 448664 2116
rect 447416 1692 447468 1698
rect 447416 1634 447468 1640
rect 448244 1692 448296 1698
rect 448244 1634 448296 1640
rect 447428 480 447456 1634
rect 448624 480 448652 2110
rect 449452 2106 449480 4420
rect 450648 2310 450676 4420
rect 450636 2304 450688 2310
rect 450636 2246 450688 2252
rect 451844 2242 451872 4420
rect 452948 2310 452976 4420
rect 452108 2304 452160 2310
rect 452108 2246 452160 2252
rect 452936 2304 452988 2310
rect 452936 2246 452988 2252
rect 451832 2236 451884 2242
rect 451832 2178 451884 2184
rect 449440 2100 449492 2106
rect 449440 2042 449492 2048
rect 450912 2100 450964 2106
rect 450912 2042 450964 2048
rect 449808 1692 449860 1698
rect 449808 1634 449860 1640
rect 449820 480 449848 1634
rect 450924 480 450952 2042
rect 452120 480 452148 2246
rect 453304 2236 453356 2242
rect 453304 2178 453356 2184
rect 453316 480 453344 2178
rect 454144 2174 454172 4420
rect 454500 2304 454552 2310
rect 454500 2246 454552 2252
rect 454132 2168 454184 2174
rect 454132 2110 454184 2116
rect 454512 480 454540 2246
rect 455340 2106 455368 4420
rect 455696 2168 455748 2174
rect 455696 2110 455748 2116
rect 455328 2100 455380 2106
rect 455328 2042 455380 2048
rect 455708 480 455736 2110
rect 456444 1562 456472 4420
rect 456892 2100 456944 2106
rect 456892 2042 456944 2048
rect 456432 1556 456484 1562
rect 456432 1498 456484 1504
rect 456904 480 456932 2042
rect 457640 1494 457668 4420
rect 458836 2242 458864 4420
rect 458824 2236 458876 2242
rect 458824 2178 458876 2184
rect 459940 1902 459968 4420
rect 460388 2236 460440 2242
rect 460388 2178 460440 2184
rect 459928 1896 459980 1902
rect 459928 1838 459980 1844
rect 458088 1556 458140 1562
rect 458088 1498 458140 1504
rect 457628 1488 457680 1494
rect 457628 1430 457680 1436
rect 458100 480 458128 1498
rect 459192 1488 459244 1494
rect 459192 1430 459244 1436
rect 459204 480 459232 1430
rect 460400 480 460428 2178
rect 461136 1494 461164 4420
rect 461584 1896 461636 1902
rect 461584 1838 461636 1844
rect 461124 1488 461176 1494
rect 461124 1430 461176 1436
rect 461596 480 461624 1838
rect 462332 1766 462360 4420
rect 463436 2242 463464 4420
rect 463424 2236 463476 2242
rect 463424 2178 463476 2184
rect 462320 1760 462372 1766
rect 462320 1702 462372 1708
rect 463976 1760 464028 1766
rect 463976 1702 464028 1708
rect 462780 1488 462832 1494
rect 462780 1430 462832 1436
rect 462792 480 462820 1430
rect 463988 480 464016 1702
rect 464632 1494 464660 4420
rect 465172 2236 465224 2242
rect 465172 2178 465224 2184
rect 464620 1488 464672 1494
rect 464620 1430 464672 1436
rect 465184 480 465212 2178
rect 465828 1562 465856 4420
rect 466932 2242 466960 4420
rect 466920 2236 466972 2242
rect 466920 2178 466972 2184
rect 468128 1630 468156 4420
rect 468668 2236 468720 2242
rect 468668 2178 468720 2184
rect 468116 1624 468168 1630
rect 468116 1566 468168 1572
rect 465816 1556 465868 1562
rect 465816 1498 465868 1504
rect 467472 1556 467524 1562
rect 467472 1498 467524 1504
rect 466276 1488 466328 1494
rect 466276 1430 466328 1436
rect 466288 480 466316 1430
rect 467484 480 467512 1498
rect 468680 480 468708 2178
rect 469324 1562 469352 4420
rect 470428 2786 470456 4420
rect 470416 2780 470468 2786
rect 470416 2722 470468 2728
rect 471624 2242 471652 4420
rect 472256 2848 472308 2854
rect 472256 2790 472308 2796
rect 471612 2236 471664 2242
rect 471612 2178 471664 2184
rect 469864 1624 469916 1630
rect 469864 1566 469916 1572
rect 469312 1556 469364 1562
rect 469312 1498 469364 1504
rect 469876 480 469904 1566
rect 471060 1556 471112 1562
rect 471060 1498 471112 1504
rect 471072 480 471100 1498
rect 472268 480 472296 2790
rect 472820 1698 472848 4420
rect 473924 2242 473952 4420
rect 473452 2236 473504 2242
rect 473452 2178 473504 2184
rect 473912 2236 473964 2242
rect 473912 2178 473964 2184
rect 472808 1692 472860 1698
rect 472808 1634 472860 1640
rect 473464 480 473492 2178
rect 475120 1698 475148 4420
rect 476316 2242 476344 4420
rect 475752 2236 475804 2242
rect 475752 2178 475804 2184
rect 476304 2236 476356 2242
rect 476304 2178 476356 2184
rect 474556 1692 474608 1698
rect 474556 1634 474608 1640
rect 475108 1692 475160 1698
rect 475108 1634 475160 1640
rect 474568 480 474596 1634
rect 475764 480 475792 2178
rect 476948 1692 477000 1698
rect 476948 1634 477000 1640
rect 476960 480 476988 1634
rect 477512 1562 477540 4420
rect 478616 2786 478644 4420
rect 478604 2780 478656 2786
rect 478604 2722 478656 2728
rect 479812 2242 479840 4420
rect 480536 2848 480588 2854
rect 480536 2790 480588 2796
rect 478144 2236 478196 2242
rect 478144 2178 478196 2184
rect 479800 2236 479852 2242
rect 479800 2178 479852 2184
rect 477500 1556 477552 1562
rect 477500 1498 477552 1504
rect 478156 480 478184 2178
rect 479340 1556 479392 1562
rect 479340 1498 479392 1504
rect 479352 480 479380 1498
rect 480548 480 480576 2790
rect 481008 1630 481036 4420
rect 481732 2236 481784 2242
rect 481732 2178 481784 2184
rect 480996 1624 481048 1630
rect 480996 1566 481048 1572
rect 481744 480 481772 2178
rect 482112 1766 482140 4420
rect 483308 2242 483336 4420
rect 483296 2236 483348 2242
rect 483296 2178 483348 2184
rect 482100 1760 482152 1766
rect 482100 1702 482152 1708
rect 484032 1760 484084 1766
rect 484032 1702 484084 1708
rect 482836 1624 482888 1630
rect 482836 1566 482888 1572
rect 482848 480 482876 1566
rect 484044 480 484072 1702
rect 484504 1630 484532 4420
rect 485608 2786 485636 4420
rect 485596 2780 485648 2786
rect 485596 2722 485648 2728
rect 486804 2310 486832 4420
rect 487620 2848 487672 2854
rect 487620 2790 487672 2796
rect 486792 2304 486844 2310
rect 486792 2246 486844 2252
rect 485228 2236 485280 2242
rect 485228 2178 485280 2184
rect 484492 1624 484544 1630
rect 484492 1566 484544 1572
rect 485240 480 485268 2178
rect 486424 1624 486476 1630
rect 486424 1566 486476 1572
rect 486436 480 486464 1566
rect 487632 480 487660 2790
rect 488000 2242 488028 4420
rect 488816 2304 488868 2310
rect 488816 2246 488868 2252
rect 487988 2236 488040 2242
rect 487988 2178 488040 2184
rect 488828 480 488856 2246
rect 489104 1970 489132 4420
rect 489920 2236 489972 2242
rect 489920 2178 489972 2184
rect 489092 1964 489144 1970
rect 489092 1906 489144 1912
rect 489932 480 489960 2178
rect 490300 1834 490328 4420
rect 491116 1964 491168 1970
rect 491116 1906 491168 1912
rect 490288 1828 490340 1834
rect 490288 1770 490340 1776
rect 491128 480 491156 1906
rect 491496 1766 491524 4420
rect 492600 2938 492628 4420
rect 492600 2910 492720 2938
rect 492692 2854 492720 2910
rect 492680 2848 492732 2854
rect 492680 2790 492732 2796
rect 493796 2786 493824 4420
rect 494704 2848 494756 2854
rect 494704 2790 494756 2796
rect 493784 2780 493836 2786
rect 493784 2722 493836 2728
rect 492312 1828 492364 1834
rect 492312 1770 492364 1776
rect 491484 1760 491536 1766
rect 491484 1702 491536 1708
rect 492324 480 492352 1770
rect 493508 1760 493560 1766
rect 493508 1702 493560 1708
rect 493520 480 493548 1702
rect 494716 480 494744 2790
rect 494992 2310 495020 4420
rect 495900 2848 495952 2854
rect 495900 2790 495952 2796
rect 494980 2304 495032 2310
rect 494980 2246 495032 2252
rect 495912 480 495940 2790
rect 496096 2242 496124 4420
rect 497292 2310 497320 4420
rect 497096 2304 497148 2310
rect 497096 2246 497148 2252
rect 497280 2304 497332 2310
rect 497280 2246 497332 2252
rect 496084 2236 496136 2242
rect 496084 2178 496136 2184
rect 497108 480 497136 2246
rect 498200 2236 498252 2242
rect 498200 2178 498252 2184
rect 498212 480 498240 2178
rect 498488 1834 498516 4420
rect 499396 2304 499448 2310
rect 499396 2246 499448 2252
rect 498476 1828 498528 1834
rect 498476 1770 498528 1776
rect 499408 480 499436 2246
rect 499592 1766 499620 4420
rect 500788 2786 500816 4420
rect 500776 2780 500828 2786
rect 500776 2722 500828 2728
rect 501984 2242 502012 4420
rect 502984 2848 503036 2854
rect 502984 2790 503036 2796
rect 501972 2236 502024 2242
rect 501972 2178 502024 2184
rect 500592 1828 500644 1834
rect 500592 1770 500644 1776
rect 499580 1760 499632 1766
rect 499580 1702 499632 1708
rect 500604 480 500632 1770
rect 501788 1760 501840 1766
rect 501788 1702 501840 1708
rect 501800 480 501828 1702
rect 502996 480 503024 2790
rect 503180 2786 503208 4420
rect 503168 2780 503220 2786
rect 503168 2722 503220 2728
rect 504284 2242 504312 4420
rect 505376 2848 505428 2854
rect 505376 2790 505428 2796
rect 504180 2236 504232 2242
rect 504180 2178 504232 2184
rect 504272 2236 504324 2242
rect 504272 2178 504324 2184
rect 504192 480 504220 2178
rect 505388 480 505416 2790
rect 505480 1834 505508 4420
rect 506676 2242 506704 4420
rect 507780 2938 507808 4420
rect 507780 2910 507900 2938
rect 507872 2854 507900 2910
rect 507860 2848 507912 2854
rect 507860 2790 507912 2796
rect 508976 2242 509004 4420
rect 510068 2848 510120 2854
rect 510068 2790 510120 2796
rect 506480 2236 506532 2242
rect 506480 2178 506532 2184
rect 506664 2236 506716 2242
rect 506664 2178 506716 2184
rect 508872 2236 508924 2242
rect 508872 2178 508924 2184
rect 508964 2236 509016 2242
rect 508964 2178 509016 2184
rect 505468 1828 505520 1834
rect 505468 1770 505520 1776
rect 506492 480 506520 2178
rect 507676 1828 507728 1834
rect 507676 1770 507728 1776
rect 507688 480 507716 1770
rect 508884 480 508912 2178
rect 510080 480 510108 2790
rect 510172 2786 510200 4420
rect 510160 2780 510212 2786
rect 510160 2722 510212 2728
rect 511276 2378 511304 4420
rect 512472 2938 512500 4420
rect 512472 2910 512592 2938
rect 512460 2848 512512 2854
rect 512460 2790 512512 2796
rect 511264 2372 511316 2378
rect 511264 2314 511316 2320
rect 511264 2236 511316 2242
rect 511264 2178 511316 2184
rect 511276 480 511304 2178
rect 512472 480 512500 2790
rect 512564 2242 512592 2910
rect 513564 2372 513616 2378
rect 513564 2314 513616 2320
rect 512552 2236 512604 2242
rect 512552 2178 512604 2184
rect 513576 480 513604 2314
rect 513668 1970 513696 4420
rect 514772 2378 514800 4420
rect 515968 2786 515996 4420
rect 517164 2786 517192 4420
rect 515956 2780 516008 2786
rect 515956 2722 516008 2728
rect 517152 2780 517204 2786
rect 517152 2722 517204 2728
rect 514760 2372 514812 2378
rect 514760 2314 514812 2320
rect 517152 2372 517204 2378
rect 517152 2314 517204 2320
rect 514760 2236 514812 2242
rect 514760 2178 514812 2184
rect 513656 1964 513708 1970
rect 513656 1906 513708 1912
rect 514772 480 514800 2178
rect 515956 1964 516008 1970
rect 515956 1906 516008 1912
rect 515968 480 515996 1906
rect 517164 480 517192 2314
rect 518268 2242 518296 4420
rect 518348 2848 518400 2854
rect 518348 2790 518400 2796
rect 518256 2236 518308 2242
rect 518256 2178 518308 2184
rect 518360 480 518388 2790
rect 519464 2786 519492 4420
rect 519544 2848 519596 2854
rect 519544 2790 519596 2796
rect 519452 2780 519504 2786
rect 519452 2722 519504 2728
rect 519556 480 519584 2790
rect 520660 2310 520688 4420
rect 520648 2304 520700 2310
rect 520648 2246 520700 2252
rect 521764 2242 521792 4420
rect 522960 2938 522988 4420
rect 522960 2910 523080 2938
rect 523052 2854 523080 2910
rect 521844 2848 521896 2854
rect 521844 2790 521896 2796
rect 523040 2848 523092 2854
rect 523040 2790 523092 2796
rect 520740 2236 520792 2242
rect 520740 2178 520792 2184
rect 521752 2236 521804 2242
rect 521752 2178 521804 2184
rect 520752 480 520780 2178
rect 521856 480 521884 2790
rect 524156 2786 524184 4420
rect 524144 2780 524196 2786
rect 524144 2722 524196 2728
rect 525260 2718 525288 4420
rect 525432 2848 525484 2854
rect 525432 2790 525484 2796
rect 525248 2712 525300 2718
rect 525248 2654 525300 2660
rect 523040 2304 523092 2310
rect 523040 2246 523092 2252
rect 523052 480 523080 2246
rect 524236 2236 524288 2242
rect 524236 2178 524288 2184
rect 524248 480 524276 2178
rect 525444 480 525472 2790
rect 526456 2310 526484 4420
rect 526628 2848 526680 2854
rect 526628 2790 526680 2796
rect 526444 2304 526496 2310
rect 526444 2246 526496 2252
rect 526640 480 526668 2790
rect 527652 2242 527680 4420
rect 527824 2848 527876 2854
rect 527824 2790 527876 2796
rect 527640 2236 527692 2242
rect 527640 2178 527692 2184
rect 527836 480 527864 2790
rect 528848 1970 528876 4420
rect 529020 2304 529072 2310
rect 529020 2246 529072 2252
rect 528836 1964 528888 1970
rect 528836 1906 528888 1912
rect 529032 480 529060 2246
rect 529952 1834 529980 4420
rect 531148 2786 531176 4420
rect 531136 2780 531188 2786
rect 531136 2722 531188 2728
rect 532344 2718 532372 4420
rect 532332 2712 532384 2718
rect 532332 2654 532384 2660
rect 533448 2242 533476 4420
rect 533712 2848 533764 2854
rect 533712 2790 533764 2796
rect 530124 2236 530176 2242
rect 530124 2178 530176 2184
rect 533436 2236 533488 2242
rect 533436 2178 533488 2184
rect 529940 1828 529992 1834
rect 529940 1770 529992 1776
rect 530136 480 530164 2178
rect 531320 1964 531372 1970
rect 531320 1906 531372 1912
rect 531332 480 531360 1906
rect 532516 1828 532568 1834
rect 532516 1770 532568 1776
rect 532528 480 532556 1770
rect 533724 480 533752 2790
rect 534644 2786 534672 4420
rect 534908 2848 534960 2854
rect 534908 2790 534960 2796
rect 534632 2780 534684 2786
rect 534632 2722 534684 2728
rect 534920 480 534948 2790
rect 535840 2310 535868 4420
rect 536944 2310 536972 4420
rect 538140 2938 538168 4420
rect 538140 2910 538260 2938
rect 538232 2854 538260 2910
rect 537208 2848 537260 2854
rect 537208 2790 537260 2796
rect 538220 2848 538272 2854
rect 538220 2790 538272 2796
rect 535828 2304 535880 2310
rect 535828 2246 535880 2252
rect 536932 2304 536984 2310
rect 536932 2246 536984 2252
rect 536104 2236 536156 2242
rect 536104 2178 536156 2184
rect 536116 480 536144 2178
rect 537220 480 537248 2790
rect 539336 2786 539364 4420
rect 540440 2922 540468 4420
rect 540428 2916 540480 2922
rect 540428 2858 540480 2864
rect 540796 2848 540848 2854
rect 540796 2790 540848 2796
rect 539324 2780 539376 2786
rect 539324 2722 539376 2728
rect 539600 2304 539652 2310
rect 539600 2246 539652 2252
rect 538404 2236 538456 2242
rect 538404 2178 538456 2184
rect 538416 480 538444 2178
rect 539612 480 539640 2246
rect 540808 480 540836 2790
rect 541636 2786 541664 4420
rect 541992 2848 542044 2854
rect 541992 2790 542044 2796
rect 541624 2780 541676 2786
rect 541624 2722 541676 2728
rect 542004 480 542032 2790
rect 542832 2786 542860 4420
rect 543188 2916 543240 2922
rect 543188 2858 543240 2864
rect 542820 2780 542872 2786
rect 542820 2722 542872 2728
rect 543200 480 543228 2858
rect 543936 2242 543964 4420
rect 544384 2848 544436 2854
rect 544384 2790 544436 2796
rect 543924 2236 543976 2242
rect 543924 2178 543976 2184
rect 544396 480 544424 2790
rect 545132 2310 545160 4420
rect 545488 2848 545540 2854
rect 545488 2790 545540 2796
rect 545120 2304 545172 2310
rect 545120 2246 545172 2252
rect 545500 480 545528 2790
rect 546328 2786 546356 4420
rect 547432 2922 547460 4420
rect 547420 2916 547472 2922
rect 547420 2858 547472 2864
rect 548628 2786 548656 4420
rect 549076 2848 549128 2854
rect 549076 2790 549128 2796
rect 546316 2780 546368 2786
rect 546316 2722 546368 2728
rect 548616 2780 548668 2786
rect 548616 2722 548668 2728
rect 547880 2304 547932 2310
rect 547880 2246 547932 2252
rect 546684 2236 546736 2242
rect 546684 2178 546736 2184
rect 546696 480 546724 2178
rect 547892 480 547920 2246
rect 549088 480 549116 2790
rect 549824 2718 549852 4420
rect 550272 2916 550324 2922
rect 550272 2858 550324 2864
rect 549812 2712 549864 2718
rect 549812 2654 549864 2660
rect 550284 480 550312 2858
rect 550928 2242 550956 4420
rect 551468 2848 551520 2854
rect 551468 2790 551520 2796
rect 550916 2236 550968 2242
rect 550916 2178 550968 2184
rect 551480 480 551508 2790
rect 552124 2786 552152 4420
rect 553320 2904 553348 4420
rect 553400 2916 553452 2922
rect 553320 2876 553400 2904
rect 553400 2858 553452 2864
rect 552664 2848 552716 2854
rect 552664 2790 552716 2796
rect 552112 2780 552164 2786
rect 552112 2722 552164 2728
rect 552676 480 552704 2790
rect 554516 2718 554544 4420
rect 554964 2848 555016 2854
rect 554964 2790 555016 2796
rect 554504 2712 554556 2718
rect 554504 2654 554556 2660
rect 553768 2236 553820 2242
rect 553768 2178 553820 2184
rect 553780 480 553808 2178
rect 554976 480 555004 2790
rect 555620 2786 555648 4420
rect 556160 2916 556212 2922
rect 556160 2858 556212 2864
rect 555608 2780 555660 2786
rect 555608 2722 555660 2728
rect 556172 480 556200 2858
rect 556816 2242 556844 4420
rect 557356 2848 557408 2854
rect 557356 2790 557408 2796
rect 556804 2236 556856 2242
rect 556804 2178 556856 2184
rect 557368 480 557396 2790
rect 558012 2786 558040 4420
rect 558552 2848 558604 2854
rect 558552 2790 558604 2796
rect 558000 2780 558052 2786
rect 558000 2722 558052 2728
rect 558564 480 558592 2790
rect 559116 2310 559144 4420
rect 560312 2786 560340 4420
rect 561508 2938 561536 4420
rect 561508 2922 561720 2938
rect 561508 2916 561732 2922
rect 561508 2910 561680 2916
rect 561680 2858 561732 2864
rect 560852 2848 560904 2854
rect 560852 2790 560904 2796
rect 560300 2780 560352 2786
rect 560300 2722 560352 2728
rect 559104 2304 559156 2310
rect 559104 2246 559156 2252
rect 559748 2236 559800 2242
rect 559748 2178 559800 2184
rect 559760 480 559788 2178
rect 560864 480 560892 2790
rect 562612 2718 562640 4420
rect 563244 2848 563296 2854
rect 563244 2790 563296 2796
rect 562600 2712 562652 2718
rect 562600 2654 562652 2660
rect 562048 2304 562100 2310
rect 562048 2246 562100 2252
rect 562060 480 562088 2246
rect 563256 480 563284 2790
rect 563808 2650 563836 4420
rect 564440 2916 564492 2922
rect 564440 2858 564492 2864
rect 563796 2644 563848 2650
rect 563796 2586 563848 2592
rect 564452 480 564480 2858
rect 565004 2242 565032 4420
rect 565636 2848 565688 2854
rect 565636 2790 565688 2796
rect 564992 2236 565044 2242
rect 564992 2178 565044 2184
rect 565648 480 565676 2790
rect 566108 2786 566136 4420
rect 566832 2848 566884 2854
rect 566832 2790 566884 2796
rect 566096 2780 566148 2786
rect 566096 2722 566148 2728
rect 566844 480 566872 2790
rect 567304 2786 567332 4420
rect 568500 2938 568528 4420
rect 568500 2922 568620 2938
rect 568500 2916 568632 2922
rect 568500 2910 568580 2916
rect 568580 2858 568632 2864
rect 569132 2848 569184 2854
rect 569132 2790 569184 2796
rect 567292 2780 567344 2786
rect 567292 2722 567344 2728
rect 568028 2236 568080 2242
rect 568028 2178 568080 2184
rect 568040 480 568068 2178
rect 569144 480 569172 2790
rect 569604 2718 569632 4420
rect 570800 2990 570828 4420
rect 570788 2984 570840 2990
rect 570788 2926 570840 2932
rect 571524 2916 571576 2922
rect 571524 2858 571576 2864
rect 570328 2848 570380 2854
rect 570328 2790 570380 2796
rect 569592 2712 569644 2718
rect 569592 2654 569644 2660
rect 570340 480 570368 2790
rect 571536 480 571564 2858
rect 571996 2786 572024 4420
rect 572720 2848 572772 2854
rect 572720 2790 572772 2796
rect 571984 2780 572036 2786
rect 571984 2722 572036 2728
rect 572732 480 572760 2790
rect 573100 2174 573128 4420
rect 573916 2984 573968 2990
rect 573916 2926 573968 2932
rect 573088 2168 573140 2174
rect 573088 2110 573140 2116
rect 573928 480 573956 2926
rect 574296 2786 574324 4420
rect 575112 2848 575164 2854
rect 575112 2790 575164 2796
rect 574284 2780 574336 2786
rect 574284 2722 574336 2728
rect 575124 480 575152 2790
rect 575492 2242 575520 4420
rect 575480 2236 575532 2242
rect 575480 2178 575532 2184
rect 576308 2168 576360 2174
rect 576308 2110 576360 2116
rect 576320 480 576348 2110
rect 576596 2106 576624 4420
rect 577412 2848 577464 2854
rect 577412 2790 577464 2796
rect 576584 2100 576636 2106
rect 576584 2042 576636 2048
rect 577424 480 577452 2790
rect 577792 2786 577820 4420
rect 577780 2780 577832 2786
rect 577780 2722 577832 2728
rect 578988 2242 579016 4420
rect 582576 4146 582604 701150
rect 582746 698048 582802 698057
rect 582746 697983 582802 697992
rect 582654 697640 582710 697649
rect 582654 697575 582710 697584
rect 582668 298761 582696 697575
rect 582760 404977 582788 697983
rect 582838 697368 582894 697377
rect 582838 697303 582894 697312
rect 582852 484673 582880 697303
rect 582930 696960 582986 696969
rect 582930 696895 582986 696904
rect 582944 591025 582972 696895
rect 582930 591016 582986 591025
rect 582930 590951 582986 590960
rect 583392 537872 583444 537878
rect 583390 537840 583392 537849
rect 583444 537840 583446 537849
rect 583390 537775 583446 537784
rect 582838 484664 582894 484673
rect 582838 484599 582894 484608
rect 583392 431656 583444 431662
rect 583390 431624 583392 431633
rect 583444 431624 583446 431633
rect 583390 431559 583446 431568
rect 583392 418328 583444 418334
rect 583390 418296 583392 418305
rect 583444 418296 583446 418305
rect 583390 418231 583446 418240
rect 582746 404968 582802 404977
rect 582746 404903 582802 404912
rect 583392 351960 583444 351966
rect 583390 351928 583392 351937
rect 583444 351928 583446 351937
rect 583390 351863 583446 351872
rect 583392 325304 583444 325310
rect 583390 325272 583392 325281
rect 583444 325272 583446 325281
rect 583390 325207 583446 325216
rect 583392 312112 583444 312118
rect 583390 312080 583392 312089
rect 583444 312080 583446 312089
rect 583390 312015 583446 312024
rect 582654 298752 582710 298761
rect 582654 298687 582710 298696
rect 583300 272264 583352 272270
rect 583298 272232 583300 272241
rect 583352 272232 583354 272241
rect 583298 272167 583354 272176
rect 583208 245608 583260 245614
rect 583206 245576 583208 245585
rect 583260 245576 583262 245585
rect 583206 245511 583262 245520
rect 583116 232416 583168 232422
rect 583114 232384 583116 232393
rect 583168 232384 583170 232393
rect 583114 232319 583170 232328
rect 583024 205760 583076 205766
rect 583022 205728 583024 205737
rect 583076 205728 583078 205737
rect 583022 205663 583078 205672
rect 582932 192568 582984 192574
rect 582930 192536 582932 192545
rect 582984 192536 582986 192545
rect 582930 192471 582986 192480
rect 582840 179240 582892 179246
rect 582838 179208 582840 179217
rect 582892 179208 582894 179217
rect 582838 179143 582894 179152
rect 582748 165912 582800 165918
rect 582746 165880 582748 165889
rect 582800 165880 582802 165889
rect 582746 165815 582802 165824
rect 582656 152720 582708 152726
rect 582654 152688 582656 152697
rect 582708 152688 582710 152697
rect 582654 152623 582710 152632
rect 582656 126064 582708 126070
rect 582654 126032 582656 126041
rect 582708 126032 582710 126041
rect 582654 125967 582710 125976
rect 582656 112872 582708 112878
rect 582654 112840 582656 112849
rect 582708 112840 582710 112849
rect 582654 112775 582710 112784
rect 582564 4140 582616 4146
rect 582564 4082 582616 4088
rect 582196 2848 582248 2854
rect 582196 2790 582248 2796
rect 578608 2236 578660 2242
rect 578608 2178 578660 2184
rect 578976 2236 579028 2242
rect 578976 2178 579028 2184
rect 578620 480 578648 2178
rect 581000 2100 581052 2106
rect 581000 2042 581052 2048
rect 581012 480 581040 2042
rect 582208 480 582236 2790
rect 583392 2236 583444 2242
rect 583392 2178 583444 2184
rect 583404 480 583432 2178
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 294 701392 350 701448
rect 846 697040 902 697096
rect 1490 684256 1546 684312
rect 1582 658144 1638 658200
rect 1674 632032 1730 632088
rect 846 606056 902 606112
rect 1766 579944 1822 580000
rect 754 553832 810 553888
rect 2042 701664 2098 701720
rect 1950 698128 2006 698184
rect 1858 527856 1914 527912
rect 1950 475632 2006 475688
rect 662 449520 718 449576
rect 570 345344 626 345400
rect 570 267144 626 267200
rect 570 214920 626 214976
rect 570 136720 626 136776
rect 202 111152 258 111208
rect 110 71848 166 71904
rect 2318 697448 2374 697504
rect 4526 701256 4582 701312
rect 2502 697720 2558 697776
rect 2410 423544 2466 423600
rect 2686 697856 2742 697912
rect 2594 501744 2650 501800
rect 3054 619112 3110 619168
rect 3422 700304 3478 700360
rect 3238 566888 3294 566944
rect 3146 514800 3202 514856
rect 2778 462576 2834 462632
rect 2686 397432 2742 397488
rect 2502 371320 2558 371376
rect 2318 319232 2374 319288
rect 2778 306212 2780 306232
rect 2780 306212 2832 306232
rect 2832 306212 2834 306232
rect 2778 306176 2834 306212
rect 3330 410488 3386 410544
rect 3238 254088 3294 254144
rect 2226 241032 2282 241088
rect 2134 162832 2190 162888
rect 2042 58520 2098 58576
rect 18 32952 74 33008
rect 3514 698400 3570 698456
rect 3698 671200 3754 671256
rect 3606 97552 3662 97608
rect 3514 84632 3570 84688
rect 4802 358400 4858 358456
rect 27066 699760 27122 699816
rect 62394 699896 62450 699952
rect 107750 700032 107806 700088
rect 218058 701528 218114 701584
rect 223854 700168 223910 700224
rect 526534 701392 526590 701448
rect 531594 701528 531650 701584
rect 556802 701256 556858 701312
rect 554778 700304 554834 700360
rect 561862 701664 561918 701720
rect 580446 699896 580502 699952
rect 143354 699080 143410 699136
rect 163594 699080 163650 699136
rect 193770 699080 193826 699136
rect 390098 699080 390154 699136
rect 430762 699080 430818 699136
rect 450726 699080 450782 699136
rect 461030 699080 461086 699136
rect 476210 699080 476266 699136
rect 541346 699080 541402 699136
rect 17222 698944 17278 699000
rect 112994 698944 113050 699000
rect 132682 698944 132738 699000
rect 579894 697176 579950 697232
rect 579894 696904 579950 696960
rect 579986 683848 580042 683904
rect 579158 644000 579214 644056
rect 580078 630808 580134 630864
rect 580262 698944 580318 699000
rect 580170 577632 580226 577688
rect 4066 293120 4122 293176
rect 3974 201864 4030 201920
rect 3882 188808 3938 188864
rect 3790 149776 3846 149832
rect 580630 700032 580686 700088
rect 580538 365064 580594 365120
rect 581550 670656 581606 670712
rect 580906 524456 580962 524512
rect 580814 471416 580870 471472
rect 580722 378392 580778 378448
rect 580630 258848 580686 258904
rect 580446 139304 580502 139360
rect 580354 99456 580410 99512
rect 580262 59608 580318 59664
rect 3698 45464 3754 45520
rect 3422 19352 3478 19408
rect 582470 699760 582526 699816
rect 582378 698264 582434 698320
rect 582286 617480 582342 617536
rect 582194 564304 582250 564360
rect 582102 511264 582158 511320
rect 582010 458088 582066 458144
rect 581918 219000 581974 219056
rect 581826 86128 581882 86184
rect 581734 46280 581790 46336
rect 582470 72936 582526 72992
rect 582470 33108 582526 33144
rect 582470 33088 582472 33108
rect 582472 33088 582524 33108
rect 582524 33088 582526 33108
rect 582378 19760 582434 19816
rect 581642 6568 581698 6624
rect 3422 6432 3478 6488
rect 582746 697992 582802 698048
rect 582654 697584 582710 697640
rect 582838 697312 582894 697368
rect 582930 696904 582986 696960
rect 582930 590960 582986 591016
rect 583390 537820 583392 537840
rect 583392 537820 583444 537840
rect 583444 537820 583446 537840
rect 583390 537784 583446 537820
rect 582838 484608 582894 484664
rect 583390 431604 583392 431624
rect 583392 431604 583444 431624
rect 583444 431604 583446 431624
rect 583390 431568 583446 431604
rect 583390 418276 583392 418296
rect 583392 418276 583444 418296
rect 583444 418276 583446 418296
rect 583390 418240 583446 418276
rect 582746 404912 582802 404968
rect 583390 351908 583392 351928
rect 583392 351908 583444 351928
rect 583444 351908 583446 351928
rect 583390 351872 583446 351908
rect 583390 325252 583392 325272
rect 583392 325252 583444 325272
rect 583444 325252 583446 325272
rect 583390 325216 583446 325252
rect 583390 312060 583392 312080
rect 583392 312060 583444 312080
rect 583444 312060 583446 312080
rect 583390 312024 583446 312060
rect 582654 298696 582710 298752
rect 583298 272212 583300 272232
rect 583300 272212 583352 272232
rect 583352 272212 583354 272232
rect 583298 272176 583354 272212
rect 583206 245556 583208 245576
rect 583208 245556 583260 245576
rect 583260 245556 583262 245576
rect 583206 245520 583262 245556
rect 583114 232364 583116 232384
rect 583116 232364 583168 232384
rect 583168 232364 583170 232384
rect 583114 232328 583170 232364
rect 583022 205708 583024 205728
rect 583024 205708 583076 205728
rect 583076 205708 583078 205728
rect 583022 205672 583078 205708
rect 582930 192516 582932 192536
rect 582932 192516 582984 192536
rect 582984 192516 582986 192536
rect 582930 192480 582986 192516
rect 582838 179188 582840 179208
rect 582840 179188 582892 179208
rect 582892 179188 582894 179208
rect 582838 179152 582894 179188
rect 582746 165860 582748 165880
rect 582748 165860 582800 165880
rect 582800 165860 582802 165880
rect 582746 165824 582802 165860
rect 582654 152668 582656 152688
rect 582656 152668 582708 152688
rect 582708 152668 582710 152688
rect 582654 152632 582710 152668
rect 582654 126012 582656 126032
rect 582656 126012 582708 126032
rect 582708 126012 582710 126032
rect 582654 125976 582710 126012
rect 582654 112820 582656 112840
rect 582656 112820 582708 112840
rect 582708 112820 582710 112840
rect 582654 112784 582710 112820
<< metal3 >>
rect 2037 701722 2103 701725
rect 561857 701722 561923 701725
rect 2037 701720 561923 701722
rect 2037 701664 2042 701720
rect 2098 701664 561862 701720
rect 561918 701664 561923 701720
rect 2037 701662 561923 701664
rect 2037 701659 2103 701662
rect 561857 701659 561923 701662
rect 218053 701586 218119 701589
rect 531589 701586 531655 701589
rect 218053 701584 531655 701586
rect 218053 701528 218058 701584
rect 218114 701528 531594 701584
rect 531650 701528 531655 701584
rect 218053 701526 531655 701528
rect 218053 701523 218119 701526
rect 531589 701523 531655 701526
rect 289 701450 355 701453
rect 526529 701450 526595 701453
rect 289 701448 526595 701450
rect 289 701392 294 701448
rect 350 701392 526534 701448
rect 526590 701392 526595 701448
rect 289 701390 526595 701392
rect 289 701387 355 701390
rect 526529 701387 526595 701390
rect 4521 701314 4587 701317
rect 556797 701314 556863 701317
rect 4521 701312 556863 701314
rect 4521 701256 4526 701312
rect 4582 701256 556802 701312
rect 556858 701256 556863 701312
rect 4521 701254 556863 701256
rect 4521 701251 4587 701254
rect 556797 701251 556863 701254
rect 3417 700362 3483 700365
rect 554773 700362 554839 700365
rect 3417 700360 554839 700362
rect 3417 700304 3422 700360
rect 3478 700304 554778 700360
rect 554834 700304 554839 700360
rect 3417 700302 554839 700304
rect 3417 700299 3483 700302
rect 554773 700299 554839 700302
rect 223849 700226 223915 700229
rect 255262 700226 255268 700228
rect 223849 700224 255268 700226
rect 223849 700168 223854 700224
rect 223910 700168 255268 700224
rect 223849 700166 255268 700168
rect 223849 700163 223915 700166
rect 255262 700164 255268 700166
rect 255332 700164 255338 700228
rect 107745 700090 107811 700093
rect 580625 700090 580691 700093
rect 107745 700088 580691 700090
rect 107745 700032 107750 700088
rect 107806 700032 580630 700088
rect 580686 700032 580691 700088
rect 107745 700030 580691 700032
rect 107745 700027 107811 700030
rect 580625 700027 580691 700030
rect 62389 699954 62455 699957
rect 580441 699954 580507 699957
rect 62389 699952 580507 699954
rect 62389 699896 62394 699952
rect 62450 699896 580446 699952
rect 580502 699896 580507 699952
rect 62389 699894 580507 699896
rect 62389 699891 62455 699894
rect 580441 699891 580507 699894
rect 27061 699818 27127 699821
rect 582465 699818 582531 699821
rect 27061 699816 582531 699818
rect 27061 699760 27066 699816
rect 27122 699760 582470 699816
rect 582526 699760 582531 699816
rect 27061 699758 582531 699760
rect 27061 699755 27127 699758
rect 582465 699755 582531 699758
rect 143349 699140 143415 699141
rect 163589 699140 163655 699141
rect 193765 699140 193831 699141
rect 143349 699136 143396 699140
rect 143460 699138 143466 699140
rect 143349 699080 143354 699136
rect 143349 699076 143396 699080
rect 143460 699078 143506 699138
rect 163589 699136 163636 699140
rect 163700 699138 163706 699140
rect 163589 699080 163594 699136
rect 143460 699076 143466 699078
rect 163589 699076 163636 699080
rect 163700 699078 163746 699138
rect 193765 699136 193812 699140
rect 193876 699138 193882 699140
rect 193765 699080 193770 699136
rect 163700 699076 163706 699078
rect 193765 699076 193812 699080
rect 193876 699078 193922 699138
rect 193876 699076 193882 699078
rect 389398 699076 389404 699140
rect 389468 699138 389474 699140
rect 390093 699138 390159 699141
rect 389468 699136 390159 699138
rect 389468 699080 390098 699136
rect 390154 699080 390159 699136
rect 389468 699078 390159 699080
rect 389468 699076 389474 699078
rect 143349 699075 143415 699076
rect 163589 699075 163655 699076
rect 193765 699075 193831 699076
rect 390093 699075 390159 699078
rect 430614 699076 430620 699140
rect 430684 699138 430690 699140
rect 430757 699138 430823 699141
rect 450721 699140 450787 699141
rect 461025 699140 461091 699141
rect 450670 699138 450676 699140
rect 430684 699136 430823 699138
rect 430684 699080 430762 699136
rect 430818 699080 430823 699136
rect 430684 699078 430823 699080
rect 450630 699078 450676 699138
rect 450740 699136 450787 699140
rect 460974 699138 460980 699140
rect 450782 699080 450787 699136
rect 430684 699076 430690 699078
rect 430757 699075 430823 699078
rect 450670 699076 450676 699078
rect 450740 699076 450787 699080
rect 460934 699078 460980 699138
rect 461044 699136 461091 699140
rect 461086 699080 461091 699136
rect 460974 699076 460980 699078
rect 461044 699076 461091 699080
rect 476062 699076 476068 699140
rect 476132 699138 476138 699140
rect 476205 699138 476271 699141
rect 476132 699136 476271 699138
rect 476132 699080 476210 699136
rect 476266 699080 476271 699136
rect 476132 699078 476271 699080
rect 476132 699076 476138 699078
rect 450721 699075 450787 699076
rect 461025 699075 461091 699076
rect 476205 699075 476271 699078
rect 539910 699076 539916 699140
rect 539980 699138 539986 699140
rect 541341 699138 541407 699141
rect 539980 699136 541407 699138
rect 539980 699080 541346 699136
rect 541402 699080 541407 699136
rect 539980 699078 541407 699080
rect 539980 699076 539986 699078
rect 541341 699075 541407 699078
rect 17217 699002 17283 699005
rect 112989 699004 113055 699005
rect 21582 699002 21588 699004
rect 17217 699000 21588 699002
rect 17217 698944 17222 699000
rect 17278 698944 21588 699000
rect 17217 698942 21588 698944
rect 17217 698939 17283 698942
rect 21582 698940 21588 698942
rect 21652 698940 21658 699004
rect 112989 699000 113036 699004
rect 113100 699002 113106 699004
rect 132677 699002 132743 699005
rect 580257 699002 580323 699005
rect 112989 698944 112994 699000
rect 112989 698940 113036 698944
rect 113100 698942 113146 699002
rect 132677 699000 580323 699002
rect 132677 698944 132682 699000
rect 132738 698944 580262 699000
rect 580318 698944 580323 699000
rect 132677 698942 580323 698944
rect 113100 698940 113106 698942
rect 112989 698939 113055 698940
rect 132677 698939 132743 698942
rect 580257 698939 580323 698942
rect 258574 698730 258580 698732
rect 258030 698670 258580 698730
rect 255262 698532 255268 698596
rect 255332 698594 255338 698596
rect 258030 698594 258090 698670
rect 258574 698668 258580 698670
rect 258644 698668 258650 698732
rect 267774 698668 267780 698732
rect 267844 698730 267850 698732
rect 383510 698730 383516 698732
rect 267844 698670 383516 698730
rect 267844 698668 267850 698670
rect 383510 698668 383516 698670
rect 383580 698668 383586 698732
rect 255332 698534 258090 698594
rect 255332 698532 255338 698534
rect 258390 698532 258396 698596
rect 258460 698594 258466 698596
rect 268142 698594 268148 698596
rect 258460 698534 268148 698594
rect 258460 698532 258466 698534
rect 268142 698532 268148 698534
rect 268212 698532 268218 698596
rect 276974 698532 276980 698596
rect 277044 698594 277050 698596
rect 277710 698594 277716 698596
rect 277044 698534 277716 698594
rect 277044 698532 277050 698534
rect 277710 698532 277716 698534
rect 277780 698532 277786 698596
rect 284886 698532 284892 698596
rect 284956 698594 284962 698596
rect 288014 698594 288020 698596
rect 284956 698534 288020 698594
rect 284956 698532 284962 698534
rect 288014 698532 288020 698534
rect 288084 698532 288090 698596
rect 296294 698532 296300 698596
rect 296364 698594 296370 698596
rect 297030 698594 297036 698596
rect 296364 698534 297036 698594
rect 296364 698532 296370 698534
rect 297030 698532 297036 698534
rect 297100 698532 297106 698596
rect 304206 698532 304212 698596
rect 304276 698594 304282 698596
rect 307334 698594 307340 698596
rect 304276 698534 307340 698594
rect 304276 698532 304282 698534
rect 307334 698532 307340 698534
rect 307404 698532 307410 698596
rect 315614 698532 315620 698596
rect 315684 698594 315690 698596
rect 316350 698594 316356 698596
rect 315684 698534 316356 698594
rect 315684 698532 315690 698534
rect 316350 698532 316356 698534
rect 316420 698532 316426 698596
rect 323526 698532 323532 698596
rect 323596 698594 323602 698596
rect 326654 698594 326660 698596
rect 323596 698534 326660 698594
rect 323596 698532 323602 698534
rect 326654 698532 326660 698534
rect 326724 698532 326730 698596
rect 334934 698532 334940 698596
rect 335004 698594 335010 698596
rect 335670 698594 335676 698596
rect 335004 698534 335676 698594
rect 335004 698532 335010 698534
rect 335670 698532 335676 698534
rect 335740 698532 335746 698596
rect 342846 698532 342852 698596
rect 342916 698594 342922 698596
rect 345974 698594 345980 698596
rect 342916 698534 345980 698594
rect 342916 698532 342922 698534
rect 345974 698532 345980 698534
rect 346044 698532 346050 698596
rect 354254 698532 354260 698596
rect 354324 698594 354330 698596
rect 354990 698594 354996 698596
rect 354324 698534 354996 698594
rect 354324 698532 354330 698534
rect 354990 698532 354996 698534
rect 355060 698532 355066 698596
rect 362166 698532 362172 698596
rect 362236 698594 362242 698596
rect 365294 698594 365300 698596
rect 362236 698534 365300 698594
rect 362236 698532 362242 698534
rect 365294 698532 365300 698534
rect 365364 698532 365370 698596
rect 373574 698532 373580 698596
rect 373644 698594 373650 698596
rect 374310 698594 374316 698596
rect 373644 698534 374316 698594
rect 373644 698532 373650 698534
rect 374310 698532 374316 698534
rect 374380 698532 374386 698596
rect 382958 698532 382964 698596
rect 383028 698594 383034 698596
rect 389398 698594 389404 698596
rect 383028 698534 389404 698594
rect 383028 698532 383034 698534
rect 389398 698532 389404 698534
rect 389468 698532 389474 698596
rect 3509 698458 3575 698461
rect 539910 698458 539916 698460
rect 3509 698456 539916 698458
rect 3509 698400 3514 698456
rect 3570 698400 539916 698456
rect 3509 698398 539916 698400
rect 3509 698395 3575 698398
rect 539910 698396 539916 698398
rect 539980 698396 539986 698460
rect 21582 698260 21588 698324
rect 21652 698322 21658 698324
rect 267774 698322 267780 698324
rect 21652 698262 267780 698322
rect 21652 698260 21658 698262
rect 267774 698260 267780 698262
rect 267844 698260 267850 698324
rect 267958 698260 267964 698324
rect 268028 698322 268034 698324
rect 277158 698322 277164 698324
rect 268028 698262 277164 698322
rect 268028 698260 268034 698262
rect 277158 698260 277164 698262
rect 277228 698260 277234 698324
rect 277526 698260 277532 698324
rect 277596 698322 277602 698324
rect 284886 698322 284892 698324
rect 277596 698262 284892 698322
rect 277596 698260 277602 698262
rect 284886 698260 284892 698262
rect 284956 698260 284962 698324
rect 286726 698260 286732 698324
rect 286796 698322 286802 698324
rect 287830 698322 287836 698324
rect 286796 698262 287836 698322
rect 286796 698260 286802 698262
rect 287830 698260 287836 698262
rect 287900 698260 287906 698324
rect 288014 698260 288020 698324
rect 288084 698322 288090 698324
rect 296478 698322 296484 698324
rect 288084 698262 296484 698322
rect 288084 698260 288090 698262
rect 296478 698260 296484 698262
rect 296548 698260 296554 698324
rect 296846 698260 296852 698324
rect 296916 698322 296922 698324
rect 304206 698322 304212 698324
rect 296916 698262 304212 698322
rect 296916 698260 296922 698262
rect 304206 698260 304212 698262
rect 304276 698260 304282 698324
rect 306046 698260 306052 698324
rect 306116 698322 306122 698324
rect 307150 698322 307156 698324
rect 306116 698262 307156 698322
rect 306116 698260 306122 698262
rect 307150 698260 307156 698262
rect 307220 698260 307226 698324
rect 307334 698260 307340 698324
rect 307404 698322 307410 698324
rect 315798 698322 315804 698324
rect 307404 698262 315804 698322
rect 307404 698260 307410 698262
rect 315798 698260 315804 698262
rect 315868 698260 315874 698324
rect 316166 698260 316172 698324
rect 316236 698322 316242 698324
rect 323526 698322 323532 698324
rect 316236 698262 323532 698322
rect 316236 698260 316242 698262
rect 323526 698260 323532 698262
rect 323596 698260 323602 698324
rect 325366 698260 325372 698324
rect 325436 698322 325442 698324
rect 326470 698322 326476 698324
rect 325436 698262 326476 698322
rect 325436 698260 325442 698262
rect 326470 698260 326476 698262
rect 326540 698260 326546 698324
rect 326654 698260 326660 698324
rect 326724 698322 326730 698324
rect 335118 698322 335124 698324
rect 326724 698262 335124 698322
rect 326724 698260 326730 698262
rect 335118 698260 335124 698262
rect 335188 698260 335194 698324
rect 335486 698260 335492 698324
rect 335556 698322 335562 698324
rect 342846 698322 342852 698324
rect 335556 698262 342852 698322
rect 335556 698260 335562 698262
rect 342846 698260 342852 698262
rect 342916 698260 342922 698324
rect 344686 698260 344692 698324
rect 344756 698322 344762 698324
rect 345790 698322 345796 698324
rect 344756 698262 345796 698322
rect 344756 698260 344762 698262
rect 345790 698260 345796 698262
rect 345860 698260 345866 698324
rect 345974 698260 345980 698324
rect 346044 698322 346050 698324
rect 354438 698322 354444 698324
rect 346044 698262 354444 698322
rect 346044 698260 346050 698262
rect 354438 698260 354444 698262
rect 354508 698260 354514 698324
rect 354806 698260 354812 698324
rect 354876 698322 354882 698324
rect 362166 698322 362172 698324
rect 354876 698262 362172 698322
rect 354876 698260 354882 698262
rect 362166 698260 362172 698262
rect 362236 698260 362242 698324
rect 364006 698260 364012 698324
rect 364076 698322 364082 698324
rect 365110 698322 365116 698324
rect 364076 698262 365116 698322
rect 364076 698260 364082 698262
rect 365110 698260 365116 698262
rect 365180 698260 365186 698324
rect 365294 698260 365300 698324
rect 365364 698322 365370 698324
rect 373758 698322 373764 698324
rect 365364 698262 373764 698322
rect 365364 698260 365370 698262
rect 373758 698260 373764 698262
rect 373828 698260 373834 698324
rect 374126 698260 374132 698324
rect 374196 698322 374202 698324
rect 383142 698322 383148 698324
rect 374196 698262 383148 698322
rect 374196 698260 374202 698262
rect 383142 698260 383148 698262
rect 383212 698260 383218 698324
rect 383510 698260 383516 698324
rect 383580 698322 383586 698324
rect 582373 698322 582439 698325
rect 383580 698320 582439 698322
rect 383580 698264 582378 698320
rect 582434 698264 582439 698320
rect 383580 698262 582439 698264
rect 383580 698260 383586 698262
rect 582373 698259 582439 698262
rect 1945 698186 2011 698189
rect 286174 698186 286180 698188
rect 1945 698184 286180 698186
rect 1945 698128 1950 698184
rect 2006 698128 286180 698184
rect 1945 698126 286180 698128
rect 1945 698123 2011 698126
rect 286174 698124 286180 698126
rect 286244 698124 286250 698188
rect 286726 698124 286732 698188
rect 286796 698186 286802 698188
rect 305494 698186 305500 698188
rect 286796 698126 305500 698186
rect 286796 698124 286802 698126
rect 305494 698124 305500 698126
rect 305564 698124 305570 698188
rect 306046 698124 306052 698188
rect 306116 698186 306122 698188
rect 324814 698186 324820 698188
rect 306116 698126 324820 698186
rect 306116 698124 306122 698126
rect 324814 698124 324820 698126
rect 324884 698124 324890 698188
rect 325366 698124 325372 698188
rect 325436 698186 325442 698188
rect 344134 698186 344140 698188
rect 325436 698126 344140 698186
rect 325436 698124 325442 698126
rect 344134 698124 344140 698126
rect 344204 698124 344210 698188
rect 344686 698124 344692 698188
rect 344756 698186 344762 698188
rect 363454 698186 363460 698188
rect 344756 698126 363460 698186
rect 344756 698124 344762 698126
rect 363454 698124 363460 698126
rect 363524 698124 363530 698188
rect 364006 698124 364012 698188
rect 364076 698186 364082 698188
rect 430614 698186 430620 698188
rect 364076 698126 430620 698186
rect 364076 698124 364082 698126
rect 430614 698124 430620 698126
rect 430684 698124 430690 698188
rect 143390 697988 143396 698052
rect 143460 698050 143466 698052
rect 143460 697990 277410 698050
rect 143460 697988 143466 697990
rect 2681 697914 2747 697917
rect 267774 697914 267780 697916
rect 2681 697912 267780 697914
rect 2681 697856 2686 697912
rect 2742 697856 267780 697912
rect 2681 697854 267780 697856
rect 2681 697851 2747 697854
rect 267774 697852 267780 697854
rect 267844 697852 267850 697916
rect 268142 697852 268148 697916
rect 268212 697914 268218 697916
rect 276974 697914 276980 697916
rect 268212 697854 276980 697914
rect 268212 697852 268218 697854
rect 276974 697852 276980 697854
rect 277044 697852 277050 697916
rect 277350 697914 277410 697990
rect 277710 697988 277716 698052
rect 277780 698050 277786 698052
rect 286358 698050 286364 698052
rect 277780 697990 286364 698050
rect 277780 697988 277786 697990
rect 286358 697988 286364 697990
rect 286428 697988 286434 698052
rect 287654 697990 296730 698050
rect 287654 697914 287714 697990
rect 277350 697854 287714 697914
rect 287830 697852 287836 697916
rect 287900 697914 287906 697916
rect 296294 697914 296300 697916
rect 287900 697854 296300 697914
rect 287900 697852 287906 697854
rect 296294 697852 296300 697854
rect 296364 697852 296370 697916
rect 296670 697914 296730 697990
rect 297030 697988 297036 698052
rect 297100 698050 297106 698052
rect 305678 698050 305684 698052
rect 297100 697990 305684 698050
rect 297100 697988 297106 697990
rect 305678 697988 305684 697990
rect 305748 697988 305754 698052
rect 306974 697990 316050 698050
rect 306974 697914 307034 697990
rect 296670 697854 307034 697914
rect 307150 697852 307156 697916
rect 307220 697914 307226 697916
rect 315614 697914 315620 697916
rect 307220 697854 315620 697914
rect 307220 697852 307226 697854
rect 315614 697852 315620 697854
rect 315684 697852 315690 697916
rect 315990 697914 316050 697990
rect 316350 697988 316356 698052
rect 316420 698050 316426 698052
rect 324998 698050 325004 698052
rect 316420 697990 325004 698050
rect 316420 697988 316426 697990
rect 324998 697988 325004 697990
rect 325068 697988 325074 698052
rect 326294 697990 335370 698050
rect 326294 697914 326354 697990
rect 315990 697854 326354 697914
rect 326470 697852 326476 697916
rect 326540 697914 326546 697916
rect 334934 697914 334940 697916
rect 326540 697854 334940 697914
rect 326540 697852 326546 697854
rect 334934 697852 334940 697854
rect 335004 697852 335010 697916
rect 335310 697914 335370 697990
rect 335670 697988 335676 698052
rect 335740 698050 335746 698052
rect 344318 698050 344324 698052
rect 335740 697990 344324 698050
rect 335740 697988 335746 697990
rect 344318 697988 344324 697990
rect 344388 697988 344394 698052
rect 345614 697990 354690 698050
rect 345614 697914 345674 697990
rect 335310 697854 345674 697914
rect 345790 697852 345796 697916
rect 345860 697914 345866 697916
rect 354254 697914 354260 697916
rect 345860 697854 354260 697914
rect 345860 697852 345866 697854
rect 354254 697852 354260 697854
rect 354324 697852 354330 697916
rect 354630 697914 354690 697990
rect 354990 697988 354996 698052
rect 355060 698050 355066 698052
rect 363638 698050 363644 698052
rect 355060 697990 363644 698050
rect 355060 697988 355066 697990
rect 363638 697988 363644 697990
rect 363708 697988 363714 698052
rect 364934 697990 374010 698050
rect 364934 697914 364994 697990
rect 354630 697854 364994 697914
rect 365110 697852 365116 697916
rect 365180 697914 365186 697916
rect 373574 697914 373580 697916
rect 365180 697854 373580 697914
rect 365180 697852 365186 697854
rect 373574 697852 373580 697854
rect 373644 697852 373650 697916
rect 373950 697914 374010 697990
rect 374310 697988 374316 698052
rect 374380 698050 374386 698052
rect 382958 698050 382964 698052
rect 374380 697990 382964 698050
rect 374380 697988 374386 697990
rect 382958 697988 382964 697990
rect 383028 697988 383034 698052
rect 582741 698050 582807 698053
rect 383334 698048 582807 698050
rect 383334 697992 582746 698048
rect 582802 697992 582807 698048
rect 383334 697990 582807 697992
rect 383334 697914 383394 697990
rect 582741 697987 582807 697990
rect 373950 697854 383394 697914
rect 383510 697852 383516 697916
rect 383580 697914 383586 697916
rect 450670 697914 450676 697916
rect 383580 697854 450676 697914
rect 383580 697852 383586 697854
rect 450670 697852 450676 697854
rect 450740 697852 450746 697916
rect 2497 697778 2563 697781
rect 460974 697778 460980 697780
rect 2497 697776 460980 697778
rect 2497 697720 2502 697776
rect 2558 697720 460980 697776
rect 2497 697718 460980 697720
rect 2497 697715 2563 697718
rect 460974 697716 460980 697718
rect 461044 697716 461050 697780
rect 113030 697580 113036 697644
rect 113100 697642 113106 697644
rect 582649 697642 582715 697645
rect 113100 697640 582715 697642
rect 113100 697584 582654 697640
rect 582710 697584 582715 697640
rect 113100 697582 582715 697584
rect 113100 697580 113106 697582
rect 582649 697579 582715 697582
rect 2313 697506 2379 697509
rect 476062 697506 476068 697508
rect 2313 697504 476068 697506
rect -960 697220 480 697460
rect 2313 697448 2318 697504
rect 2374 697448 476068 697504
rect 2313 697446 476068 697448
rect 2313 697443 2379 697446
rect 476062 697444 476068 697446
rect 476132 697444 476138 697508
rect 163630 697308 163636 697372
rect 163700 697370 163706 697372
rect 582833 697370 582899 697373
rect 163700 697368 582899 697370
rect 163700 697312 582838 697368
rect 582894 697312 582899 697368
rect 163700 697310 582899 697312
rect 163700 697308 163706 697310
rect 582833 697307 582899 697310
rect 193806 697172 193812 697236
rect 193876 697234 193882 697236
rect 579889 697234 579955 697237
rect 583520 697234 584960 697324
rect 193876 697232 579955 697234
rect 193876 697176 579894 697232
rect 579950 697176 579955 697232
rect 193876 697174 579955 697176
rect 193876 697172 193882 697174
rect 579889 697171 579955 697174
rect 580214 697174 584960 697234
rect 841 697098 907 697101
rect 258022 697098 258028 697100
rect 841 697096 258028 697098
rect 841 697040 846 697096
rect 902 697040 258028 697096
rect 841 697038 258028 697040
rect 841 697035 907 697038
rect 258022 697036 258028 697038
rect 258092 697036 258098 697100
rect 258574 697036 258580 697100
rect 258644 697098 258650 697100
rect 580214 697098 580274 697174
rect 258644 697038 580274 697098
rect 583520 697084 584960 697174
rect 258644 697036 258650 697038
rect 579889 696962 579955 696965
rect 582925 696962 582991 696965
rect 579889 696960 582991 696962
rect 579889 696904 579894 696960
rect 579950 696904 582930 696960
rect 582986 696904 582991 696960
rect 579889 696902 582991 696904
rect 579889 696899 579955 696902
rect 582925 696899 582991 696902
rect -960 684314 480 684404
rect 1485 684314 1551 684317
rect -960 684312 1551 684314
rect -960 684256 1490 684312
rect 1546 684256 1551 684312
rect -960 684254 1551 684256
rect -960 684164 480 684254
rect 1485 684251 1551 684254
rect 579981 683906 580047 683909
rect 583520 683906 584960 683996
rect 579981 683904 584960 683906
rect 579981 683848 579986 683904
rect 580042 683848 584960 683904
rect 579981 683846 584960 683848
rect 579981 683843 580047 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3693 671258 3759 671261
rect -960 671256 3759 671258
rect -960 671200 3698 671256
rect 3754 671200 3759 671256
rect -960 671198 3759 671200
rect -960 671108 480 671198
rect 3693 671195 3759 671198
rect 581545 670714 581611 670717
rect 583520 670714 584960 670804
rect 581545 670712 584960 670714
rect 581545 670656 581550 670712
rect 581606 670656 584960 670712
rect 581545 670654 584960 670656
rect 581545 670651 581611 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 1577 658202 1643 658205
rect -960 658200 1643 658202
rect -960 658144 1582 658200
rect 1638 658144 1643 658200
rect -960 658142 1643 658144
rect -960 658052 480 658142
rect 1577 658139 1643 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 579153 644058 579219 644061
rect 583520 644058 584960 644148
rect 579153 644056 584960 644058
rect 579153 644000 579158 644056
rect 579214 644000 584960 644056
rect 579153 643998 584960 644000
rect 579153 643995 579219 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 1669 632090 1735 632093
rect -960 632088 1735 632090
rect -960 632032 1674 632088
rect 1730 632032 1735 632088
rect -960 632030 1735 632032
rect -960 631940 480 632030
rect 1669 632027 1735 632030
rect 580073 630866 580139 630869
rect 583520 630866 584960 630956
rect 580073 630864 584960 630866
rect 580073 630808 580078 630864
rect 580134 630808 584960 630864
rect 580073 630806 584960 630808
rect 580073 630803 580139 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3049 619170 3115 619173
rect -960 619168 3115 619170
rect -960 619112 3054 619168
rect 3110 619112 3115 619168
rect -960 619110 3115 619112
rect -960 619020 480 619110
rect 3049 619107 3115 619110
rect 582281 617538 582347 617541
rect 583520 617538 584960 617628
rect 582281 617536 584960 617538
rect 582281 617480 582286 617536
rect 582342 617480 584960 617536
rect 582281 617478 584960 617480
rect 582281 617475 582347 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 841 606114 907 606117
rect -960 606112 907 606114
rect -960 606056 846 606112
rect 902 606056 907 606112
rect -960 606054 907 606056
rect -960 605964 480 606054
rect 841 606051 907 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 582925 591018 582991 591021
rect 583520 591018 584960 591108
rect 582925 591016 584960 591018
rect 582925 590960 582930 591016
rect 582986 590960 584960 591016
rect 582925 590958 584960 590960
rect 582925 590955 582991 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 1761 580002 1827 580005
rect -960 580000 1827 580002
rect -960 579944 1766 580000
rect 1822 579944 1827 580000
rect -960 579942 1827 579944
rect -960 579852 480 579942
rect 1761 579939 1827 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 582189 564362 582255 564365
rect 583520 564362 584960 564452
rect 582189 564360 584960 564362
rect 582189 564304 582194 564360
rect 582250 564304 584960 564360
rect 582189 564302 584960 564304
rect 582189 564299 582255 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 749 553890 815 553893
rect -960 553888 815 553890
rect -960 553832 754 553888
rect 810 553832 815 553888
rect -960 553830 815 553832
rect -960 553740 480 553830
rect 749 553827 815 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583385 537842 583451 537845
rect 583520 537842 584960 537932
rect 583385 537840 584960 537842
rect 583385 537784 583390 537840
rect 583446 537784 584960 537840
rect 583385 537782 584960 537784
rect 583385 537779 583451 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 1853 527914 1919 527917
rect -960 527912 1919 527914
rect -960 527856 1858 527912
rect 1914 527856 1919 527912
rect -960 527854 1919 527856
rect -960 527764 480 527854
rect 1853 527851 1919 527854
rect 580901 524514 580967 524517
rect 583520 524514 584960 524604
rect 580901 524512 584960 524514
rect 580901 524456 580906 524512
rect 580962 524456 584960 524512
rect 580901 524454 584960 524456
rect 580901 524451 580967 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3141 514858 3207 514861
rect -960 514856 3207 514858
rect -960 514800 3146 514856
rect 3202 514800 3207 514856
rect -960 514798 3207 514800
rect -960 514708 480 514798
rect 3141 514795 3207 514798
rect 582097 511322 582163 511325
rect 583520 511322 584960 511412
rect 582097 511320 584960 511322
rect 582097 511264 582102 511320
rect 582158 511264 584960 511320
rect 582097 511262 584960 511264
rect 582097 511259 582163 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2589 501802 2655 501805
rect -960 501800 2655 501802
rect -960 501744 2594 501800
rect 2650 501744 2655 501800
rect -960 501742 2655 501744
rect -960 501652 480 501742
rect 2589 501739 2655 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 582833 484666 582899 484669
rect 583520 484666 584960 484756
rect 582833 484664 584960 484666
rect 582833 484608 582838 484664
rect 582894 484608 584960 484664
rect 582833 484606 584960 484608
rect 582833 484603 582899 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 1945 475690 2011 475693
rect -960 475688 2011 475690
rect -960 475632 1950 475688
rect 2006 475632 2011 475688
rect -960 475630 2011 475632
rect -960 475540 480 475630
rect 1945 475627 2011 475630
rect 580809 471474 580875 471477
rect 583520 471474 584960 471564
rect 580809 471472 584960 471474
rect 580809 471416 580814 471472
rect 580870 471416 584960 471472
rect 580809 471414 584960 471416
rect 580809 471411 580875 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 582005 458146 582071 458149
rect 583520 458146 584960 458236
rect 582005 458144 584960 458146
rect 582005 458088 582010 458144
rect 582066 458088 584960 458144
rect 582005 458086 584960 458088
rect 582005 458083 582071 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 657 449578 723 449581
rect -960 449576 723 449578
rect -960 449520 662 449576
rect 718 449520 723 449576
rect -960 449518 723 449520
rect -960 449428 480 449518
rect 657 449515 723 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583385 431626 583451 431629
rect 583520 431626 584960 431716
rect 583385 431624 584960 431626
rect 583385 431568 583390 431624
rect 583446 431568 584960 431624
rect 583385 431566 584960 431568
rect 583385 431563 583451 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2405 423602 2471 423605
rect -960 423600 2471 423602
rect -960 423544 2410 423600
rect 2466 423544 2471 423600
rect -960 423542 2471 423544
rect -960 423452 480 423542
rect 2405 423539 2471 423542
rect 583385 418298 583451 418301
rect 583520 418298 584960 418388
rect 583385 418296 584960 418298
rect 583385 418240 583390 418296
rect 583446 418240 584960 418296
rect 583385 418238 584960 418240
rect 583385 418235 583451 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 582741 404970 582807 404973
rect 583520 404970 584960 405060
rect 582741 404968 584960 404970
rect 582741 404912 582746 404968
rect 582802 404912 584960 404968
rect 582741 404910 584960 404912
rect 582741 404907 582807 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 2681 397490 2747 397493
rect -960 397488 2747 397490
rect -960 397432 2686 397488
rect 2742 397432 2747 397488
rect -960 397430 2747 397432
rect -960 397340 480 397430
rect 2681 397427 2747 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580717 378450 580783 378453
rect 583520 378450 584960 378540
rect 580717 378448 584960 378450
rect 580717 378392 580722 378448
rect 580778 378392 584960 378448
rect 580717 378390 584960 378392
rect 580717 378387 580783 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2497 371378 2563 371381
rect -960 371376 2563 371378
rect -960 371320 2502 371376
rect 2558 371320 2563 371376
rect -960 371318 2563 371320
rect -960 371228 480 371318
rect 2497 371315 2563 371318
rect 580533 365122 580599 365125
rect 583520 365122 584960 365212
rect 580533 365120 584960 365122
rect 580533 365064 580538 365120
rect 580594 365064 584960 365120
rect 580533 365062 584960 365064
rect 580533 365059 580599 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 4797 358458 4863 358461
rect -960 358456 4863 358458
rect -960 358400 4802 358456
rect 4858 358400 4863 358456
rect -960 358398 4863 358400
rect -960 358308 480 358398
rect 4797 358395 4863 358398
rect 583385 351930 583451 351933
rect 583520 351930 584960 352020
rect 583385 351928 584960 351930
rect 583385 351872 583390 351928
rect 583446 351872 584960 351928
rect 583385 351870 584960 351872
rect 583385 351867 583451 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 565 345402 631 345405
rect -960 345400 631 345402
rect -960 345344 570 345400
rect 626 345344 631 345400
rect -960 345342 631 345344
rect -960 345252 480 345342
rect 565 345339 631 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583385 325274 583451 325277
rect 583520 325274 584960 325364
rect 583385 325272 584960 325274
rect 583385 325216 583390 325272
rect 583446 325216 584960 325272
rect 583385 325214 584960 325216
rect 583385 325211 583451 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2313 319290 2379 319293
rect -960 319288 2379 319290
rect -960 319232 2318 319288
rect 2374 319232 2379 319288
rect -960 319230 2379 319232
rect -960 319140 480 319230
rect 2313 319227 2379 319230
rect 583385 312082 583451 312085
rect 583520 312082 584960 312172
rect 583385 312080 584960 312082
rect 583385 312024 583390 312080
rect 583446 312024 584960 312080
rect 583385 312022 584960 312024
rect 583385 312019 583451 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 2773 306234 2839 306237
rect -960 306232 2839 306234
rect -960 306176 2778 306232
rect 2834 306176 2839 306232
rect -960 306174 2839 306176
rect -960 306084 480 306174
rect 2773 306171 2839 306174
rect 582649 298754 582715 298757
rect 583520 298754 584960 298844
rect 582649 298752 584960 298754
rect 582649 298696 582654 298752
rect 582710 298696 584960 298752
rect 582649 298694 584960 298696
rect 582649 298691 582715 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 4061 293178 4127 293181
rect -960 293176 4127 293178
rect -960 293120 4066 293176
rect 4122 293120 4127 293176
rect -960 293118 4127 293120
rect -960 293028 480 293118
rect 4061 293115 4127 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583293 272234 583359 272237
rect 583520 272234 584960 272324
rect 583293 272232 584960 272234
rect 583293 272176 583298 272232
rect 583354 272176 584960 272232
rect 583293 272174 584960 272176
rect 583293 272171 583359 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 565 267202 631 267205
rect -960 267200 631 267202
rect -960 267144 570 267200
rect 626 267144 631 267200
rect -960 267142 631 267144
rect -960 267052 480 267142
rect 565 267139 631 267142
rect 580625 258906 580691 258909
rect 583520 258906 584960 258996
rect 580625 258904 584960 258906
rect 580625 258848 580630 258904
rect 580686 258848 584960 258904
rect 580625 258846 584960 258848
rect 580625 258843 580691 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3233 254146 3299 254149
rect -960 254144 3299 254146
rect -960 254088 3238 254144
rect 3294 254088 3299 254144
rect -960 254086 3299 254088
rect -960 253996 480 254086
rect 3233 254083 3299 254086
rect 583201 245578 583267 245581
rect 583520 245578 584960 245668
rect 583201 245576 584960 245578
rect 583201 245520 583206 245576
rect 583262 245520 584960 245576
rect 583201 245518 584960 245520
rect 583201 245515 583267 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2221 241090 2287 241093
rect -960 241088 2287 241090
rect -960 241032 2226 241088
rect 2282 241032 2287 241088
rect -960 241030 2287 241032
rect -960 240940 480 241030
rect 2221 241027 2287 241030
rect 583109 232386 583175 232389
rect 583520 232386 584960 232476
rect 583109 232384 584960 232386
rect 583109 232328 583114 232384
rect 583170 232328 584960 232384
rect 583109 232326 584960 232328
rect 583109 232323 583175 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 581913 219058 581979 219061
rect 583520 219058 584960 219148
rect 581913 219056 584960 219058
rect 581913 219000 581918 219056
rect 581974 219000 584960 219056
rect 581913 218998 584960 219000
rect 581913 218995 581979 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 565 214978 631 214981
rect -960 214976 631 214978
rect -960 214920 570 214976
rect 626 214920 631 214976
rect -960 214918 631 214920
rect -960 214828 480 214918
rect 565 214915 631 214918
rect 583017 205730 583083 205733
rect 583520 205730 584960 205820
rect 583017 205728 584960 205730
rect 583017 205672 583022 205728
rect 583078 205672 584960 205728
rect 583017 205670 584960 205672
rect 583017 205667 583083 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3969 201922 4035 201925
rect -960 201920 4035 201922
rect -960 201864 3974 201920
rect 4030 201864 4035 201920
rect -960 201862 4035 201864
rect -960 201772 480 201862
rect 3969 201859 4035 201862
rect 582925 192538 582991 192541
rect 583520 192538 584960 192628
rect 582925 192536 584960 192538
rect 582925 192480 582930 192536
rect 582986 192480 584960 192536
rect 582925 192478 584960 192480
rect 582925 192475 582991 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3877 188866 3943 188869
rect -960 188864 3943 188866
rect -960 188808 3882 188864
rect 3938 188808 3943 188864
rect -960 188806 3943 188808
rect -960 188716 480 188806
rect 3877 188803 3943 188806
rect 582833 179210 582899 179213
rect 583520 179210 584960 179300
rect 582833 179208 584960 179210
rect 582833 179152 582838 179208
rect 582894 179152 584960 179208
rect 582833 179150 584960 179152
rect 582833 179147 582899 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 582741 165882 582807 165885
rect 583520 165882 584960 165972
rect 582741 165880 584960 165882
rect 582741 165824 582746 165880
rect 582802 165824 584960 165880
rect 582741 165822 584960 165824
rect 582741 165819 582807 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2129 162890 2195 162893
rect -960 162888 2195 162890
rect -960 162832 2134 162888
rect 2190 162832 2195 162888
rect -960 162830 2195 162832
rect -960 162740 480 162830
rect 2129 162827 2195 162830
rect 582649 152690 582715 152693
rect 583520 152690 584960 152780
rect 582649 152688 584960 152690
rect 582649 152632 582654 152688
rect 582710 152632 584960 152688
rect 582649 152630 584960 152632
rect 582649 152627 582715 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3785 149834 3851 149837
rect -960 149832 3851 149834
rect -960 149776 3790 149832
rect 3846 149776 3851 149832
rect -960 149774 3851 149776
rect -960 149684 480 149774
rect 3785 149771 3851 149774
rect 580441 139362 580507 139365
rect 583520 139362 584960 139452
rect 580441 139360 584960 139362
rect 580441 139304 580446 139360
rect 580502 139304 584960 139360
rect 580441 139302 584960 139304
rect 580441 139299 580507 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 565 136778 631 136781
rect -960 136776 631 136778
rect -960 136720 570 136776
rect 626 136720 631 136776
rect -960 136718 631 136720
rect -960 136628 480 136718
rect 565 136715 631 136718
rect 582649 126034 582715 126037
rect 583520 126034 584960 126124
rect 582649 126032 584960 126034
rect 582649 125976 582654 126032
rect 582710 125976 584960 126032
rect 582649 125974 584960 125976
rect 582649 125971 582715 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 582649 112842 582715 112845
rect 583520 112842 584960 112932
rect 582649 112840 584960 112842
rect 582649 112784 582654 112840
rect 582710 112784 584960 112840
rect 582649 112782 584960 112784
rect 582649 112779 582715 112782
rect 583520 112692 584960 112782
rect 197 111210 263 111213
rect 197 111208 306 111210
rect 197 111152 202 111208
rect 258 111152 306 111208
rect 197 111147 306 111152
rect 246 110802 306 111147
rect 246 110756 674 110802
rect -960 110742 674 110756
rect -960 110666 480 110742
rect 614 110666 674 110742
rect -960 110606 674 110666
rect -960 110516 480 110606
rect 580349 99514 580415 99517
rect 583520 99514 584960 99604
rect 580349 99512 584960 99514
rect 580349 99456 580354 99512
rect 580410 99456 584960 99512
rect 580349 99454 584960 99456
rect 580349 99451 580415 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3601 97610 3667 97613
rect -960 97608 3667 97610
rect -960 97552 3606 97608
rect 3662 97552 3667 97608
rect -960 97550 3667 97552
rect -960 97460 480 97550
rect 3601 97547 3667 97550
rect 581821 86186 581887 86189
rect 583520 86186 584960 86276
rect 581821 86184 584960 86186
rect 581821 86128 581826 86184
rect 581882 86128 584960 86184
rect 581821 86126 584960 86128
rect 581821 86123 581887 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 582465 72994 582531 72997
rect 583520 72994 584960 73084
rect 582465 72992 584960 72994
rect 582465 72936 582470 72992
rect 582526 72936 584960 72992
rect 582465 72934 584960 72936
rect 582465 72931 582531 72934
rect 583520 72844 584960 72934
rect 105 71906 171 71909
rect 62 71904 171 71906
rect 62 71848 110 71904
rect 166 71848 171 71904
rect 62 71843 171 71848
rect 62 71770 122 71843
rect 62 71724 674 71770
rect -960 71710 674 71724
rect -960 71634 480 71710
rect 614 71634 674 71710
rect -960 71574 674 71634
rect -960 71484 480 71574
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2037 58578 2103 58581
rect -960 58576 2103 58578
rect -960 58520 2042 58576
rect 2098 58520 2103 58576
rect -960 58518 2103 58520
rect -960 58428 480 58518
rect 2037 58515 2103 58518
rect 581729 46338 581795 46341
rect 583520 46338 584960 46428
rect 581729 46336 584960 46338
rect 581729 46280 581734 46336
rect 581790 46280 584960 46336
rect 581729 46278 584960 46280
rect 581729 46275 581795 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3693 45522 3759 45525
rect -960 45520 3759 45522
rect -960 45464 3698 45520
rect 3754 45464 3759 45520
rect -960 45462 3759 45464
rect -960 45372 480 45462
rect 3693 45459 3759 45462
rect 582465 33146 582531 33149
rect 583520 33146 584960 33236
rect 582465 33144 584960 33146
rect 582465 33088 582470 33144
rect 582526 33088 584960 33144
rect 582465 33086 584960 33088
rect 582465 33083 582531 33086
rect 13 33010 79 33013
rect 13 33008 122 33010
rect 13 32952 18 33008
rect 74 32952 122 33008
rect 583520 32996 584960 33086
rect 13 32947 122 32952
rect 62 32602 122 32947
rect 62 32556 674 32602
rect -960 32542 674 32556
rect -960 32466 480 32542
rect 614 32466 674 32542
rect -960 32406 674 32466
rect -960 32316 480 32406
rect 582373 19818 582439 19821
rect 583520 19818 584960 19908
rect 582373 19816 584960 19818
rect 582373 19760 582378 19816
rect 582434 19760 584960 19816
rect 582373 19758 584960 19760
rect 582373 19755 582439 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 581637 6626 581703 6629
rect 583520 6626 584960 6716
rect 581637 6624 584960 6626
rect -960 6490 480 6580
rect 581637 6568 581642 6624
rect 581698 6568 584960 6624
rect 581637 6566 584960 6568
rect 581637 6563 581703 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 255268 700164 255332 700228
rect 143396 699136 143460 699140
rect 143396 699080 143410 699136
rect 143410 699080 143460 699136
rect 143396 699076 143460 699080
rect 163636 699136 163700 699140
rect 163636 699080 163650 699136
rect 163650 699080 163700 699136
rect 163636 699076 163700 699080
rect 193812 699136 193876 699140
rect 193812 699080 193826 699136
rect 193826 699080 193876 699136
rect 193812 699076 193876 699080
rect 389404 699076 389468 699140
rect 430620 699076 430684 699140
rect 450676 699136 450740 699140
rect 450676 699080 450726 699136
rect 450726 699080 450740 699136
rect 450676 699076 450740 699080
rect 460980 699136 461044 699140
rect 460980 699080 461030 699136
rect 461030 699080 461044 699136
rect 460980 699076 461044 699080
rect 476068 699076 476132 699140
rect 539916 699076 539980 699140
rect 21588 698940 21652 699004
rect 113036 699000 113100 699004
rect 113036 698944 113050 699000
rect 113050 698944 113100 699000
rect 113036 698940 113100 698944
rect 255268 698532 255332 698596
rect 258580 698668 258644 698732
rect 267780 698668 267844 698732
rect 383516 698668 383580 698732
rect 258396 698532 258460 698596
rect 268148 698532 268212 698596
rect 276980 698532 277044 698596
rect 277716 698532 277780 698596
rect 284892 698532 284956 698596
rect 288020 698532 288084 698596
rect 296300 698532 296364 698596
rect 297036 698532 297100 698596
rect 304212 698532 304276 698596
rect 307340 698532 307404 698596
rect 315620 698532 315684 698596
rect 316356 698532 316420 698596
rect 323532 698532 323596 698596
rect 326660 698532 326724 698596
rect 334940 698532 335004 698596
rect 335676 698532 335740 698596
rect 342852 698532 342916 698596
rect 345980 698532 346044 698596
rect 354260 698532 354324 698596
rect 354996 698532 355060 698596
rect 362172 698532 362236 698596
rect 365300 698532 365364 698596
rect 373580 698532 373644 698596
rect 374316 698532 374380 698596
rect 382964 698532 383028 698596
rect 389404 698532 389468 698596
rect 539916 698396 539980 698460
rect 21588 698260 21652 698324
rect 267780 698260 267844 698324
rect 267964 698260 268028 698324
rect 277164 698260 277228 698324
rect 277532 698260 277596 698324
rect 284892 698260 284956 698324
rect 286732 698260 286796 698324
rect 287836 698260 287900 698324
rect 288020 698260 288084 698324
rect 296484 698260 296548 698324
rect 296852 698260 296916 698324
rect 304212 698260 304276 698324
rect 306052 698260 306116 698324
rect 307156 698260 307220 698324
rect 307340 698260 307404 698324
rect 315804 698260 315868 698324
rect 316172 698260 316236 698324
rect 323532 698260 323596 698324
rect 325372 698260 325436 698324
rect 326476 698260 326540 698324
rect 326660 698260 326724 698324
rect 335124 698260 335188 698324
rect 335492 698260 335556 698324
rect 342852 698260 342916 698324
rect 344692 698260 344756 698324
rect 345796 698260 345860 698324
rect 345980 698260 346044 698324
rect 354444 698260 354508 698324
rect 354812 698260 354876 698324
rect 362172 698260 362236 698324
rect 364012 698260 364076 698324
rect 365116 698260 365180 698324
rect 365300 698260 365364 698324
rect 373764 698260 373828 698324
rect 374132 698260 374196 698324
rect 383148 698260 383212 698324
rect 383516 698260 383580 698324
rect 286180 698124 286244 698188
rect 286732 698124 286796 698188
rect 305500 698124 305564 698188
rect 306052 698124 306116 698188
rect 324820 698124 324884 698188
rect 325372 698124 325436 698188
rect 344140 698124 344204 698188
rect 344692 698124 344756 698188
rect 363460 698124 363524 698188
rect 364012 698124 364076 698188
rect 430620 698124 430684 698188
rect 143396 697988 143460 698052
rect 267780 697852 267844 697916
rect 268148 697852 268212 697916
rect 276980 697852 277044 697916
rect 277716 697988 277780 698052
rect 286364 697988 286428 698052
rect 287836 697852 287900 697916
rect 296300 697852 296364 697916
rect 297036 697988 297100 698052
rect 305684 697988 305748 698052
rect 307156 697852 307220 697916
rect 315620 697852 315684 697916
rect 316356 697988 316420 698052
rect 325004 697988 325068 698052
rect 326476 697852 326540 697916
rect 334940 697852 335004 697916
rect 335676 697988 335740 698052
rect 344324 697988 344388 698052
rect 345796 697852 345860 697916
rect 354260 697852 354324 697916
rect 354996 697988 355060 698052
rect 363644 697988 363708 698052
rect 365116 697852 365180 697916
rect 373580 697852 373644 697916
rect 374316 697988 374380 698052
rect 382964 697988 383028 698052
rect 383516 697852 383580 697916
rect 450676 697852 450740 697916
rect 460980 697716 461044 697780
rect 113036 697580 113100 697644
rect 476068 697444 476132 697508
rect 163636 697308 163700 697372
rect 193812 697172 193876 697236
rect 258028 697036 258092 697100
rect 258580 697036 258644 697100
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 701600 2414 704282
rect 5514 701600 6134 706202
rect 9234 701600 9854 708122
rect 12954 701600 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 701600 20414 705242
rect 23514 701600 24134 707162
rect 27234 701600 27854 709082
rect 30954 701600 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 701600 38414 704282
rect 41514 701600 42134 706202
rect 45234 701600 45854 708122
rect 48954 701600 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 701600 56414 705242
rect 59514 701600 60134 707162
rect 63234 701600 63854 709082
rect 66954 701600 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 701600 74414 704282
rect 77514 701600 78134 706202
rect 81234 701600 81854 708122
rect 84954 701600 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 701600 92414 705242
rect 95514 701600 96134 707162
rect 99234 701600 99854 709082
rect 102954 701600 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 701600 110414 704282
rect 113514 701600 114134 706202
rect 117234 701600 117854 708122
rect 120954 701600 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 701600 128414 705242
rect 131514 701600 132134 707162
rect 135234 701600 135854 709082
rect 138954 701600 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 701600 146414 704282
rect 149514 701600 150134 706202
rect 153234 701600 153854 708122
rect 156954 701600 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 701600 164414 705242
rect 167514 701600 168134 707162
rect 171234 701600 171854 709082
rect 174954 701600 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 701600 182414 704282
rect 185514 701600 186134 706202
rect 189234 701600 189854 708122
rect 192954 701600 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 701600 200414 705242
rect 203514 701600 204134 707162
rect 207234 701600 207854 709082
rect 210954 701600 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 701600 218414 704282
rect 221514 701600 222134 706202
rect 225234 701600 225854 708122
rect 228954 701600 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 701600 236414 705242
rect 239514 701600 240134 707162
rect 243234 701600 243854 709082
rect 246954 701600 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 701600 254414 704282
rect 257514 701600 258134 706202
rect 261234 701600 261854 708122
rect 264954 701600 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 701600 272414 705242
rect 275514 701600 276134 707162
rect 279234 701600 279854 709082
rect 282954 701600 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 701600 290414 704282
rect 293514 701600 294134 706202
rect 297234 701600 297854 708122
rect 300954 701600 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 701600 308414 705242
rect 311514 701600 312134 707162
rect 315234 701600 315854 709082
rect 318954 701600 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 701600 326414 704282
rect 329514 701600 330134 706202
rect 333234 701600 333854 708122
rect 336954 701600 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 701600 344414 705242
rect 347514 701600 348134 707162
rect 351234 701600 351854 709082
rect 354954 701600 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 701600 362414 704282
rect 365514 701600 366134 706202
rect 369234 701600 369854 708122
rect 372954 701600 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 701600 380414 705242
rect 383514 701600 384134 707162
rect 387234 701600 387854 709082
rect 390954 701600 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 701600 398414 704282
rect 401514 701600 402134 706202
rect 405234 701600 405854 708122
rect 408954 701600 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 701600 416414 705242
rect 419514 701600 420134 707162
rect 423234 701600 423854 709082
rect 426954 701600 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 701600 434414 704282
rect 437514 701600 438134 706202
rect 441234 701600 441854 708122
rect 444954 701600 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 701600 452414 705242
rect 455514 701600 456134 707162
rect 459234 701600 459854 709082
rect 462954 701600 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 701600 470414 704282
rect 473514 701600 474134 706202
rect 477234 701600 477854 708122
rect 480954 701600 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 701600 488414 705242
rect 491514 701600 492134 707162
rect 495234 701600 495854 709082
rect 498954 701600 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 701600 506414 704282
rect 509514 701600 510134 706202
rect 513234 701600 513854 708122
rect 516954 701600 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 701600 524414 705242
rect 527514 701600 528134 707162
rect 531234 701600 531854 709082
rect 534954 701600 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 701600 542414 704282
rect 545514 701600 546134 706202
rect 549234 701600 549854 708122
rect 552954 701600 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 701600 560414 705242
rect 563514 701600 564134 707162
rect 567234 701600 567854 709082
rect 570954 701600 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 701600 578414 704282
rect 581514 701600 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 255267 700228 255333 700229
rect 255267 700164 255268 700228
rect 255332 700164 255333 700228
rect 255267 700163 255333 700164
rect 143395 699140 143461 699141
rect 143395 699076 143396 699140
rect 143460 699076 143461 699140
rect 143395 699075 143461 699076
rect 163635 699140 163701 699141
rect 163635 699076 163636 699140
rect 163700 699076 163701 699140
rect 163635 699075 163701 699076
rect 193811 699140 193877 699141
rect 193811 699076 193812 699140
rect 193876 699076 193877 699140
rect 193811 699075 193877 699076
rect 21587 699004 21653 699005
rect 21587 698940 21588 699004
rect 21652 698940 21653 699004
rect 21587 698939 21653 698940
rect 113035 699004 113101 699005
rect 113035 698940 113036 699004
rect 113100 698940 113101 699004
rect 113035 698939 113101 698940
rect 21590 698325 21650 698939
rect 21587 698324 21653 698325
rect 21587 698260 21588 698324
rect 21652 698260 21653 698324
rect 21587 698259 21653 698260
rect 113038 697645 113098 698939
rect 143398 698053 143458 699075
rect 143395 698052 143461 698053
rect 143395 697988 143396 698052
rect 143460 697988 143461 698052
rect 143395 697987 143461 697988
rect 113035 697644 113101 697645
rect 113035 697580 113036 697644
rect 113100 697580 113101 697644
rect 113035 697579 113101 697580
rect 163638 697373 163698 699075
rect 163635 697372 163701 697373
rect 163635 697308 163636 697372
rect 163700 697308 163701 697372
rect 163635 697307 163701 697308
rect 193814 697237 193874 699075
rect 255270 698597 255330 700163
rect 389403 699140 389469 699141
rect 389403 699076 389404 699140
rect 389468 699076 389469 699140
rect 389403 699075 389469 699076
rect 430619 699140 430685 699141
rect 430619 699076 430620 699140
rect 430684 699076 430685 699140
rect 430619 699075 430685 699076
rect 450675 699140 450741 699141
rect 450675 699076 450676 699140
rect 450740 699076 450741 699140
rect 450675 699075 450741 699076
rect 460979 699140 461045 699141
rect 460979 699076 460980 699140
rect 461044 699076 461045 699140
rect 460979 699075 461045 699076
rect 476067 699140 476133 699141
rect 476067 699076 476068 699140
rect 476132 699076 476133 699140
rect 476067 699075 476133 699076
rect 539915 699140 539981 699141
rect 539915 699076 539916 699140
rect 539980 699076 539981 699140
rect 539915 699075 539981 699076
rect 258579 698732 258645 698733
rect 258579 698668 258580 698732
rect 258644 698668 258645 698732
rect 258579 698667 258645 698668
rect 267779 698732 267845 698733
rect 267779 698668 267780 698732
rect 267844 698668 267845 698732
rect 267779 698667 267845 698668
rect 383515 698732 383581 698733
rect 383515 698668 383516 698732
rect 383580 698668 383581 698732
rect 383515 698667 383581 698668
rect 255267 698596 255333 698597
rect 255267 698532 255268 698596
rect 255332 698532 255333 698596
rect 255267 698531 255333 698532
rect 258395 698596 258461 698597
rect 258395 698532 258396 698596
rect 258460 698532 258461 698596
rect 258395 698531 258461 698532
rect 258398 697370 258458 698531
rect 258030 697310 258458 697370
rect 193811 697236 193877 697237
rect 193811 697172 193812 697236
rect 193876 697172 193877 697236
rect 193811 697171 193877 697172
rect 258030 697101 258090 697310
rect 258582 697101 258642 698667
rect 267782 698325 267842 698667
rect 268147 698596 268213 698597
rect 268147 698532 268148 698596
rect 268212 698532 268213 698596
rect 268147 698531 268213 698532
rect 276979 698596 277045 698597
rect 276979 698532 276980 698596
rect 277044 698532 277045 698596
rect 276979 698531 277045 698532
rect 277715 698596 277781 698597
rect 277715 698532 277716 698596
rect 277780 698532 277781 698596
rect 277715 698531 277781 698532
rect 284891 698596 284957 698597
rect 284891 698532 284892 698596
rect 284956 698532 284957 698596
rect 284891 698531 284957 698532
rect 288019 698596 288085 698597
rect 288019 698532 288020 698596
rect 288084 698532 288085 698596
rect 288019 698531 288085 698532
rect 296299 698596 296365 698597
rect 296299 698532 296300 698596
rect 296364 698532 296365 698596
rect 296299 698531 296365 698532
rect 297035 698596 297101 698597
rect 297035 698532 297036 698596
rect 297100 698532 297101 698596
rect 297035 698531 297101 698532
rect 304211 698596 304277 698597
rect 304211 698532 304212 698596
rect 304276 698532 304277 698596
rect 304211 698531 304277 698532
rect 307339 698596 307405 698597
rect 307339 698532 307340 698596
rect 307404 698532 307405 698596
rect 307339 698531 307405 698532
rect 315619 698596 315685 698597
rect 315619 698532 315620 698596
rect 315684 698532 315685 698596
rect 315619 698531 315685 698532
rect 316355 698596 316421 698597
rect 316355 698532 316356 698596
rect 316420 698532 316421 698596
rect 316355 698531 316421 698532
rect 323531 698596 323597 698597
rect 323531 698532 323532 698596
rect 323596 698532 323597 698596
rect 323531 698531 323597 698532
rect 326659 698596 326725 698597
rect 326659 698532 326660 698596
rect 326724 698532 326725 698596
rect 326659 698531 326725 698532
rect 334939 698596 335005 698597
rect 334939 698532 334940 698596
rect 335004 698532 335005 698596
rect 334939 698531 335005 698532
rect 335675 698596 335741 698597
rect 335675 698532 335676 698596
rect 335740 698532 335741 698596
rect 335675 698531 335741 698532
rect 342851 698596 342917 698597
rect 342851 698532 342852 698596
rect 342916 698532 342917 698596
rect 342851 698531 342917 698532
rect 345979 698596 346045 698597
rect 345979 698532 345980 698596
rect 346044 698532 346045 698596
rect 345979 698531 346045 698532
rect 354259 698596 354325 698597
rect 354259 698532 354260 698596
rect 354324 698532 354325 698596
rect 354259 698531 354325 698532
rect 354995 698596 355061 698597
rect 354995 698532 354996 698596
rect 355060 698532 355061 698596
rect 354995 698531 355061 698532
rect 362171 698596 362237 698597
rect 362171 698532 362172 698596
rect 362236 698532 362237 698596
rect 362171 698531 362237 698532
rect 365299 698596 365365 698597
rect 365299 698532 365300 698596
rect 365364 698532 365365 698596
rect 365299 698531 365365 698532
rect 373579 698596 373645 698597
rect 373579 698532 373580 698596
rect 373644 698532 373645 698596
rect 373579 698531 373645 698532
rect 374315 698596 374381 698597
rect 374315 698532 374316 698596
rect 374380 698532 374381 698596
rect 374315 698531 374381 698532
rect 382963 698596 383029 698597
rect 382963 698532 382964 698596
rect 383028 698532 383029 698596
rect 382963 698531 383029 698532
rect 267779 698324 267845 698325
rect 267779 698260 267780 698324
rect 267844 698260 267845 698324
rect 267779 698259 267845 698260
rect 267963 698324 268029 698325
rect 267963 698260 267964 698324
rect 268028 698260 268029 698324
rect 267963 698259 268029 698260
rect 267966 698050 268026 698259
rect 267782 697990 268026 698050
rect 267782 697917 267842 697990
rect 268150 697917 268210 698531
rect 276982 697917 277042 698531
rect 277163 698324 277229 698325
rect 277163 698260 277164 698324
rect 277228 698260 277229 698324
rect 277163 698259 277229 698260
rect 277531 698324 277597 698325
rect 277531 698260 277532 698324
rect 277596 698260 277597 698324
rect 277531 698259 277597 698260
rect 277166 698050 277226 698259
rect 277534 698050 277594 698259
rect 277718 698053 277778 698531
rect 284894 698325 284954 698531
rect 288022 698325 288082 698531
rect 284891 698324 284957 698325
rect 284891 698260 284892 698324
rect 284956 698260 284957 698324
rect 286731 698324 286797 698325
rect 286731 698310 286732 698324
rect 284891 698259 284957 698260
rect 286550 698260 286732 698310
rect 286796 698260 286797 698324
rect 286550 698259 286797 698260
rect 287835 698324 287901 698325
rect 287835 698260 287836 698324
rect 287900 698260 287901 698324
rect 287835 698259 287901 698260
rect 288019 698324 288085 698325
rect 288019 698260 288020 698324
rect 288084 698260 288085 698324
rect 288019 698259 288085 698260
rect 286550 698250 286794 698259
rect 286179 698188 286245 698189
rect 286179 698124 286180 698188
rect 286244 698124 286245 698188
rect 286179 698123 286245 698124
rect 277166 697990 277594 698050
rect 277715 698052 277781 698053
rect 277715 697988 277716 698052
rect 277780 697988 277781 698052
rect 277715 697987 277781 697988
rect 267779 697916 267845 697917
rect 267779 697852 267780 697916
rect 267844 697852 267845 697916
rect 267779 697851 267845 697852
rect 268147 697916 268213 697917
rect 268147 697852 268148 697916
rect 268212 697852 268213 697916
rect 268147 697851 268213 697852
rect 276979 697916 277045 697917
rect 276979 697852 276980 697916
rect 277044 697852 277045 697916
rect 286182 697914 286242 698123
rect 286363 698052 286429 698053
rect 286363 697988 286364 698052
rect 286428 698050 286429 698052
rect 286550 698050 286610 698250
rect 286731 698188 286797 698189
rect 286731 698124 286732 698188
rect 286796 698124 286797 698188
rect 286731 698123 286797 698124
rect 286428 697990 286610 698050
rect 286428 697988 286429 697990
rect 286363 697987 286429 697988
rect 286734 697914 286794 698123
rect 287838 697917 287898 698259
rect 296302 697917 296362 698531
rect 296483 698324 296549 698325
rect 296483 698260 296484 698324
rect 296548 698260 296549 698324
rect 296483 698259 296549 698260
rect 296851 698324 296917 698325
rect 296851 698260 296852 698324
rect 296916 698260 296917 698324
rect 296851 698259 296917 698260
rect 296486 698050 296546 698259
rect 296854 698050 296914 698259
rect 297038 698053 297098 698531
rect 304214 698325 304274 698531
rect 307342 698325 307402 698531
rect 304211 698324 304277 698325
rect 304211 698260 304212 698324
rect 304276 698260 304277 698324
rect 306051 698324 306117 698325
rect 306051 698310 306052 698324
rect 304211 698259 304277 698260
rect 305870 698260 306052 698310
rect 306116 698260 306117 698324
rect 305870 698259 306117 698260
rect 307155 698324 307221 698325
rect 307155 698260 307156 698324
rect 307220 698260 307221 698324
rect 307155 698259 307221 698260
rect 307339 698324 307405 698325
rect 307339 698260 307340 698324
rect 307404 698260 307405 698324
rect 307339 698259 307405 698260
rect 305870 698250 306114 698259
rect 305499 698188 305565 698189
rect 305499 698124 305500 698188
rect 305564 698124 305565 698188
rect 305499 698123 305565 698124
rect 296486 697990 296914 698050
rect 297035 698052 297101 698053
rect 297035 697988 297036 698052
rect 297100 697988 297101 698052
rect 297035 697987 297101 697988
rect 286182 697854 286794 697914
rect 287835 697916 287901 697917
rect 276979 697851 277045 697852
rect 287835 697852 287836 697916
rect 287900 697852 287901 697916
rect 287835 697851 287901 697852
rect 296299 697916 296365 697917
rect 296299 697852 296300 697916
rect 296364 697852 296365 697916
rect 305502 697914 305562 698123
rect 305683 698052 305749 698053
rect 305683 697988 305684 698052
rect 305748 698050 305749 698052
rect 305870 698050 305930 698250
rect 306051 698188 306117 698189
rect 306051 698124 306052 698188
rect 306116 698124 306117 698188
rect 306051 698123 306117 698124
rect 305748 697990 305930 698050
rect 305748 697988 305749 697990
rect 305683 697987 305749 697988
rect 306054 697914 306114 698123
rect 307158 697917 307218 698259
rect 315622 697917 315682 698531
rect 315803 698324 315869 698325
rect 315803 698260 315804 698324
rect 315868 698260 315869 698324
rect 315803 698259 315869 698260
rect 316171 698324 316237 698325
rect 316171 698260 316172 698324
rect 316236 698260 316237 698324
rect 316171 698259 316237 698260
rect 315806 698050 315866 698259
rect 316174 698050 316234 698259
rect 316358 698053 316418 698531
rect 323534 698325 323594 698531
rect 326662 698325 326722 698531
rect 323531 698324 323597 698325
rect 323531 698260 323532 698324
rect 323596 698260 323597 698324
rect 325371 698324 325437 698325
rect 325371 698310 325372 698324
rect 323531 698259 323597 698260
rect 325190 698260 325372 698310
rect 325436 698260 325437 698324
rect 325190 698259 325437 698260
rect 326475 698324 326541 698325
rect 326475 698260 326476 698324
rect 326540 698260 326541 698324
rect 326475 698259 326541 698260
rect 326659 698324 326725 698325
rect 326659 698260 326660 698324
rect 326724 698260 326725 698324
rect 326659 698259 326725 698260
rect 325190 698250 325434 698259
rect 324819 698188 324885 698189
rect 324819 698124 324820 698188
rect 324884 698124 324885 698188
rect 324819 698123 324885 698124
rect 315806 697990 316234 698050
rect 316355 698052 316421 698053
rect 316355 697988 316356 698052
rect 316420 697988 316421 698052
rect 316355 697987 316421 697988
rect 305502 697854 306114 697914
rect 307155 697916 307221 697917
rect 296299 697851 296365 697852
rect 307155 697852 307156 697916
rect 307220 697852 307221 697916
rect 307155 697851 307221 697852
rect 315619 697916 315685 697917
rect 315619 697852 315620 697916
rect 315684 697852 315685 697916
rect 324822 697914 324882 698123
rect 325003 698052 325069 698053
rect 325003 697988 325004 698052
rect 325068 698050 325069 698052
rect 325190 698050 325250 698250
rect 325371 698188 325437 698189
rect 325371 698124 325372 698188
rect 325436 698124 325437 698188
rect 325371 698123 325437 698124
rect 325068 697990 325250 698050
rect 325068 697988 325069 697990
rect 325003 697987 325069 697988
rect 325374 697914 325434 698123
rect 326478 697917 326538 698259
rect 334942 697917 335002 698531
rect 335123 698324 335189 698325
rect 335123 698260 335124 698324
rect 335188 698260 335189 698324
rect 335123 698259 335189 698260
rect 335491 698324 335557 698325
rect 335491 698260 335492 698324
rect 335556 698260 335557 698324
rect 335491 698259 335557 698260
rect 335126 698050 335186 698259
rect 335494 698050 335554 698259
rect 335678 698053 335738 698531
rect 342854 698325 342914 698531
rect 345982 698325 346042 698531
rect 342851 698324 342917 698325
rect 342851 698260 342852 698324
rect 342916 698260 342917 698324
rect 344691 698324 344757 698325
rect 344691 698310 344692 698324
rect 342851 698259 342917 698260
rect 344510 698260 344692 698310
rect 344756 698260 344757 698324
rect 344510 698259 344757 698260
rect 345795 698324 345861 698325
rect 345795 698260 345796 698324
rect 345860 698260 345861 698324
rect 345795 698259 345861 698260
rect 345979 698324 346045 698325
rect 345979 698260 345980 698324
rect 346044 698260 346045 698324
rect 345979 698259 346045 698260
rect 344510 698250 344754 698259
rect 344139 698188 344205 698189
rect 344139 698124 344140 698188
rect 344204 698124 344205 698188
rect 344139 698123 344205 698124
rect 335126 697990 335554 698050
rect 335675 698052 335741 698053
rect 335675 697988 335676 698052
rect 335740 697988 335741 698052
rect 335675 697987 335741 697988
rect 324822 697854 325434 697914
rect 326475 697916 326541 697917
rect 315619 697851 315685 697852
rect 326475 697852 326476 697916
rect 326540 697852 326541 697916
rect 326475 697851 326541 697852
rect 334939 697916 335005 697917
rect 334939 697852 334940 697916
rect 335004 697852 335005 697916
rect 344142 697914 344202 698123
rect 344323 698052 344389 698053
rect 344323 697988 344324 698052
rect 344388 698050 344389 698052
rect 344510 698050 344570 698250
rect 344691 698188 344757 698189
rect 344691 698124 344692 698188
rect 344756 698124 344757 698188
rect 344691 698123 344757 698124
rect 344388 697990 344570 698050
rect 344388 697988 344389 697990
rect 344323 697987 344389 697988
rect 344694 697914 344754 698123
rect 345798 697917 345858 698259
rect 354262 697917 354322 698531
rect 354443 698324 354509 698325
rect 354443 698260 354444 698324
rect 354508 698260 354509 698324
rect 354443 698259 354509 698260
rect 354811 698324 354877 698325
rect 354811 698260 354812 698324
rect 354876 698260 354877 698324
rect 354811 698259 354877 698260
rect 354446 698050 354506 698259
rect 354814 698050 354874 698259
rect 354998 698053 355058 698531
rect 362174 698325 362234 698531
rect 365302 698325 365362 698531
rect 362171 698324 362237 698325
rect 362171 698260 362172 698324
rect 362236 698260 362237 698324
rect 364011 698324 364077 698325
rect 364011 698310 364012 698324
rect 362171 698259 362237 698260
rect 363830 698260 364012 698310
rect 364076 698260 364077 698324
rect 363830 698259 364077 698260
rect 365115 698324 365181 698325
rect 365115 698260 365116 698324
rect 365180 698260 365181 698324
rect 365115 698259 365181 698260
rect 365299 698324 365365 698325
rect 365299 698260 365300 698324
rect 365364 698260 365365 698324
rect 365299 698259 365365 698260
rect 363830 698250 364074 698259
rect 363459 698188 363525 698189
rect 363459 698124 363460 698188
rect 363524 698124 363525 698188
rect 363459 698123 363525 698124
rect 354446 697990 354874 698050
rect 354995 698052 355061 698053
rect 354995 697988 354996 698052
rect 355060 697988 355061 698052
rect 354995 697987 355061 697988
rect 344142 697854 344754 697914
rect 345795 697916 345861 697917
rect 334939 697851 335005 697852
rect 345795 697852 345796 697916
rect 345860 697852 345861 697916
rect 345795 697851 345861 697852
rect 354259 697916 354325 697917
rect 354259 697852 354260 697916
rect 354324 697852 354325 697916
rect 363462 697914 363522 698123
rect 363643 698052 363709 698053
rect 363643 697988 363644 698052
rect 363708 698050 363709 698052
rect 363830 698050 363890 698250
rect 364011 698188 364077 698189
rect 364011 698124 364012 698188
rect 364076 698124 364077 698188
rect 364011 698123 364077 698124
rect 363708 697990 363890 698050
rect 363708 697988 363709 697990
rect 363643 697987 363709 697988
rect 364014 697914 364074 698123
rect 365118 697917 365178 698259
rect 373582 697917 373642 698531
rect 373763 698324 373829 698325
rect 373763 698260 373764 698324
rect 373828 698260 373829 698324
rect 373763 698259 373829 698260
rect 374131 698324 374197 698325
rect 374131 698260 374132 698324
rect 374196 698260 374197 698324
rect 374131 698259 374197 698260
rect 373766 698050 373826 698259
rect 374134 698050 374194 698259
rect 374318 698053 374378 698531
rect 382966 698053 383026 698531
rect 383518 698325 383578 698667
rect 389406 698597 389466 699075
rect 389403 698596 389469 698597
rect 389403 698532 389404 698596
rect 389468 698532 389469 698596
rect 389403 698531 389469 698532
rect 383147 698324 383213 698325
rect 383147 698260 383148 698324
rect 383212 698260 383213 698324
rect 383147 698259 383213 698260
rect 383515 698324 383581 698325
rect 383515 698260 383516 698324
rect 383580 698260 383581 698324
rect 383515 698259 383581 698260
rect 373766 697990 374194 698050
rect 374315 698052 374381 698053
rect 374315 697988 374316 698052
rect 374380 697988 374381 698052
rect 374315 697987 374381 697988
rect 382963 698052 383029 698053
rect 382963 697988 382964 698052
rect 383028 697988 383029 698052
rect 382963 697987 383029 697988
rect 363462 697854 364074 697914
rect 365115 697916 365181 697917
rect 354259 697851 354325 697852
rect 365115 697852 365116 697916
rect 365180 697852 365181 697916
rect 365115 697851 365181 697852
rect 373579 697916 373645 697917
rect 373579 697852 373580 697916
rect 373644 697852 373645 697916
rect 383150 697914 383210 698259
rect 430622 698189 430682 699075
rect 430619 698188 430685 698189
rect 430619 698124 430620 698188
rect 430684 698124 430685 698188
rect 430619 698123 430685 698124
rect 450678 697917 450738 699075
rect 383515 697916 383581 697917
rect 383515 697914 383516 697916
rect 383150 697854 383516 697914
rect 373579 697851 373645 697852
rect 383515 697852 383516 697854
rect 383580 697852 383581 697916
rect 383515 697851 383581 697852
rect 450675 697916 450741 697917
rect 450675 697852 450676 697916
rect 450740 697852 450741 697916
rect 450675 697851 450741 697852
rect 460982 697781 461042 699075
rect 460979 697780 461045 697781
rect 460979 697716 460980 697780
rect 461044 697716 461045 697780
rect 460979 697715 461045 697716
rect 476070 697509 476130 699075
rect 539918 698461 539978 699075
rect 539915 698460 539981 698461
rect 539915 698396 539916 698460
rect 539980 698396 539981 698460
rect 539915 698395 539981 698396
rect 476067 697508 476133 697509
rect 476067 697444 476068 697508
rect 476132 697444 476133 697508
rect 476067 697443 476133 697444
rect 258027 697100 258093 697101
rect 258027 697036 258028 697100
rect 258092 697036 258093 697100
rect 258027 697035 258093 697036
rect 258579 697100 258645 697101
rect 258579 697036 258580 697100
rect 258644 697036 258645 697100
rect 258579 697035 258645 697036
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect 8608 687454 8928 687486
rect 8608 687218 8650 687454
rect 8886 687218 8928 687454
rect 8608 687134 8928 687218
rect 8608 686898 8650 687134
rect 8886 686898 8928 687134
rect 8608 686866 8928 686898
rect 39328 687454 39648 687486
rect 39328 687218 39370 687454
rect 39606 687218 39648 687454
rect 39328 687134 39648 687218
rect 39328 686898 39370 687134
rect 39606 686898 39648 687134
rect 39328 686866 39648 686898
rect 70048 687454 70368 687486
rect 70048 687218 70090 687454
rect 70326 687218 70368 687454
rect 70048 687134 70368 687218
rect 70048 686898 70090 687134
rect 70326 686898 70368 687134
rect 70048 686866 70368 686898
rect 100768 687454 101088 687486
rect 100768 687218 100810 687454
rect 101046 687218 101088 687454
rect 100768 687134 101088 687218
rect 100768 686898 100810 687134
rect 101046 686898 101088 687134
rect 100768 686866 101088 686898
rect 131488 687454 131808 687486
rect 131488 687218 131530 687454
rect 131766 687218 131808 687454
rect 131488 687134 131808 687218
rect 131488 686898 131530 687134
rect 131766 686898 131808 687134
rect 131488 686866 131808 686898
rect 162208 687454 162528 687486
rect 162208 687218 162250 687454
rect 162486 687218 162528 687454
rect 162208 687134 162528 687218
rect 162208 686898 162250 687134
rect 162486 686898 162528 687134
rect 162208 686866 162528 686898
rect 192928 687454 193248 687486
rect 192928 687218 192970 687454
rect 193206 687218 193248 687454
rect 192928 687134 193248 687218
rect 192928 686898 192970 687134
rect 193206 686898 193248 687134
rect 192928 686866 193248 686898
rect 223648 687454 223968 687486
rect 223648 687218 223690 687454
rect 223926 687218 223968 687454
rect 223648 687134 223968 687218
rect 223648 686898 223690 687134
rect 223926 686898 223968 687134
rect 223648 686866 223968 686898
rect 254368 687454 254688 687486
rect 254368 687218 254410 687454
rect 254646 687218 254688 687454
rect 254368 687134 254688 687218
rect 254368 686898 254410 687134
rect 254646 686898 254688 687134
rect 254368 686866 254688 686898
rect 285088 687454 285408 687486
rect 285088 687218 285130 687454
rect 285366 687218 285408 687454
rect 285088 687134 285408 687218
rect 285088 686898 285130 687134
rect 285366 686898 285408 687134
rect 285088 686866 285408 686898
rect 315808 687454 316128 687486
rect 315808 687218 315850 687454
rect 316086 687218 316128 687454
rect 315808 687134 316128 687218
rect 315808 686898 315850 687134
rect 316086 686898 316128 687134
rect 315808 686866 316128 686898
rect 346528 687454 346848 687486
rect 346528 687218 346570 687454
rect 346806 687218 346848 687454
rect 346528 687134 346848 687218
rect 346528 686898 346570 687134
rect 346806 686898 346848 687134
rect 346528 686866 346848 686898
rect 377248 687454 377568 687486
rect 377248 687218 377290 687454
rect 377526 687218 377568 687454
rect 377248 687134 377568 687218
rect 377248 686898 377290 687134
rect 377526 686898 377568 687134
rect 377248 686866 377568 686898
rect 407968 687454 408288 687486
rect 407968 687218 408010 687454
rect 408246 687218 408288 687454
rect 407968 687134 408288 687218
rect 407968 686898 408010 687134
rect 408246 686898 408288 687134
rect 407968 686866 408288 686898
rect 438688 687454 439008 687486
rect 438688 687218 438730 687454
rect 438966 687218 439008 687454
rect 438688 687134 439008 687218
rect 438688 686898 438730 687134
rect 438966 686898 439008 687134
rect 438688 686866 439008 686898
rect 469408 687454 469728 687486
rect 469408 687218 469450 687454
rect 469686 687218 469728 687454
rect 469408 687134 469728 687218
rect 469408 686898 469450 687134
rect 469686 686898 469728 687134
rect 469408 686866 469728 686898
rect 500128 687454 500448 687486
rect 500128 687218 500170 687454
rect 500406 687218 500448 687454
rect 500128 687134 500448 687218
rect 500128 686898 500170 687134
rect 500406 686898 500448 687134
rect 500128 686866 500448 686898
rect 530848 687454 531168 687486
rect 530848 687218 530890 687454
rect 531126 687218 531168 687454
rect 530848 687134 531168 687218
rect 530848 686898 530890 687134
rect 531126 686898 531168 687134
rect 530848 686866 531168 686898
rect 561568 687454 561888 687486
rect 561568 687218 561610 687454
rect 561846 687218 561888 687454
rect 561568 687134 561888 687218
rect 561568 686898 561610 687134
rect 561846 686898 561888 687134
rect 561568 686866 561888 686898
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 23968 669454 24288 669486
rect 23968 669218 24010 669454
rect 24246 669218 24288 669454
rect 23968 669134 24288 669218
rect 23968 668898 24010 669134
rect 24246 668898 24288 669134
rect 23968 668866 24288 668898
rect 54688 669454 55008 669486
rect 54688 669218 54730 669454
rect 54966 669218 55008 669454
rect 54688 669134 55008 669218
rect 54688 668898 54730 669134
rect 54966 668898 55008 669134
rect 54688 668866 55008 668898
rect 85408 669454 85728 669486
rect 85408 669218 85450 669454
rect 85686 669218 85728 669454
rect 85408 669134 85728 669218
rect 85408 668898 85450 669134
rect 85686 668898 85728 669134
rect 85408 668866 85728 668898
rect 116128 669454 116448 669486
rect 116128 669218 116170 669454
rect 116406 669218 116448 669454
rect 116128 669134 116448 669218
rect 116128 668898 116170 669134
rect 116406 668898 116448 669134
rect 116128 668866 116448 668898
rect 146848 669454 147168 669486
rect 146848 669218 146890 669454
rect 147126 669218 147168 669454
rect 146848 669134 147168 669218
rect 146848 668898 146890 669134
rect 147126 668898 147168 669134
rect 146848 668866 147168 668898
rect 177568 669454 177888 669486
rect 177568 669218 177610 669454
rect 177846 669218 177888 669454
rect 177568 669134 177888 669218
rect 177568 668898 177610 669134
rect 177846 668898 177888 669134
rect 177568 668866 177888 668898
rect 208288 669454 208608 669486
rect 208288 669218 208330 669454
rect 208566 669218 208608 669454
rect 208288 669134 208608 669218
rect 208288 668898 208330 669134
rect 208566 668898 208608 669134
rect 208288 668866 208608 668898
rect 239008 669454 239328 669486
rect 239008 669218 239050 669454
rect 239286 669218 239328 669454
rect 239008 669134 239328 669218
rect 239008 668898 239050 669134
rect 239286 668898 239328 669134
rect 239008 668866 239328 668898
rect 269728 669454 270048 669486
rect 269728 669218 269770 669454
rect 270006 669218 270048 669454
rect 269728 669134 270048 669218
rect 269728 668898 269770 669134
rect 270006 668898 270048 669134
rect 269728 668866 270048 668898
rect 300448 669454 300768 669486
rect 300448 669218 300490 669454
rect 300726 669218 300768 669454
rect 300448 669134 300768 669218
rect 300448 668898 300490 669134
rect 300726 668898 300768 669134
rect 300448 668866 300768 668898
rect 331168 669454 331488 669486
rect 331168 669218 331210 669454
rect 331446 669218 331488 669454
rect 331168 669134 331488 669218
rect 331168 668898 331210 669134
rect 331446 668898 331488 669134
rect 331168 668866 331488 668898
rect 361888 669454 362208 669486
rect 361888 669218 361930 669454
rect 362166 669218 362208 669454
rect 361888 669134 362208 669218
rect 361888 668898 361930 669134
rect 362166 668898 362208 669134
rect 361888 668866 362208 668898
rect 392608 669454 392928 669486
rect 392608 669218 392650 669454
rect 392886 669218 392928 669454
rect 392608 669134 392928 669218
rect 392608 668898 392650 669134
rect 392886 668898 392928 669134
rect 392608 668866 392928 668898
rect 423328 669454 423648 669486
rect 423328 669218 423370 669454
rect 423606 669218 423648 669454
rect 423328 669134 423648 669218
rect 423328 668898 423370 669134
rect 423606 668898 423648 669134
rect 423328 668866 423648 668898
rect 454048 669454 454368 669486
rect 454048 669218 454090 669454
rect 454326 669218 454368 669454
rect 454048 669134 454368 669218
rect 454048 668898 454090 669134
rect 454326 668898 454368 669134
rect 454048 668866 454368 668898
rect 484768 669454 485088 669486
rect 484768 669218 484810 669454
rect 485046 669218 485088 669454
rect 484768 669134 485088 669218
rect 484768 668898 484810 669134
rect 485046 668898 485088 669134
rect 484768 668866 485088 668898
rect 515488 669454 515808 669486
rect 515488 669218 515530 669454
rect 515766 669218 515808 669454
rect 515488 669134 515808 669218
rect 515488 668898 515530 669134
rect 515766 668898 515808 669134
rect 515488 668866 515808 668898
rect 546208 669454 546528 669486
rect 546208 669218 546250 669454
rect 546486 669218 546528 669454
rect 546208 669134 546528 669218
rect 546208 668898 546250 669134
rect 546486 668898 546528 669134
rect 546208 668866 546528 668898
rect 576928 669454 577248 669486
rect 576928 669218 576970 669454
rect 577206 669218 577248 669454
rect 576928 669134 577248 669218
rect 576928 668898 576970 669134
rect 577206 668898 577248 669134
rect 576928 668866 577248 668898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect 8608 651454 8928 651486
rect 8608 651218 8650 651454
rect 8886 651218 8928 651454
rect 8608 651134 8928 651218
rect 8608 650898 8650 651134
rect 8886 650898 8928 651134
rect 8608 650866 8928 650898
rect 39328 651454 39648 651486
rect 39328 651218 39370 651454
rect 39606 651218 39648 651454
rect 39328 651134 39648 651218
rect 39328 650898 39370 651134
rect 39606 650898 39648 651134
rect 39328 650866 39648 650898
rect 70048 651454 70368 651486
rect 70048 651218 70090 651454
rect 70326 651218 70368 651454
rect 70048 651134 70368 651218
rect 70048 650898 70090 651134
rect 70326 650898 70368 651134
rect 70048 650866 70368 650898
rect 100768 651454 101088 651486
rect 100768 651218 100810 651454
rect 101046 651218 101088 651454
rect 100768 651134 101088 651218
rect 100768 650898 100810 651134
rect 101046 650898 101088 651134
rect 100768 650866 101088 650898
rect 131488 651454 131808 651486
rect 131488 651218 131530 651454
rect 131766 651218 131808 651454
rect 131488 651134 131808 651218
rect 131488 650898 131530 651134
rect 131766 650898 131808 651134
rect 131488 650866 131808 650898
rect 162208 651454 162528 651486
rect 162208 651218 162250 651454
rect 162486 651218 162528 651454
rect 162208 651134 162528 651218
rect 162208 650898 162250 651134
rect 162486 650898 162528 651134
rect 162208 650866 162528 650898
rect 192928 651454 193248 651486
rect 192928 651218 192970 651454
rect 193206 651218 193248 651454
rect 192928 651134 193248 651218
rect 192928 650898 192970 651134
rect 193206 650898 193248 651134
rect 192928 650866 193248 650898
rect 223648 651454 223968 651486
rect 223648 651218 223690 651454
rect 223926 651218 223968 651454
rect 223648 651134 223968 651218
rect 223648 650898 223690 651134
rect 223926 650898 223968 651134
rect 223648 650866 223968 650898
rect 254368 651454 254688 651486
rect 254368 651218 254410 651454
rect 254646 651218 254688 651454
rect 254368 651134 254688 651218
rect 254368 650898 254410 651134
rect 254646 650898 254688 651134
rect 254368 650866 254688 650898
rect 285088 651454 285408 651486
rect 285088 651218 285130 651454
rect 285366 651218 285408 651454
rect 285088 651134 285408 651218
rect 285088 650898 285130 651134
rect 285366 650898 285408 651134
rect 285088 650866 285408 650898
rect 315808 651454 316128 651486
rect 315808 651218 315850 651454
rect 316086 651218 316128 651454
rect 315808 651134 316128 651218
rect 315808 650898 315850 651134
rect 316086 650898 316128 651134
rect 315808 650866 316128 650898
rect 346528 651454 346848 651486
rect 346528 651218 346570 651454
rect 346806 651218 346848 651454
rect 346528 651134 346848 651218
rect 346528 650898 346570 651134
rect 346806 650898 346848 651134
rect 346528 650866 346848 650898
rect 377248 651454 377568 651486
rect 377248 651218 377290 651454
rect 377526 651218 377568 651454
rect 377248 651134 377568 651218
rect 377248 650898 377290 651134
rect 377526 650898 377568 651134
rect 377248 650866 377568 650898
rect 407968 651454 408288 651486
rect 407968 651218 408010 651454
rect 408246 651218 408288 651454
rect 407968 651134 408288 651218
rect 407968 650898 408010 651134
rect 408246 650898 408288 651134
rect 407968 650866 408288 650898
rect 438688 651454 439008 651486
rect 438688 651218 438730 651454
rect 438966 651218 439008 651454
rect 438688 651134 439008 651218
rect 438688 650898 438730 651134
rect 438966 650898 439008 651134
rect 438688 650866 439008 650898
rect 469408 651454 469728 651486
rect 469408 651218 469450 651454
rect 469686 651218 469728 651454
rect 469408 651134 469728 651218
rect 469408 650898 469450 651134
rect 469686 650898 469728 651134
rect 469408 650866 469728 650898
rect 500128 651454 500448 651486
rect 500128 651218 500170 651454
rect 500406 651218 500448 651454
rect 500128 651134 500448 651218
rect 500128 650898 500170 651134
rect 500406 650898 500448 651134
rect 500128 650866 500448 650898
rect 530848 651454 531168 651486
rect 530848 651218 530890 651454
rect 531126 651218 531168 651454
rect 530848 651134 531168 651218
rect 530848 650898 530890 651134
rect 531126 650898 531168 651134
rect 530848 650866 531168 650898
rect 561568 651454 561888 651486
rect 561568 651218 561610 651454
rect 561846 651218 561888 651454
rect 561568 651134 561888 651218
rect 561568 650898 561610 651134
rect 561846 650898 561888 651134
rect 561568 650866 561888 650898
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 23968 633454 24288 633486
rect 23968 633218 24010 633454
rect 24246 633218 24288 633454
rect 23968 633134 24288 633218
rect 23968 632898 24010 633134
rect 24246 632898 24288 633134
rect 23968 632866 24288 632898
rect 54688 633454 55008 633486
rect 54688 633218 54730 633454
rect 54966 633218 55008 633454
rect 54688 633134 55008 633218
rect 54688 632898 54730 633134
rect 54966 632898 55008 633134
rect 54688 632866 55008 632898
rect 85408 633454 85728 633486
rect 85408 633218 85450 633454
rect 85686 633218 85728 633454
rect 85408 633134 85728 633218
rect 85408 632898 85450 633134
rect 85686 632898 85728 633134
rect 85408 632866 85728 632898
rect 116128 633454 116448 633486
rect 116128 633218 116170 633454
rect 116406 633218 116448 633454
rect 116128 633134 116448 633218
rect 116128 632898 116170 633134
rect 116406 632898 116448 633134
rect 116128 632866 116448 632898
rect 146848 633454 147168 633486
rect 146848 633218 146890 633454
rect 147126 633218 147168 633454
rect 146848 633134 147168 633218
rect 146848 632898 146890 633134
rect 147126 632898 147168 633134
rect 146848 632866 147168 632898
rect 177568 633454 177888 633486
rect 177568 633218 177610 633454
rect 177846 633218 177888 633454
rect 177568 633134 177888 633218
rect 177568 632898 177610 633134
rect 177846 632898 177888 633134
rect 177568 632866 177888 632898
rect 208288 633454 208608 633486
rect 208288 633218 208330 633454
rect 208566 633218 208608 633454
rect 208288 633134 208608 633218
rect 208288 632898 208330 633134
rect 208566 632898 208608 633134
rect 208288 632866 208608 632898
rect 239008 633454 239328 633486
rect 239008 633218 239050 633454
rect 239286 633218 239328 633454
rect 239008 633134 239328 633218
rect 239008 632898 239050 633134
rect 239286 632898 239328 633134
rect 239008 632866 239328 632898
rect 269728 633454 270048 633486
rect 269728 633218 269770 633454
rect 270006 633218 270048 633454
rect 269728 633134 270048 633218
rect 269728 632898 269770 633134
rect 270006 632898 270048 633134
rect 269728 632866 270048 632898
rect 300448 633454 300768 633486
rect 300448 633218 300490 633454
rect 300726 633218 300768 633454
rect 300448 633134 300768 633218
rect 300448 632898 300490 633134
rect 300726 632898 300768 633134
rect 300448 632866 300768 632898
rect 331168 633454 331488 633486
rect 331168 633218 331210 633454
rect 331446 633218 331488 633454
rect 331168 633134 331488 633218
rect 331168 632898 331210 633134
rect 331446 632898 331488 633134
rect 331168 632866 331488 632898
rect 361888 633454 362208 633486
rect 361888 633218 361930 633454
rect 362166 633218 362208 633454
rect 361888 633134 362208 633218
rect 361888 632898 361930 633134
rect 362166 632898 362208 633134
rect 361888 632866 362208 632898
rect 392608 633454 392928 633486
rect 392608 633218 392650 633454
rect 392886 633218 392928 633454
rect 392608 633134 392928 633218
rect 392608 632898 392650 633134
rect 392886 632898 392928 633134
rect 392608 632866 392928 632898
rect 423328 633454 423648 633486
rect 423328 633218 423370 633454
rect 423606 633218 423648 633454
rect 423328 633134 423648 633218
rect 423328 632898 423370 633134
rect 423606 632898 423648 633134
rect 423328 632866 423648 632898
rect 454048 633454 454368 633486
rect 454048 633218 454090 633454
rect 454326 633218 454368 633454
rect 454048 633134 454368 633218
rect 454048 632898 454090 633134
rect 454326 632898 454368 633134
rect 454048 632866 454368 632898
rect 484768 633454 485088 633486
rect 484768 633218 484810 633454
rect 485046 633218 485088 633454
rect 484768 633134 485088 633218
rect 484768 632898 484810 633134
rect 485046 632898 485088 633134
rect 484768 632866 485088 632898
rect 515488 633454 515808 633486
rect 515488 633218 515530 633454
rect 515766 633218 515808 633454
rect 515488 633134 515808 633218
rect 515488 632898 515530 633134
rect 515766 632898 515808 633134
rect 515488 632866 515808 632898
rect 546208 633454 546528 633486
rect 546208 633218 546250 633454
rect 546486 633218 546528 633454
rect 546208 633134 546528 633218
rect 546208 632898 546250 633134
rect 546486 632898 546528 633134
rect 546208 632866 546528 632898
rect 576928 633454 577248 633486
rect 576928 633218 576970 633454
rect 577206 633218 577248 633454
rect 576928 633134 577248 633218
rect 576928 632898 576970 633134
rect 577206 632898 577248 633134
rect 576928 632866 577248 632898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect 8608 615454 8928 615486
rect 8608 615218 8650 615454
rect 8886 615218 8928 615454
rect 8608 615134 8928 615218
rect 8608 614898 8650 615134
rect 8886 614898 8928 615134
rect 8608 614866 8928 614898
rect 39328 615454 39648 615486
rect 39328 615218 39370 615454
rect 39606 615218 39648 615454
rect 39328 615134 39648 615218
rect 39328 614898 39370 615134
rect 39606 614898 39648 615134
rect 39328 614866 39648 614898
rect 70048 615454 70368 615486
rect 70048 615218 70090 615454
rect 70326 615218 70368 615454
rect 70048 615134 70368 615218
rect 70048 614898 70090 615134
rect 70326 614898 70368 615134
rect 70048 614866 70368 614898
rect 100768 615454 101088 615486
rect 100768 615218 100810 615454
rect 101046 615218 101088 615454
rect 100768 615134 101088 615218
rect 100768 614898 100810 615134
rect 101046 614898 101088 615134
rect 100768 614866 101088 614898
rect 131488 615454 131808 615486
rect 131488 615218 131530 615454
rect 131766 615218 131808 615454
rect 131488 615134 131808 615218
rect 131488 614898 131530 615134
rect 131766 614898 131808 615134
rect 131488 614866 131808 614898
rect 162208 615454 162528 615486
rect 162208 615218 162250 615454
rect 162486 615218 162528 615454
rect 162208 615134 162528 615218
rect 162208 614898 162250 615134
rect 162486 614898 162528 615134
rect 162208 614866 162528 614898
rect 192928 615454 193248 615486
rect 192928 615218 192970 615454
rect 193206 615218 193248 615454
rect 192928 615134 193248 615218
rect 192928 614898 192970 615134
rect 193206 614898 193248 615134
rect 192928 614866 193248 614898
rect 223648 615454 223968 615486
rect 223648 615218 223690 615454
rect 223926 615218 223968 615454
rect 223648 615134 223968 615218
rect 223648 614898 223690 615134
rect 223926 614898 223968 615134
rect 223648 614866 223968 614898
rect 254368 615454 254688 615486
rect 254368 615218 254410 615454
rect 254646 615218 254688 615454
rect 254368 615134 254688 615218
rect 254368 614898 254410 615134
rect 254646 614898 254688 615134
rect 254368 614866 254688 614898
rect 285088 615454 285408 615486
rect 285088 615218 285130 615454
rect 285366 615218 285408 615454
rect 285088 615134 285408 615218
rect 285088 614898 285130 615134
rect 285366 614898 285408 615134
rect 285088 614866 285408 614898
rect 315808 615454 316128 615486
rect 315808 615218 315850 615454
rect 316086 615218 316128 615454
rect 315808 615134 316128 615218
rect 315808 614898 315850 615134
rect 316086 614898 316128 615134
rect 315808 614866 316128 614898
rect 346528 615454 346848 615486
rect 346528 615218 346570 615454
rect 346806 615218 346848 615454
rect 346528 615134 346848 615218
rect 346528 614898 346570 615134
rect 346806 614898 346848 615134
rect 346528 614866 346848 614898
rect 377248 615454 377568 615486
rect 377248 615218 377290 615454
rect 377526 615218 377568 615454
rect 377248 615134 377568 615218
rect 377248 614898 377290 615134
rect 377526 614898 377568 615134
rect 377248 614866 377568 614898
rect 407968 615454 408288 615486
rect 407968 615218 408010 615454
rect 408246 615218 408288 615454
rect 407968 615134 408288 615218
rect 407968 614898 408010 615134
rect 408246 614898 408288 615134
rect 407968 614866 408288 614898
rect 438688 615454 439008 615486
rect 438688 615218 438730 615454
rect 438966 615218 439008 615454
rect 438688 615134 439008 615218
rect 438688 614898 438730 615134
rect 438966 614898 439008 615134
rect 438688 614866 439008 614898
rect 469408 615454 469728 615486
rect 469408 615218 469450 615454
rect 469686 615218 469728 615454
rect 469408 615134 469728 615218
rect 469408 614898 469450 615134
rect 469686 614898 469728 615134
rect 469408 614866 469728 614898
rect 500128 615454 500448 615486
rect 500128 615218 500170 615454
rect 500406 615218 500448 615454
rect 500128 615134 500448 615218
rect 500128 614898 500170 615134
rect 500406 614898 500448 615134
rect 500128 614866 500448 614898
rect 530848 615454 531168 615486
rect 530848 615218 530890 615454
rect 531126 615218 531168 615454
rect 530848 615134 531168 615218
rect 530848 614898 530890 615134
rect 531126 614898 531168 615134
rect 530848 614866 531168 614898
rect 561568 615454 561888 615486
rect 561568 615218 561610 615454
rect 561846 615218 561888 615454
rect 561568 615134 561888 615218
rect 561568 614898 561610 615134
rect 561846 614898 561888 615134
rect 561568 614866 561888 614898
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 23968 597454 24288 597486
rect 23968 597218 24010 597454
rect 24246 597218 24288 597454
rect 23968 597134 24288 597218
rect 23968 596898 24010 597134
rect 24246 596898 24288 597134
rect 23968 596866 24288 596898
rect 54688 597454 55008 597486
rect 54688 597218 54730 597454
rect 54966 597218 55008 597454
rect 54688 597134 55008 597218
rect 54688 596898 54730 597134
rect 54966 596898 55008 597134
rect 54688 596866 55008 596898
rect 85408 597454 85728 597486
rect 85408 597218 85450 597454
rect 85686 597218 85728 597454
rect 85408 597134 85728 597218
rect 85408 596898 85450 597134
rect 85686 596898 85728 597134
rect 85408 596866 85728 596898
rect 116128 597454 116448 597486
rect 116128 597218 116170 597454
rect 116406 597218 116448 597454
rect 116128 597134 116448 597218
rect 116128 596898 116170 597134
rect 116406 596898 116448 597134
rect 116128 596866 116448 596898
rect 146848 597454 147168 597486
rect 146848 597218 146890 597454
rect 147126 597218 147168 597454
rect 146848 597134 147168 597218
rect 146848 596898 146890 597134
rect 147126 596898 147168 597134
rect 146848 596866 147168 596898
rect 177568 597454 177888 597486
rect 177568 597218 177610 597454
rect 177846 597218 177888 597454
rect 177568 597134 177888 597218
rect 177568 596898 177610 597134
rect 177846 596898 177888 597134
rect 177568 596866 177888 596898
rect 208288 597454 208608 597486
rect 208288 597218 208330 597454
rect 208566 597218 208608 597454
rect 208288 597134 208608 597218
rect 208288 596898 208330 597134
rect 208566 596898 208608 597134
rect 208288 596866 208608 596898
rect 239008 597454 239328 597486
rect 239008 597218 239050 597454
rect 239286 597218 239328 597454
rect 239008 597134 239328 597218
rect 239008 596898 239050 597134
rect 239286 596898 239328 597134
rect 239008 596866 239328 596898
rect 269728 597454 270048 597486
rect 269728 597218 269770 597454
rect 270006 597218 270048 597454
rect 269728 597134 270048 597218
rect 269728 596898 269770 597134
rect 270006 596898 270048 597134
rect 269728 596866 270048 596898
rect 300448 597454 300768 597486
rect 300448 597218 300490 597454
rect 300726 597218 300768 597454
rect 300448 597134 300768 597218
rect 300448 596898 300490 597134
rect 300726 596898 300768 597134
rect 300448 596866 300768 596898
rect 331168 597454 331488 597486
rect 331168 597218 331210 597454
rect 331446 597218 331488 597454
rect 331168 597134 331488 597218
rect 331168 596898 331210 597134
rect 331446 596898 331488 597134
rect 331168 596866 331488 596898
rect 361888 597454 362208 597486
rect 361888 597218 361930 597454
rect 362166 597218 362208 597454
rect 361888 597134 362208 597218
rect 361888 596898 361930 597134
rect 362166 596898 362208 597134
rect 361888 596866 362208 596898
rect 392608 597454 392928 597486
rect 392608 597218 392650 597454
rect 392886 597218 392928 597454
rect 392608 597134 392928 597218
rect 392608 596898 392650 597134
rect 392886 596898 392928 597134
rect 392608 596866 392928 596898
rect 423328 597454 423648 597486
rect 423328 597218 423370 597454
rect 423606 597218 423648 597454
rect 423328 597134 423648 597218
rect 423328 596898 423370 597134
rect 423606 596898 423648 597134
rect 423328 596866 423648 596898
rect 454048 597454 454368 597486
rect 454048 597218 454090 597454
rect 454326 597218 454368 597454
rect 454048 597134 454368 597218
rect 454048 596898 454090 597134
rect 454326 596898 454368 597134
rect 454048 596866 454368 596898
rect 484768 597454 485088 597486
rect 484768 597218 484810 597454
rect 485046 597218 485088 597454
rect 484768 597134 485088 597218
rect 484768 596898 484810 597134
rect 485046 596898 485088 597134
rect 484768 596866 485088 596898
rect 515488 597454 515808 597486
rect 515488 597218 515530 597454
rect 515766 597218 515808 597454
rect 515488 597134 515808 597218
rect 515488 596898 515530 597134
rect 515766 596898 515808 597134
rect 515488 596866 515808 596898
rect 546208 597454 546528 597486
rect 546208 597218 546250 597454
rect 546486 597218 546528 597454
rect 546208 597134 546528 597218
rect 546208 596898 546250 597134
rect 546486 596898 546528 597134
rect 546208 596866 546528 596898
rect 576928 597454 577248 597486
rect 576928 597218 576970 597454
rect 577206 597218 577248 597454
rect 576928 597134 577248 597218
rect 576928 596898 576970 597134
rect 577206 596898 577248 597134
rect 576928 596866 577248 596898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect 8608 579454 8928 579486
rect 8608 579218 8650 579454
rect 8886 579218 8928 579454
rect 8608 579134 8928 579218
rect 8608 578898 8650 579134
rect 8886 578898 8928 579134
rect 8608 578866 8928 578898
rect 39328 579454 39648 579486
rect 39328 579218 39370 579454
rect 39606 579218 39648 579454
rect 39328 579134 39648 579218
rect 39328 578898 39370 579134
rect 39606 578898 39648 579134
rect 39328 578866 39648 578898
rect 70048 579454 70368 579486
rect 70048 579218 70090 579454
rect 70326 579218 70368 579454
rect 70048 579134 70368 579218
rect 70048 578898 70090 579134
rect 70326 578898 70368 579134
rect 70048 578866 70368 578898
rect 100768 579454 101088 579486
rect 100768 579218 100810 579454
rect 101046 579218 101088 579454
rect 100768 579134 101088 579218
rect 100768 578898 100810 579134
rect 101046 578898 101088 579134
rect 100768 578866 101088 578898
rect 131488 579454 131808 579486
rect 131488 579218 131530 579454
rect 131766 579218 131808 579454
rect 131488 579134 131808 579218
rect 131488 578898 131530 579134
rect 131766 578898 131808 579134
rect 131488 578866 131808 578898
rect 162208 579454 162528 579486
rect 162208 579218 162250 579454
rect 162486 579218 162528 579454
rect 162208 579134 162528 579218
rect 162208 578898 162250 579134
rect 162486 578898 162528 579134
rect 162208 578866 162528 578898
rect 192928 579454 193248 579486
rect 192928 579218 192970 579454
rect 193206 579218 193248 579454
rect 192928 579134 193248 579218
rect 192928 578898 192970 579134
rect 193206 578898 193248 579134
rect 192928 578866 193248 578898
rect 223648 579454 223968 579486
rect 223648 579218 223690 579454
rect 223926 579218 223968 579454
rect 223648 579134 223968 579218
rect 223648 578898 223690 579134
rect 223926 578898 223968 579134
rect 223648 578866 223968 578898
rect 254368 579454 254688 579486
rect 254368 579218 254410 579454
rect 254646 579218 254688 579454
rect 254368 579134 254688 579218
rect 254368 578898 254410 579134
rect 254646 578898 254688 579134
rect 254368 578866 254688 578898
rect 285088 579454 285408 579486
rect 285088 579218 285130 579454
rect 285366 579218 285408 579454
rect 285088 579134 285408 579218
rect 285088 578898 285130 579134
rect 285366 578898 285408 579134
rect 285088 578866 285408 578898
rect 315808 579454 316128 579486
rect 315808 579218 315850 579454
rect 316086 579218 316128 579454
rect 315808 579134 316128 579218
rect 315808 578898 315850 579134
rect 316086 578898 316128 579134
rect 315808 578866 316128 578898
rect 346528 579454 346848 579486
rect 346528 579218 346570 579454
rect 346806 579218 346848 579454
rect 346528 579134 346848 579218
rect 346528 578898 346570 579134
rect 346806 578898 346848 579134
rect 346528 578866 346848 578898
rect 377248 579454 377568 579486
rect 377248 579218 377290 579454
rect 377526 579218 377568 579454
rect 377248 579134 377568 579218
rect 377248 578898 377290 579134
rect 377526 578898 377568 579134
rect 377248 578866 377568 578898
rect 407968 579454 408288 579486
rect 407968 579218 408010 579454
rect 408246 579218 408288 579454
rect 407968 579134 408288 579218
rect 407968 578898 408010 579134
rect 408246 578898 408288 579134
rect 407968 578866 408288 578898
rect 438688 579454 439008 579486
rect 438688 579218 438730 579454
rect 438966 579218 439008 579454
rect 438688 579134 439008 579218
rect 438688 578898 438730 579134
rect 438966 578898 439008 579134
rect 438688 578866 439008 578898
rect 469408 579454 469728 579486
rect 469408 579218 469450 579454
rect 469686 579218 469728 579454
rect 469408 579134 469728 579218
rect 469408 578898 469450 579134
rect 469686 578898 469728 579134
rect 469408 578866 469728 578898
rect 500128 579454 500448 579486
rect 500128 579218 500170 579454
rect 500406 579218 500448 579454
rect 500128 579134 500448 579218
rect 500128 578898 500170 579134
rect 500406 578898 500448 579134
rect 500128 578866 500448 578898
rect 530848 579454 531168 579486
rect 530848 579218 530890 579454
rect 531126 579218 531168 579454
rect 530848 579134 531168 579218
rect 530848 578898 530890 579134
rect 531126 578898 531168 579134
rect 530848 578866 531168 578898
rect 561568 579454 561888 579486
rect 561568 579218 561610 579454
rect 561846 579218 561888 579454
rect 561568 579134 561888 579218
rect 561568 578898 561610 579134
rect 561846 578898 561888 579134
rect 561568 578866 561888 578898
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 23968 561454 24288 561486
rect 23968 561218 24010 561454
rect 24246 561218 24288 561454
rect 23968 561134 24288 561218
rect 23968 560898 24010 561134
rect 24246 560898 24288 561134
rect 23968 560866 24288 560898
rect 54688 561454 55008 561486
rect 54688 561218 54730 561454
rect 54966 561218 55008 561454
rect 54688 561134 55008 561218
rect 54688 560898 54730 561134
rect 54966 560898 55008 561134
rect 54688 560866 55008 560898
rect 85408 561454 85728 561486
rect 85408 561218 85450 561454
rect 85686 561218 85728 561454
rect 85408 561134 85728 561218
rect 85408 560898 85450 561134
rect 85686 560898 85728 561134
rect 85408 560866 85728 560898
rect 116128 561454 116448 561486
rect 116128 561218 116170 561454
rect 116406 561218 116448 561454
rect 116128 561134 116448 561218
rect 116128 560898 116170 561134
rect 116406 560898 116448 561134
rect 116128 560866 116448 560898
rect 146848 561454 147168 561486
rect 146848 561218 146890 561454
rect 147126 561218 147168 561454
rect 146848 561134 147168 561218
rect 146848 560898 146890 561134
rect 147126 560898 147168 561134
rect 146848 560866 147168 560898
rect 177568 561454 177888 561486
rect 177568 561218 177610 561454
rect 177846 561218 177888 561454
rect 177568 561134 177888 561218
rect 177568 560898 177610 561134
rect 177846 560898 177888 561134
rect 177568 560866 177888 560898
rect 208288 561454 208608 561486
rect 208288 561218 208330 561454
rect 208566 561218 208608 561454
rect 208288 561134 208608 561218
rect 208288 560898 208330 561134
rect 208566 560898 208608 561134
rect 208288 560866 208608 560898
rect 239008 561454 239328 561486
rect 239008 561218 239050 561454
rect 239286 561218 239328 561454
rect 239008 561134 239328 561218
rect 239008 560898 239050 561134
rect 239286 560898 239328 561134
rect 239008 560866 239328 560898
rect 269728 561454 270048 561486
rect 269728 561218 269770 561454
rect 270006 561218 270048 561454
rect 269728 561134 270048 561218
rect 269728 560898 269770 561134
rect 270006 560898 270048 561134
rect 269728 560866 270048 560898
rect 300448 561454 300768 561486
rect 300448 561218 300490 561454
rect 300726 561218 300768 561454
rect 300448 561134 300768 561218
rect 300448 560898 300490 561134
rect 300726 560898 300768 561134
rect 300448 560866 300768 560898
rect 331168 561454 331488 561486
rect 331168 561218 331210 561454
rect 331446 561218 331488 561454
rect 331168 561134 331488 561218
rect 331168 560898 331210 561134
rect 331446 560898 331488 561134
rect 331168 560866 331488 560898
rect 361888 561454 362208 561486
rect 361888 561218 361930 561454
rect 362166 561218 362208 561454
rect 361888 561134 362208 561218
rect 361888 560898 361930 561134
rect 362166 560898 362208 561134
rect 361888 560866 362208 560898
rect 392608 561454 392928 561486
rect 392608 561218 392650 561454
rect 392886 561218 392928 561454
rect 392608 561134 392928 561218
rect 392608 560898 392650 561134
rect 392886 560898 392928 561134
rect 392608 560866 392928 560898
rect 423328 561454 423648 561486
rect 423328 561218 423370 561454
rect 423606 561218 423648 561454
rect 423328 561134 423648 561218
rect 423328 560898 423370 561134
rect 423606 560898 423648 561134
rect 423328 560866 423648 560898
rect 454048 561454 454368 561486
rect 454048 561218 454090 561454
rect 454326 561218 454368 561454
rect 454048 561134 454368 561218
rect 454048 560898 454090 561134
rect 454326 560898 454368 561134
rect 454048 560866 454368 560898
rect 484768 561454 485088 561486
rect 484768 561218 484810 561454
rect 485046 561218 485088 561454
rect 484768 561134 485088 561218
rect 484768 560898 484810 561134
rect 485046 560898 485088 561134
rect 484768 560866 485088 560898
rect 515488 561454 515808 561486
rect 515488 561218 515530 561454
rect 515766 561218 515808 561454
rect 515488 561134 515808 561218
rect 515488 560898 515530 561134
rect 515766 560898 515808 561134
rect 515488 560866 515808 560898
rect 546208 561454 546528 561486
rect 546208 561218 546250 561454
rect 546486 561218 546528 561454
rect 546208 561134 546528 561218
rect 546208 560898 546250 561134
rect 546486 560898 546528 561134
rect 546208 560866 546528 560898
rect 576928 561454 577248 561486
rect 576928 561218 576970 561454
rect 577206 561218 577248 561454
rect 576928 561134 577248 561218
rect 576928 560898 576970 561134
rect 577206 560898 577248 561134
rect 576928 560866 577248 560898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect 8608 543454 8928 543486
rect 8608 543218 8650 543454
rect 8886 543218 8928 543454
rect 8608 543134 8928 543218
rect 8608 542898 8650 543134
rect 8886 542898 8928 543134
rect 8608 542866 8928 542898
rect 39328 543454 39648 543486
rect 39328 543218 39370 543454
rect 39606 543218 39648 543454
rect 39328 543134 39648 543218
rect 39328 542898 39370 543134
rect 39606 542898 39648 543134
rect 39328 542866 39648 542898
rect 70048 543454 70368 543486
rect 70048 543218 70090 543454
rect 70326 543218 70368 543454
rect 70048 543134 70368 543218
rect 70048 542898 70090 543134
rect 70326 542898 70368 543134
rect 70048 542866 70368 542898
rect 100768 543454 101088 543486
rect 100768 543218 100810 543454
rect 101046 543218 101088 543454
rect 100768 543134 101088 543218
rect 100768 542898 100810 543134
rect 101046 542898 101088 543134
rect 100768 542866 101088 542898
rect 131488 543454 131808 543486
rect 131488 543218 131530 543454
rect 131766 543218 131808 543454
rect 131488 543134 131808 543218
rect 131488 542898 131530 543134
rect 131766 542898 131808 543134
rect 131488 542866 131808 542898
rect 162208 543454 162528 543486
rect 162208 543218 162250 543454
rect 162486 543218 162528 543454
rect 162208 543134 162528 543218
rect 162208 542898 162250 543134
rect 162486 542898 162528 543134
rect 162208 542866 162528 542898
rect 192928 543454 193248 543486
rect 192928 543218 192970 543454
rect 193206 543218 193248 543454
rect 192928 543134 193248 543218
rect 192928 542898 192970 543134
rect 193206 542898 193248 543134
rect 192928 542866 193248 542898
rect 223648 543454 223968 543486
rect 223648 543218 223690 543454
rect 223926 543218 223968 543454
rect 223648 543134 223968 543218
rect 223648 542898 223690 543134
rect 223926 542898 223968 543134
rect 223648 542866 223968 542898
rect 254368 543454 254688 543486
rect 254368 543218 254410 543454
rect 254646 543218 254688 543454
rect 254368 543134 254688 543218
rect 254368 542898 254410 543134
rect 254646 542898 254688 543134
rect 254368 542866 254688 542898
rect 285088 543454 285408 543486
rect 285088 543218 285130 543454
rect 285366 543218 285408 543454
rect 285088 543134 285408 543218
rect 285088 542898 285130 543134
rect 285366 542898 285408 543134
rect 285088 542866 285408 542898
rect 315808 543454 316128 543486
rect 315808 543218 315850 543454
rect 316086 543218 316128 543454
rect 315808 543134 316128 543218
rect 315808 542898 315850 543134
rect 316086 542898 316128 543134
rect 315808 542866 316128 542898
rect 346528 543454 346848 543486
rect 346528 543218 346570 543454
rect 346806 543218 346848 543454
rect 346528 543134 346848 543218
rect 346528 542898 346570 543134
rect 346806 542898 346848 543134
rect 346528 542866 346848 542898
rect 377248 543454 377568 543486
rect 377248 543218 377290 543454
rect 377526 543218 377568 543454
rect 377248 543134 377568 543218
rect 377248 542898 377290 543134
rect 377526 542898 377568 543134
rect 377248 542866 377568 542898
rect 407968 543454 408288 543486
rect 407968 543218 408010 543454
rect 408246 543218 408288 543454
rect 407968 543134 408288 543218
rect 407968 542898 408010 543134
rect 408246 542898 408288 543134
rect 407968 542866 408288 542898
rect 438688 543454 439008 543486
rect 438688 543218 438730 543454
rect 438966 543218 439008 543454
rect 438688 543134 439008 543218
rect 438688 542898 438730 543134
rect 438966 542898 439008 543134
rect 438688 542866 439008 542898
rect 469408 543454 469728 543486
rect 469408 543218 469450 543454
rect 469686 543218 469728 543454
rect 469408 543134 469728 543218
rect 469408 542898 469450 543134
rect 469686 542898 469728 543134
rect 469408 542866 469728 542898
rect 500128 543454 500448 543486
rect 500128 543218 500170 543454
rect 500406 543218 500448 543454
rect 500128 543134 500448 543218
rect 500128 542898 500170 543134
rect 500406 542898 500448 543134
rect 500128 542866 500448 542898
rect 530848 543454 531168 543486
rect 530848 543218 530890 543454
rect 531126 543218 531168 543454
rect 530848 543134 531168 543218
rect 530848 542898 530890 543134
rect 531126 542898 531168 543134
rect 530848 542866 531168 542898
rect 561568 543454 561888 543486
rect 561568 543218 561610 543454
rect 561846 543218 561888 543454
rect 561568 543134 561888 543218
rect 561568 542898 561610 543134
rect 561846 542898 561888 543134
rect 561568 542866 561888 542898
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 23968 525454 24288 525486
rect 23968 525218 24010 525454
rect 24246 525218 24288 525454
rect 23968 525134 24288 525218
rect 23968 524898 24010 525134
rect 24246 524898 24288 525134
rect 23968 524866 24288 524898
rect 54688 525454 55008 525486
rect 54688 525218 54730 525454
rect 54966 525218 55008 525454
rect 54688 525134 55008 525218
rect 54688 524898 54730 525134
rect 54966 524898 55008 525134
rect 54688 524866 55008 524898
rect 85408 525454 85728 525486
rect 85408 525218 85450 525454
rect 85686 525218 85728 525454
rect 85408 525134 85728 525218
rect 85408 524898 85450 525134
rect 85686 524898 85728 525134
rect 85408 524866 85728 524898
rect 116128 525454 116448 525486
rect 116128 525218 116170 525454
rect 116406 525218 116448 525454
rect 116128 525134 116448 525218
rect 116128 524898 116170 525134
rect 116406 524898 116448 525134
rect 116128 524866 116448 524898
rect 146848 525454 147168 525486
rect 146848 525218 146890 525454
rect 147126 525218 147168 525454
rect 146848 525134 147168 525218
rect 146848 524898 146890 525134
rect 147126 524898 147168 525134
rect 146848 524866 147168 524898
rect 177568 525454 177888 525486
rect 177568 525218 177610 525454
rect 177846 525218 177888 525454
rect 177568 525134 177888 525218
rect 177568 524898 177610 525134
rect 177846 524898 177888 525134
rect 177568 524866 177888 524898
rect 208288 525454 208608 525486
rect 208288 525218 208330 525454
rect 208566 525218 208608 525454
rect 208288 525134 208608 525218
rect 208288 524898 208330 525134
rect 208566 524898 208608 525134
rect 208288 524866 208608 524898
rect 239008 525454 239328 525486
rect 239008 525218 239050 525454
rect 239286 525218 239328 525454
rect 239008 525134 239328 525218
rect 239008 524898 239050 525134
rect 239286 524898 239328 525134
rect 239008 524866 239328 524898
rect 269728 525454 270048 525486
rect 269728 525218 269770 525454
rect 270006 525218 270048 525454
rect 269728 525134 270048 525218
rect 269728 524898 269770 525134
rect 270006 524898 270048 525134
rect 269728 524866 270048 524898
rect 300448 525454 300768 525486
rect 300448 525218 300490 525454
rect 300726 525218 300768 525454
rect 300448 525134 300768 525218
rect 300448 524898 300490 525134
rect 300726 524898 300768 525134
rect 300448 524866 300768 524898
rect 331168 525454 331488 525486
rect 331168 525218 331210 525454
rect 331446 525218 331488 525454
rect 331168 525134 331488 525218
rect 331168 524898 331210 525134
rect 331446 524898 331488 525134
rect 331168 524866 331488 524898
rect 361888 525454 362208 525486
rect 361888 525218 361930 525454
rect 362166 525218 362208 525454
rect 361888 525134 362208 525218
rect 361888 524898 361930 525134
rect 362166 524898 362208 525134
rect 361888 524866 362208 524898
rect 392608 525454 392928 525486
rect 392608 525218 392650 525454
rect 392886 525218 392928 525454
rect 392608 525134 392928 525218
rect 392608 524898 392650 525134
rect 392886 524898 392928 525134
rect 392608 524866 392928 524898
rect 423328 525454 423648 525486
rect 423328 525218 423370 525454
rect 423606 525218 423648 525454
rect 423328 525134 423648 525218
rect 423328 524898 423370 525134
rect 423606 524898 423648 525134
rect 423328 524866 423648 524898
rect 454048 525454 454368 525486
rect 454048 525218 454090 525454
rect 454326 525218 454368 525454
rect 454048 525134 454368 525218
rect 454048 524898 454090 525134
rect 454326 524898 454368 525134
rect 454048 524866 454368 524898
rect 484768 525454 485088 525486
rect 484768 525218 484810 525454
rect 485046 525218 485088 525454
rect 484768 525134 485088 525218
rect 484768 524898 484810 525134
rect 485046 524898 485088 525134
rect 484768 524866 485088 524898
rect 515488 525454 515808 525486
rect 515488 525218 515530 525454
rect 515766 525218 515808 525454
rect 515488 525134 515808 525218
rect 515488 524898 515530 525134
rect 515766 524898 515808 525134
rect 515488 524866 515808 524898
rect 546208 525454 546528 525486
rect 546208 525218 546250 525454
rect 546486 525218 546528 525454
rect 546208 525134 546528 525218
rect 546208 524898 546250 525134
rect 546486 524898 546528 525134
rect 546208 524866 546528 524898
rect 576928 525454 577248 525486
rect 576928 525218 576970 525454
rect 577206 525218 577248 525454
rect 576928 525134 577248 525218
rect 576928 524898 576970 525134
rect 577206 524898 577248 525134
rect 576928 524866 577248 524898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect 8608 507454 8928 507486
rect 8608 507218 8650 507454
rect 8886 507218 8928 507454
rect 8608 507134 8928 507218
rect 8608 506898 8650 507134
rect 8886 506898 8928 507134
rect 8608 506866 8928 506898
rect 39328 507454 39648 507486
rect 39328 507218 39370 507454
rect 39606 507218 39648 507454
rect 39328 507134 39648 507218
rect 39328 506898 39370 507134
rect 39606 506898 39648 507134
rect 39328 506866 39648 506898
rect 70048 507454 70368 507486
rect 70048 507218 70090 507454
rect 70326 507218 70368 507454
rect 70048 507134 70368 507218
rect 70048 506898 70090 507134
rect 70326 506898 70368 507134
rect 70048 506866 70368 506898
rect 100768 507454 101088 507486
rect 100768 507218 100810 507454
rect 101046 507218 101088 507454
rect 100768 507134 101088 507218
rect 100768 506898 100810 507134
rect 101046 506898 101088 507134
rect 100768 506866 101088 506898
rect 131488 507454 131808 507486
rect 131488 507218 131530 507454
rect 131766 507218 131808 507454
rect 131488 507134 131808 507218
rect 131488 506898 131530 507134
rect 131766 506898 131808 507134
rect 131488 506866 131808 506898
rect 162208 507454 162528 507486
rect 162208 507218 162250 507454
rect 162486 507218 162528 507454
rect 162208 507134 162528 507218
rect 162208 506898 162250 507134
rect 162486 506898 162528 507134
rect 162208 506866 162528 506898
rect 192928 507454 193248 507486
rect 192928 507218 192970 507454
rect 193206 507218 193248 507454
rect 192928 507134 193248 507218
rect 192928 506898 192970 507134
rect 193206 506898 193248 507134
rect 192928 506866 193248 506898
rect 223648 507454 223968 507486
rect 223648 507218 223690 507454
rect 223926 507218 223968 507454
rect 223648 507134 223968 507218
rect 223648 506898 223690 507134
rect 223926 506898 223968 507134
rect 223648 506866 223968 506898
rect 254368 507454 254688 507486
rect 254368 507218 254410 507454
rect 254646 507218 254688 507454
rect 254368 507134 254688 507218
rect 254368 506898 254410 507134
rect 254646 506898 254688 507134
rect 254368 506866 254688 506898
rect 285088 507454 285408 507486
rect 285088 507218 285130 507454
rect 285366 507218 285408 507454
rect 285088 507134 285408 507218
rect 285088 506898 285130 507134
rect 285366 506898 285408 507134
rect 285088 506866 285408 506898
rect 315808 507454 316128 507486
rect 315808 507218 315850 507454
rect 316086 507218 316128 507454
rect 315808 507134 316128 507218
rect 315808 506898 315850 507134
rect 316086 506898 316128 507134
rect 315808 506866 316128 506898
rect 346528 507454 346848 507486
rect 346528 507218 346570 507454
rect 346806 507218 346848 507454
rect 346528 507134 346848 507218
rect 346528 506898 346570 507134
rect 346806 506898 346848 507134
rect 346528 506866 346848 506898
rect 377248 507454 377568 507486
rect 377248 507218 377290 507454
rect 377526 507218 377568 507454
rect 377248 507134 377568 507218
rect 377248 506898 377290 507134
rect 377526 506898 377568 507134
rect 377248 506866 377568 506898
rect 407968 507454 408288 507486
rect 407968 507218 408010 507454
rect 408246 507218 408288 507454
rect 407968 507134 408288 507218
rect 407968 506898 408010 507134
rect 408246 506898 408288 507134
rect 407968 506866 408288 506898
rect 438688 507454 439008 507486
rect 438688 507218 438730 507454
rect 438966 507218 439008 507454
rect 438688 507134 439008 507218
rect 438688 506898 438730 507134
rect 438966 506898 439008 507134
rect 438688 506866 439008 506898
rect 469408 507454 469728 507486
rect 469408 507218 469450 507454
rect 469686 507218 469728 507454
rect 469408 507134 469728 507218
rect 469408 506898 469450 507134
rect 469686 506898 469728 507134
rect 469408 506866 469728 506898
rect 500128 507454 500448 507486
rect 500128 507218 500170 507454
rect 500406 507218 500448 507454
rect 500128 507134 500448 507218
rect 500128 506898 500170 507134
rect 500406 506898 500448 507134
rect 500128 506866 500448 506898
rect 530848 507454 531168 507486
rect 530848 507218 530890 507454
rect 531126 507218 531168 507454
rect 530848 507134 531168 507218
rect 530848 506898 530890 507134
rect 531126 506898 531168 507134
rect 530848 506866 531168 506898
rect 561568 507454 561888 507486
rect 561568 507218 561610 507454
rect 561846 507218 561888 507454
rect 561568 507134 561888 507218
rect 561568 506898 561610 507134
rect 561846 506898 561888 507134
rect 561568 506866 561888 506898
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 23968 489454 24288 489486
rect 23968 489218 24010 489454
rect 24246 489218 24288 489454
rect 23968 489134 24288 489218
rect 23968 488898 24010 489134
rect 24246 488898 24288 489134
rect 23968 488866 24288 488898
rect 54688 489454 55008 489486
rect 54688 489218 54730 489454
rect 54966 489218 55008 489454
rect 54688 489134 55008 489218
rect 54688 488898 54730 489134
rect 54966 488898 55008 489134
rect 54688 488866 55008 488898
rect 85408 489454 85728 489486
rect 85408 489218 85450 489454
rect 85686 489218 85728 489454
rect 85408 489134 85728 489218
rect 85408 488898 85450 489134
rect 85686 488898 85728 489134
rect 85408 488866 85728 488898
rect 116128 489454 116448 489486
rect 116128 489218 116170 489454
rect 116406 489218 116448 489454
rect 116128 489134 116448 489218
rect 116128 488898 116170 489134
rect 116406 488898 116448 489134
rect 116128 488866 116448 488898
rect 146848 489454 147168 489486
rect 146848 489218 146890 489454
rect 147126 489218 147168 489454
rect 146848 489134 147168 489218
rect 146848 488898 146890 489134
rect 147126 488898 147168 489134
rect 146848 488866 147168 488898
rect 177568 489454 177888 489486
rect 177568 489218 177610 489454
rect 177846 489218 177888 489454
rect 177568 489134 177888 489218
rect 177568 488898 177610 489134
rect 177846 488898 177888 489134
rect 177568 488866 177888 488898
rect 208288 489454 208608 489486
rect 208288 489218 208330 489454
rect 208566 489218 208608 489454
rect 208288 489134 208608 489218
rect 208288 488898 208330 489134
rect 208566 488898 208608 489134
rect 208288 488866 208608 488898
rect 239008 489454 239328 489486
rect 239008 489218 239050 489454
rect 239286 489218 239328 489454
rect 239008 489134 239328 489218
rect 239008 488898 239050 489134
rect 239286 488898 239328 489134
rect 239008 488866 239328 488898
rect 269728 489454 270048 489486
rect 269728 489218 269770 489454
rect 270006 489218 270048 489454
rect 269728 489134 270048 489218
rect 269728 488898 269770 489134
rect 270006 488898 270048 489134
rect 269728 488866 270048 488898
rect 300448 489454 300768 489486
rect 300448 489218 300490 489454
rect 300726 489218 300768 489454
rect 300448 489134 300768 489218
rect 300448 488898 300490 489134
rect 300726 488898 300768 489134
rect 300448 488866 300768 488898
rect 331168 489454 331488 489486
rect 331168 489218 331210 489454
rect 331446 489218 331488 489454
rect 331168 489134 331488 489218
rect 331168 488898 331210 489134
rect 331446 488898 331488 489134
rect 331168 488866 331488 488898
rect 361888 489454 362208 489486
rect 361888 489218 361930 489454
rect 362166 489218 362208 489454
rect 361888 489134 362208 489218
rect 361888 488898 361930 489134
rect 362166 488898 362208 489134
rect 361888 488866 362208 488898
rect 392608 489454 392928 489486
rect 392608 489218 392650 489454
rect 392886 489218 392928 489454
rect 392608 489134 392928 489218
rect 392608 488898 392650 489134
rect 392886 488898 392928 489134
rect 392608 488866 392928 488898
rect 423328 489454 423648 489486
rect 423328 489218 423370 489454
rect 423606 489218 423648 489454
rect 423328 489134 423648 489218
rect 423328 488898 423370 489134
rect 423606 488898 423648 489134
rect 423328 488866 423648 488898
rect 454048 489454 454368 489486
rect 454048 489218 454090 489454
rect 454326 489218 454368 489454
rect 454048 489134 454368 489218
rect 454048 488898 454090 489134
rect 454326 488898 454368 489134
rect 454048 488866 454368 488898
rect 484768 489454 485088 489486
rect 484768 489218 484810 489454
rect 485046 489218 485088 489454
rect 484768 489134 485088 489218
rect 484768 488898 484810 489134
rect 485046 488898 485088 489134
rect 484768 488866 485088 488898
rect 515488 489454 515808 489486
rect 515488 489218 515530 489454
rect 515766 489218 515808 489454
rect 515488 489134 515808 489218
rect 515488 488898 515530 489134
rect 515766 488898 515808 489134
rect 515488 488866 515808 488898
rect 546208 489454 546528 489486
rect 546208 489218 546250 489454
rect 546486 489218 546528 489454
rect 546208 489134 546528 489218
rect 546208 488898 546250 489134
rect 546486 488898 546528 489134
rect 546208 488866 546528 488898
rect 576928 489454 577248 489486
rect 576928 489218 576970 489454
rect 577206 489218 577248 489454
rect 576928 489134 577248 489218
rect 576928 488898 576970 489134
rect 577206 488898 577248 489134
rect 576928 488866 577248 488898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect 8608 471454 8928 471486
rect 8608 471218 8650 471454
rect 8886 471218 8928 471454
rect 8608 471134 8928 471218
rect 8608 470898 8650 471134
rect 8886 470898 8928 471134
rect 8608 470866 8928 470898
rect 39328 471454 39648 471486
rect 39328 471218 39370 471454
rect 39606 471218 39648 471454
rect 39328 471134 39648 471218
rect 39328 470898 39370 471134
rect 39606 470898 39648 471134
rect 39328 470866 39648 470898
rect 70048 471454 70368 471486
rect 70048 471218 70090 471454
rect 70326 471218 70368 471454
rect 70048 471134 70368 471218
rect 70048 470898 70090 471134
rect 70326 470898 70368 471134
rect 70048 470866 70368 470898
rect 100768 471454 101088 471486
rect 100768 471218 100810 471454
rect 101046 471218 101088 471454
rect 100768 471134 101088 471218
rect 100768 470898 100810 471134
rect 101046 470898 101088 471134
rect 100768 470866 101088 470898
rect 131488 471454 131808 471486
rect 131488 471218 131530 471454
rect 131766 471218 131808 471454
rect 131488 471134 131808 471218
rect 131488 470898 131530 471134
rect 131766 470898 131808 471134
rect 131488 470866 131808 470898
rect 162208 471454 162528 471486
rect 162208 471218 162250 471454
rect 162486 471218 162528 471454
rect 162208 471134 162528 471218
rect 162208 470898 162250 471134
rect 162486 470898 162528 471134
rect 162208 470866 162528 470898
rect 192928 471454 193248 471486
rect 192928 471218 192970 471454
rect 193206 471218 193248 471454
rect 192928 471134 193248 471218
rect 192928 470898 192970 471134
rect 193206 470898 193248 471134
rect 192928 470866 193248 470898
rect 223648 471454 223968 471486
rect 223648 471218 223690 471454
rect 223926 471218 223968 471454
rect 223648 471134 223968 471218
rect 223648 470898 223690 471134
rect 223926 470898 223968 471134
rect 223648 470866 223968 470898
rect 254368 471454 254688 471486
rect 254368 471218 254410 471454
rect 254646 471218 254688 471454
rect 254368 471134 254688 471218
rect 254368 470898 254410 471134
rect 254646 470898 254688 471134
rect 254368 470866 254688 470898
rect 285088 471454 285408 471486
rect 285088 471218 285130 471454
rect 285366 471218 285408 471454
rect 285088 471134 285408 471218
rect 285088 470898 285130 471134
rect 285366 470898 285408 471134
rect 285088 470866 285408 470898
rect 315808 471454 316128 471486
rect 315808 471218 315850 471454
rect 316086 471218 316128 471454
rect 315808 471134 316128 471218
rect 315808 470898 315850 471134
rect 316086 470898 316128 471134
rect 315808 470866 316128 470898
rect 346528 471454 346848 471486
rect 346528 471218 346570 471454
rect 346806 471218 346848 471454
rect 346528 471134 346848 471218
rect 346528 470898 346570 471134
rect 346806 470898 346848 471134
rect 346528 470866 346848 470898
rect 377248 471454 377568 471486
rect 377248 471218 377290 471454
rect 377526 471218 377568 471454
rect 377248 471134 377568 471218
rect 377248 470898 377290 471134
rect 377526 470898 377568 471134
rect 377248 470866 377568 470898
rect 407968 471454 408288 471486
rect 407968 471218 408010 471454
rect 408246 471218 408288 471454
rect 407968 471134 408288 471218
rect 407968 470898 408010 471134
rect 408246 470898 408288 471134
rect 407968 470866 408288 470898
rect 438688 471454 439008 471486
rect 438688 471218 438730 471454
rect 438966 471218 439008 471454
rect 438688 471134 439008 471218
rect 438688 470898 438730 471134
rect 438966 470898 439008 471134
rect 438688 470866 439008 470898
rect 469408 471454 469728 471486
rect 469408 471218 469450 471454
rect 469686 471218 469728 471454
rect 469408 471134 469728 471218
rect 469408 470898 469450 471134
rect 469686 470898 469728 471134
rect 469408 470866 469728 470898
rect 500128 471454 500448 471486
rect 500128 471218 500170 471454
rect 500406 471218 500448 471454
rect 500128 471134 500448 471218
rect 500128 470898 500170 471134
rect 500406 470898 500448 471134
rect 500128 470866 500448 470898
rect 530848 471454 531168 471486
rect 530848 471218 530890 471454
rect 531126 471218 531168 471454
rect 530848 471134 531168 471218
rect 530848 470898 530890 471134
rect 531126 470898 531168 471134
rect 530848 470866 531168 470898
rect 561568 471454 561888 471486
rect 561568 471218 561610 471454
rect 561846 471218 561888 471454
rect 561568 471134 561888 471218
rect 561568 470898 561610 471134
rect 561846 470898 561888 471134
rect 561568 470866 561888 470898
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 23968 453454 24288 453486
rect 23968 453218 24010 453454
rect 24246 453218 24288 453454
rect 23968 453134 24288 453218
rect 23968 452898 24010 453134
rect 24246 452898 24288 453134
rect 23968 452866 24288 452898
rect 54688 453454 55008 453486
rect 54688 453218 54730 453454
rect 54966 453218 55008 453454
rect 54688 453134 55008 453218
rect 54688 452898 54730 453134
rect 54966 452898 55008 453134
rect 54688 452866 55008 452898
rect 85408 453454 85728 453486
rect 85408 453218 85450 453454
rect 85686 453218 85728 453454
rect 85408 453134 85728 453218
rect 85408 452898 85450 453134
rect 85686 452898 85728 453134
rect 85408 452866 85728 452898
rect 116128 453454 116448 453486
rect 116128 453218 116170 453454
rect 116406 453218 116448 453454
rect 116128 453134 116448 453218
rect 116128 452898 116170 453134
rect 116406 452898 116448 453134
rect 116128 452866 116448 452898
rect 146848 453454 147168 453486
rect 146848 453218 146890 453454
rect 147126 453218 147168 453454
rect 146848 453134 147168 453218
rect 146848 452898 146890 453134
rect 147126 452898 147168 453134
rect 146848 452866 147168 452898
rect 177568 453454 177888 453486
rect 177568 453218 177610 453454
rect 177846 453218 177888 453454
rect 177568 453134 177888 453218
rect 177568 452898 177610 453134
rect 177846 452898 177888 453134
rect 177568 452866 177888 452898
rect 208288 453454 208608 453486
rect 208288 453218 208330 453454
rect 208566 453218 208608 453454
rect 208288 453134 208608 453218
rect 208288 452898 208330 453134
rect 208566 452898 208608 453134
rect 208288 452866 208608 452898
rect 239008 453454 239328 453486
rect 239008 453218 239050 453454
rect 239286 453218 239328 453454
rect 239008 453134 239328 453218
rect 239008 452898 239050 453134
rect 239286 452898 239328 453134
rect 239008 452866 239328 452898
rect 269728 453454 270048 453486
rect 269728 453218 269770 453454
rect 270006 453218 270048 453454
rect 269728 453134 270048 453218
rect 269728 452898 269770 453134
rect 270006 452898 270048 453134
rect 269728 452866 270048 452898
rect 300448 453454 300768 453486
rect 300448 453218 300490 453454
rect 300726 453218 300768 453454
rect 300448 453134 300768 453218
rect 300448 452898 300490 453134
rect 300726 452898 300768 453134
rect 300448 452866 300768 452898
rect 331168 453454 331488 453486
rect 331168 453218 331210 453454
rect 331446 453218 331488 453454
rect 331168 453134 331488 453218
rect 331168 452898 331210 453134
rect 331446 452898 331488 453134
rect 331168 452866 331488 452898
rect 361888 453454 362208 453486
rect 361888 453218 361930 453454
rect 362166 453218 362208 453454
rect 361888 453134 362208 453218
rect 361888 452898 361930 453134
rect 362166 452898 362208 453134
rect 361888 452866 362208 452898
rect 392608 453454 392928 453486
rect 392608 453218 392650 453454
rect 392886 453218 392928 453454
rect 392608 453134 392928 453218
rect 392608 452898 392650 453134
rect 392886 452898 392928 453134
rect 392608 452866 392928 452898
rect 423328 453454 423648 453486
rect 423328 453218 423370 453454
rect 423606 453218 423648 453454
rect 423328 453134 423648 453218
rect 423328 452898 423370 453134
rect 423606 452898 423648 453134
rect 423328 452866 423648 452898
rect 454048 453454 454368 453486
rect 454048 453218 454090 453454
rect 454326 453218 454368 453454
rect 454048 453134 454368 453218
rect 454048 452898 454090 453134
rect 454326 452898 454368 453134
rect 454048 452866 454368 452898
rect 484768 453454 485088 453486
rect 484768 453218 484810 453454
rect 485046 453218 485088 453454
rect 484768 453134 485088 453218
rect 484768 452898 484810 453134
rect 485046 452898 485088 453134
rect 484768 452866 485088 452898
rect 515488 453454 515808 453486
rect 515488 453218 515530 453454
rect 515766 453218 515808 453454
rect 515488 453134 515808 453218
rect 515488 452898 515530 453134
rect 515766 452898 515808 453134
rect 515488 452866 515808 452898
rect 546208 453454 546528 453486
rect 546208 453218 546250 453454
rect 546486 453218 546528 453454
rect 546208 453134 546528 453218
rect 546208 452898 546250 453134
rect 546486 452898 546528 453134
rect 546208 452866 546528 452898
rect 576928 453454 577248 453486
rect 576928 453218 576970 453454
rect 577206 453218 577248 453454
rect 576928 453134 577248 453218
rect 576928 452898 576970 453134
rect 577206 452898 577248 453134
rect 576928 452866 577248 452898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect 8608 435454 8928 435486
rect 8608 435218 8650 435454
rect 8886 435218 8928 435454
rect 8608 435134 8928 435218
rect 8608 434898 8650 435134
rect 8886 434898 8928 435134
rect 8608 434866 8928 434898
rect 39328 435454 39648 435486
rect 39328 435218 39370 435454
rect 39606 435218 39648 435454
rect 39328 435134 39648 435218
rect 39328 434898 39370 435134
rect 39606 434898 39648 435134
rect 39328 434866 39648 434898
rect 70048 435454 70368 435486
rect 70048 435218 70090 435454
rect 70326 435218 70368 435454
rect 70048 435134 70368 435218
rect 70048 434898 70090 435134
rect 70326 434898 70368 435134
rect 70048 434866 70368 434898
rect 100768 435454 101088 435486
rect 100768 435218 100810 435454
rect 101046 435218 101088 435454
rect 100768 435134 101088 435218
rect 100768 434898 100810 435134
rect 101046 434898 101088 435134
rect 100768 434866 101088 434898
rect 131488 435454 131808 435486
rect 131488 435218 131530 435454
rect 131766 435218 131808 435454
rect 131488 435134 131808 435218
rect 131488 434898 131530 435134
rect 131766 434898 131808 435134
rect 131488 434866 131808 434898
rect 162208 435454 162528 435486
rect 162208 435218 162250 435454
rect 162486 435218 162528 435454
rect 162208 435134 162528 435218
rect 162208 434898 162250 435134
rect 162486 434898 162528 435134
rect 162208 434866 162528 434898
rect 192928 435454 193248 435486
rect 192928 435218 192970 435454
rect 193206 435218 193248 435454
rect 192928 435134 193248 435218
rect 192928 434898 192970 435134
rect 193206 434898 193248 435134
rect 192928 434866 193248 434898
rect 223648 435454 223968 435486
rect 223648 435218 223690 435454
rect 223926 435218 223968 435454
rect 223648 435134 223968 435218
rect 223648 434898 223690 435134
rect 223926 434898 223968 435134
rect 223648 434866 223968 434898
rect 254368 435454 254688 435486
rect 254368 435218 254410 435454
rect 254646 435218 254688 435454
rect 254368 435134 254688 435218
rect 254368 434898 254410 435134
rect 254646 434898 254688 435134
rect 254368 434866 254688 434898
rect 285088 435454 285408 435486
rect 285088 435218 285130 435454
rect 285366 435218 285408 435454
rect 285088 435134 285408 435218
rect 285088 434898 285130 435134
rect 285366 434898 285408 435134
rect 285088 434866 285408 434898
rect 315808 435454 316128 435486
rect 315808 435218 315850 435454
rect 316086 435218 316128 435454
rect 315808 435134 316128 435218
rect 315808 434898 315850 435134
rect 316086 434898 316128 435134
rect 315808 434866 316128 434898
rect 346528 435454 346848 435486
rect 346528 435218 346570 435454
rect 346806 435218 346848 435454
rect 346528 435134 346848 435218
rect 346528 434898 346570 435134
rect 346806 434898 346848 435134
rect 346528 434866 346848 434898
rect 377248 435454 377568 435486
rect 377248 435218 377290 435454
rect 377526 435218 377568 435454
rect 377248 435134 377568 435218
rect 377248 434898 377290 435134
rect 377526 434898 377568 435134
rect 377248 434866 377568 434898
rect 407968 435454 408288 435486
rect 407968 435218 408010 435454
rect 408246 435218 408288 435454
rect 407968 435134 408288 435218
rect 407968 434898 408010 435134
rect 408246 434898 408288 435134
rect 407968 434866 408288 434898
rect 438688 435454 439008 435486
rect 438688 435218 438730 435454
rect 438966 435218 439008 435454
rect 438688 435134 439008 435218
rect 438688 434898 438730 435134
rect 438966 434898 439008 435134
rect 438688 434866 439008 434898
rect 469408 435454 469728 435486
rect 469408 435218 469450 435454
rect 469686 435218 469728 435454
rect 469408 435134 469728 435218
rect 469408 434898 469450 435134
rect 469686 434898 469728 435134
rect 469408 434866 469728 434898
rect 500128 435454 500448 435486
rect 500128 435218 500170 435454
rect 500406 435218 500448 435454
rect 500128 435134 500448 435218
rect 500128 434898 500170 435134
rect 500406 434898 500448 435134
rect 500128 434866 500448 434898
rect 530848 435454 531168 435486
rect 530848 435218 530890 435454
rect 531126 435218 531168 435454
rect 530848 435134 531168 435218
rect 530848 434898 530890 435134
rect 531126 434898 531168 435134
rect 530848 434866 531168 434898
rect 561568 435454 561888 435486
rect 561568 435218 561610 435454
rect 561846 435218 561888 435454
rect 561568 435134 561888 435218
rect 561568 434898 561610 435134
rect 561846 434898 561888 435134
rect 561568 434866 561888 434898
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 23968 417454 24288 417486
rect 23968 417218 24010 417454
rect 24246 417218 24288 417454
rect 23968 417134 24288 417218
rect 23968 416898 24010 417134
rect 24246 416898 24288 417134
rect 23968 416866 24288 416898
rect 54688 417454 55008 417486
rect 54688 417218 54730 417454
rect 54966 417218 55008 417454
rect 54688 417134 55008 417218
rect 54688 416898 54730 417134
rect 54966 416898 55008 417134
rect 54688 416866 55008 416898
rect 85408 417454 85728 417486
rect 85408 417218 85450 417454
rect 85686 417218 85728 417454
rect 85408 417134 85728 417218
rect 85408 416898 85450 417134
rect 85686 416898 85728 417134
rect 85408 416866 85728 416898
rect 116128 417454 116448 417486
rect 116128 417218 116170 417454
rect 116406 417218 116448 417454
rect 116128 417134 116448 417218
rect 116128 416898 116170 417134
rect 116406 416898 116448 417134
rect 116128 416866 116448 416898
rect 146848 417454 147168 417486
rect 146848 417218 146890 417454
rect 147126 417218 147168 417454
rect 146848 417134 147168 417218
rect 146848 416898 146890 417134
rect 147126 416898 147168 417134
rect 146848 416866 147168 416898
rect 177568 417454 177888 417486
rect 177568 417218 177610 417454
rect 177846 417218 177888 417454
rect 177568 417134 177888 417218
rect 177568 416898 177610 417134
rect 177846 416898 177888 417134
rect 177568 416866 177888 416898
rect 208288 417454 208608 417486
rect 208288 417218 208330 417454
rect 208566 417218 208608 417454
rect 208288 417134 208608 417218
rect 208288 416898 208330 417134
rect 208566 416898 208608 417134
rect 208288 416866 208608 416898
rect 239008 417454 239328 417486
rect 239008 417218 239050 417454
rect 239286 417218 239328 417454
rect 239008 417134 239328 417218
rect 239008 416898 239050 417134
rect 239286 416898 239328 417134
rect 239008 416866 239328 416898
rect 269728 417454 270048 417486
rect 269728 417218 269770 417454
rect 270006 417218 270048 417454
rect 269728 417134 270048 417218
rect 269728 416898 269770 417134
rect 270006 416898 270048 417134
rect 269728 416866 270048 416898
rect 300448 417454 300768 417486
rect 300448 417218 300490 417454
rect 300726 417218 300768 417454
rect 300448 417134 300768 417218
rect 300448 416898 300490 417134
rect 300726 416898 300768 417134
rect 300448 416866 300768 416898
rect 331168 417454 331488 417486
rect 331168 417218 331210 417454
rect 331446 417218 331488 417454
rect 331168 417134 331488 417218
rect 331168 416898 331210 417134
rect 331446 416898 331488 417134
rect 331168 416866 331488 416898
rect 361888 417454 362208 417486
rect 361888 417218 361930 417454
rect 362166 417218 362208 417454
rect 361888 417134 362208 417218
rect 361888 416898 361930 417134
rect 362166 416898 362208 417134
rect 361888 416866 362208 416898
rect 392608 417454 392928 417486
rect 392608 417218 392650 417454
rect 392886 417218 392928 417454
rect 392608 417134 392928 417218
rect 392608 416898 392650 417134
rect 392886 416898 392928 417134
rect 392608 416866 392928 416898
rect 423328 417454 423648 417486
rect 423328 417218 423370 417454
rect 423606 417218 423648 417454
rect 423328 417134 423648 417218
rect 423328 416898 423370 417134
rect 423606 416898 423648 417134
rect 423328 416866 423648 416898
rect 454048 417454 454368 417486
rect 454048 417218 454090 417454
rect 454326 417218 454368 417454
rect 454048 417134 454368 417218
rect 454048 416898 454090 417134
rect 454326 416898 454368 417134
rect 454048 416866 454368 416898
rect 484768 417454 485088 417486
rect 484768 417218 484810 417454
rect 485046 417218 485088 417454
rect 484768 417134 485088 417218
rect 484768 416898 484810 417134
rect 485046 416898 485088 417134
rect 484768 416866 485088 416898
rect 515488 417454 515808 417486
rect 515488 417218 515530 417454
rect 515766 417218 515808 417454
rect 515488 417134 515808 417218
rect 515488 416898 515530 417134
rect 515766 416898 515808 417134
rect 515488 416866 515808 416898
rect 546208 417454 546528 417486
rect 546208 417218 546250 417454
rect 546486 417218 546528 417454
rect 546208 417134 546528 417218
rect 546208 416898 546250 417134
rect 546486 416898 546528 417134
rect 546208 416866 546528 416898
rect 576928 417454 577248 417486
rect 576928 417218 576970 417454
rect 577206 417218 577248 417454
rect 576928 417134 577248 417218
rect 576928 416898 576970 417134
rect 577206 416898 577248 417134
rect 576928 416866 577248 416898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect 8608 399454 8928 399486
rect 8608 399218 8650 399454
rect 8886 399218 8928 399454
rect 8608 399134 8928 399218
rect 8608 398898 8650 399134
rect 8886 398898 8928 399134
rect 8608 398866 8928 398898
rect 39328 399454 39648 399486
rect 39328 399218 39370 399454
rect 39606 399218 39648 399454
rect 39328 399134 39648 399218
rect 39328 398898 39370 399134
rect 39606 398898 39648 399134
rect 39328 398866 39648 398898
rect 70048 399454 70368 399486
rect 70048 399218 70090 399454
rect 70326 399218 70368 399454
rect 70048 399134 70368 399218
rect 70048 398898 70090 399134
rect 70326 398898 70368 399134
rect 70048 398866 70368 398898
rect 100768 399454 101088 399486
rect 100768 399218 100810 399454
rect 101046 399218 101088 399454
rect 100768 399134 101088 399218
rect 100768 398898 100810 399134
rect 101046 398898 101088 399134
rect 100768 398866 101088 398898
rect 131488 399454 131808 399486
rect 131488 399218 131530 399454
rect 131766 399218 131808 399454
rect 131488 399134 131808 399218
rect 131488 398898 131530 399134
rect 131766 398898 131808 399134
rect 131488 398866 131808 398898
rect 162208 399454 162528 399486
rect 162208 399218 162250 399454
rect 162486 399218 162528 399454
rect 162208 399134 162528 399218
rect 162208 398898 162250 399134
rect 162486 398898 162528 399134
rect 162208 398866 162528 398898
rect 192928 399454 193248 399486
rect 192928 399218 192970 399454
rect 193206 399218 193248 399454
rect 192928 399134 193248 399218
rect 192928 398898 192970 399134
rect 193206 398898 193248 399134
rect 192928 398866 193248 398898
rect 223648 399454 223968 399486
rect 223648 399218 223690 399454
rect 223926 399218 223968 399454
rect 223648 399134 223968 399218
rect 223648 398898 223690 399134
rect 223926 398898 223968 399134
rect 223648 398866 223968 398898
rect 254368 399454 254688 399486
rect 254368 399218 254410 399454
rect 254646 399218 254688 399454
rect 254368 399134 254688 399218
rect 254368 398898 254410 399134
rect 254646 398898 254688 399134
rect 254368 398866 254688 398898
rect 285088 399454 285408 399486
rect 285088 399218 285130 399454
rect 285366 399218 285408 399454
rect 285088 399134 285408 399218
rect 285088 398898 285130 399134
rect 285366 398898 285408 399134
rect 285088 398866 285408 398898
rect 315808 399454 316128 399486
rect 315808 399218 315850 399454
rect 316086 399218 316128 399454
rect 315808 399134 316128 399218
rect 315808 398898 315850 399134
rect 316086 398898 316128 399134
rect 315808 398866 316128 398898
rect 346528 399454 346848 399486
rect 346528 399218 346570 399454
rect 346806 399218 346848 399454
rect 346528 399134 346848 399218
rect 346528 398898 346570 399134
rect 346806 398898 346848 399134
rect 346528 398866 346848 398898
rect 377248 399454 377568 399486
rect 377248 399218 377290 399454
rect 377526 399218 377568 399454
rect 377248 399134 377568 399218
rect 377248 398898 377290 399134
rect 377526 398898 377568 399134
rect 377248 398866 377568 398898
rect 407968 399454 408288 399486
rect 407968 399218 408010 399454
rect 408246 399218 408288 399454
rect 407968 399134 408288 399218
rect 407968 398898 408010 399134
rect 408246 398898 408288 399134
rect 407968 398866 408288 398898
rect 438688 399454 439008 399486
rect 438688 399218 438730 399454
rect 438966 399218 439008 399454
rect 438688 399134 439008 399218
rect 438688 398898 438730 399134
rect 438966 398898 439008 399134
rect 438688 398866 439008 398898
rect 469408 399454 469728 399486
rect 469408 399218 469450 399454
rect 469686 399218 469728 399454
rect 469408 399134 469728 399218
rect 469408 398898 469450 399134
rect 469686 398898 469728 399134
rect 469408 398866 469728 398898
rect 500128 399454 500448 399486
rect 500128 399218 500170 399454
rect 500406 399218 500448 399454
rect 500128 399134 500448 399218
rect 500128 398898 500170 399134
rect 500406 398898 500448 399134
rect 500128 398866 500448 398898
rect 530848 399454 531168 399486
rect 530848 399218 530890 399454
rect 531126 399218 531168 399454
rect 530848 399134 531168 399218
rect 530848 398898 530890 399134
rect 531126 398898 531168 399134
rect 530848 398866 531168 398898
rect 561568 399454 561888 399486
rect 561568 399218 561610 399454
rect 561846 399218 561888 399454
rect 561568 399134 561888 399218
rect 561568 398898 561610 399134
rect 561846 398898 561888 399134
rect 561568 398866 561888 398898
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 23968 381454 24288 381486
rect 23968 381218 24010 381454
rect 24246 381218 24288 381454
rect 23968 381134 24288 381218
rect 23968 380898 24010 381134
rect 24246 380898 24288 381134
rect 23968 380866 24288 380898
rect 54688 381454 55008 381486
rect 54688 381218 54730 381454
rect 54966 381218 55008 381454
rect 54688 381134 55008 381218
rect 54688 380898 54730 381134
rect 54966 380898 55008 381134
rect 54688 380866 55008 380898
rect 85408 381454 85728 381486
rect 85408 381218 85450 381454
rect 85686 381218 85728 381454
rect 85408 381134 85728 381218
rect 85408 380898 85450 381134
rect 85686 380898 85728 381134
rect 85408 380866 85728 380898
rect 116128 381454 116448 381486
rect 116128 381218 116170 381454
rect 116406 381218 116448 381454
rect 116128 381134 116448 381218
rect 116128 380898 116170 381134
rect 116406 380898 116448 381134
rect 116128 380866 116448 380898
rect 146848 381454 147168 381486
rect 146848 381218 146890 381454
rect 147126 381218 147168 381454
rect 146848 381134 147168 381218
rect 146848 380898 146890 381134
rect 147126 380898 147168 381134
rect 146848 380866 147168 380898
rect 177568 381454 177888 381486
rect 177568 381218 177610 381454
rect 177846 381218 177888 381454
rect 177568 381134 177888 381218
rect 177568 380898 177610 381134
rect 177846 380898 177888 381134
rect 177568 380866 177888 380898
rect 208288 381454 208608 381486
rect 208288 381218 208330 381454
rect 208566 381218 208608 381454
rect 208288 381134 208608 381218
rect 208288 380898 208330 381134
rect 208566 380898 208608 381134
rect 208288 380866 208608 380898
rect 239008 381454 239328 381486
rect 239008 381218 239050 381454
rect 239286 381218 239328 381454
rect 239008 381134 239328 381218
rect 239008 380898 239050 381134
rect 239286 380898 239328 381134
rect 239008 380866 239328 380898
rect 269728 381454 270048 381486
rect 269728 381218 269770 381454
rect 270006 381218 270048 381454
rect 269728 381134 270048 381218
rect 269728 380898 269770 381134
rect 270006 380898 270048 381134
rect 269728 380866 270048 380898
rect 300448 381454 300768 381486
rect 300448 381218 300490 381454
rect 300726 381218 300768 381454
rect 300448 381134 300768 381218
rect 300448 380898 300490 381134
rect 300726 380898 300768 381134
rect 300448 380866 300768 380898
rect 331168 381454 331488 381486
rect 331168 381218 331210 381454
rect 331446 381218 331488 381454
rect 331168 381134 331488 381218
rect 331168 380898 331210 381134
rect 331446 380898 331488 381134
rect 331168 380866 331488 380898
rect 361888 381454 362208 381486
rect 361888 381218 361930 381454
rect 362166 381218 362208 381454
rect 361888 381134 362208 381218
rect 361888 380898 361930 381134
rect 362166 380898 362208 381134
rect 361888 380866 362208 380898
rect 392608 381454 392928 381486
rect 392608 381218 392650 381454
rect 392886 381218 392928 381454
rect 392608 381134 392928 381218
rect 392608 380898 392650 381134
rect 392886 380898 392928 381134
rect 392608 380866 392928 380898
rect 423328 381454 423648 381486
rect 423328 381218 423370 381454
rect 423606 381218 423648 381454
rect 423328 381134 423648 381218
rect 423328 380898 423370 381134
rect 423606 380898 423648 381134
rect 423328 380866 423648 380898
rect 454048 381454 454368 381486
rect 454048 381218 454090 381454
rect 454326 381218 454368 381454
rect 454048 381134 454368 381218
rect 454048 380898 454090 381134
rect 454326 380898 454368 381134
rect 454048 380866 454368 380898
rect 484768 381454 485088 381486
rect 484768 381218 484810 381454
rect 485046 381218 485088 381454
rect 484768 381134 485088 381218
rect 484768 380898 484810 381134
rect 485046 380898 485088 381134
rect 484768 380866 485088 380898
rect 515488 381454 515808 381486
rect 515488 381218 515530 381454
rect 515766 381218 515808 381454
rect 515488 381134 515808 381218
rect 515488 380898 515530 381134
rect 515766 380898 515808 381134
rect 515488 380866 515808 380898
rect 546208 381454 546528 381486
rect 546208 381218 546250 381454
rect 546486 381218 546528 381454
rect 546208 381134 546528 381218
rect 546208 380898 546250 381134
rect 546486 380898 546528 381134
rect 546208 380866 546528 380898
rect 576928 381454 577248 381486
rect 576928 381218 576970 381454
rect 577206 381218 577248 381454
rect 576928 381134 577248 381218
rect 576928 380898 576970 381134
rect 577206 380898 577248 381134
rect 576928 380866 577248 380898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect 8608 363454 8928 363486
rect 8608 363218 8650 363454
rect 8886 363218 8928 363454
rect 8608 363134 8928 363218
rect 8608 362898 8650 363134
rect 8886 362898 8928 363134
rect 8608 362866 8928 362898
rect 39328 363454 39648 363486
rect 39328 363218 39370 363454
rect 39606 363218 39648 363454
rect 39328 363134 39648 363218
rect 39328 362898 39370 363134
rect 39606 362898 39648 363134
rect 39328 362866 39648 362898
rect 70048 363454 70368 363486
rect 70048 363218 70090 363454
rect 70326 363218 70368 363454
rect 70048 363134 70368 363218
rect 70048 362898 70090 363134
rect 70326 362898 70368 363134
rect 70048 362866 70368 362898
rect 100768 363454 101088 363486
rect 100768 363218 100810 363454
rect 101046 363218 101088 363454
rect 100768 363134 101088 363218
rect 100768 362898 100810 363134
rect 101046 362898 101088 363134
rect 100768 362866 101088 362898
rect 131488 363454 131808 363486
rect 131488 363218 131530 363454
rect 131766 363218 131808 363454
rect 131488 363134 131808 363218
rect 131488 362898 131530 363134
rect 131766 362898 131808 363134
rect 131488 362866 131808 362898
rect 162208 363454 162528 363486
rect 162208 363218 162250 363454
rect 162486 363218 162528 363454
rect 162208 363134 162528 363218
rect 162208 362898 162250 363134
rect 162486 362898 162528 363134
rect 162208 362866 162528 362898
rect 192928 363454 193248 363486
rect 192928 363218 192970 363454
rect 193206 363218 193248 363454
rect 192928 363134 193248 363218
rect 192928 362898 192970 363134
rect 193206 362898 193248 363134
rect 192928 362866 193248 362898
rect 223648 363454 223968 363486
rect 223648 363218 223690 363454
rect 223926 363218 223968 363454
rect 223648 363134 223968 363218
rect 223648 362898 223690 363134
rect 223926 362898 223968 363134
rect 223648 362866 223968 362898
rect 254368 363454 254688 363486
rect 254368 363218 254410 363454
rect 254646 363218 254688 363454
rect 254368 363134 254688 363218
rect 254368 362898 254410 363134
rect 254646 362898 254688 363134
rect 254368 362866 254688 362898
rect 285088 363454 285408 363486
rect 285088 363218 285130 363454
rect 285366 363218 285408 363454
rect 285088 363134 285408 363218
rect 285088 362898 285130 363134
rect 285366 362898 285408 363134
rect 285088 362866 285408 362898
rect 315808 363454 316128 363486
rect 315808 363218 315850 363454
rect 316086 363218 316128 363454
rect 315808 363134 316128 363218
rect 315808 362898 315850 363134
rect 316086 362898 316128 363134
rect 315808 362866 316128 362898
rect 346528 363454 346848 363486
rect 346528 363218 346570 363454
rect 346806 363218 346848 363454
rect 346528 363134 346848 363218
rect 346528 362898 346570 363134
rect 346806 362898 346848 363134
rect 346528 362866 346848 362898
rect 377248 363454 377568 363486
rect 377248 363218 377290 363454
rect 377526 363218 377568 363454
rect 377248 363134 377568 363218
rect 377248 362898 377290 363134
rect 377526 362898 377568 363134
rect 377248 362866 377568 362898
rect 407968 363454 408288 363486
rect 407968 363218 408010 363454
rect 408246 363218 408288 363454
rect 407968 363134 408288 363218
rect 407968 362898 408010 363134
rect 408246 362898 408288 363134
rect 407968 362866 408288 362898
rect 438688 363454 439008 363486
rect 438688 363218 438730 363454
rect 438966 363218 439008 363454
rect 438688 363134 439008 363218
rect 438688 362898 438730 363134
rect 438966 362898 439008 363134
rect 438688 362866 439008 362898
rect 469408 363454 469728 363486
rect 469408 363218 469450 363454
rect 469686 363218 469728 363454
rect 469408 363134 469728 363218
rect 469408 362898 469450 363134
rect 469686 362898 469728 363134
rect 469408 362866 469728 362898
rect 500128 363454 500448 363486
rect 500128 363218 500170 363454
rect 500406 363218 500448 363454
rect 500128 363134 500448 363218
rect 500128 362898 500170 363134
rect 500406 362898 500448 363134
rect 500128 362866 500448 362898
rect 530848 363454 531168 363486
rect 530848 363218 530890 363454
rect 531126 363218 531168 363454
rect 530848 363134 531168 363218
rect 530848 362898 530890 363134
rect 531126 362898 531168 363134
rect 530848 362866 531168 362898
rect 561568 363454 561888 363486
rect 561568 363218 561610 363454
rect 561846 363218 561888 363454
rect 561568 363134 561888 363218
rect 561568 362898 561610 363134
rect 561846 362898 561888 363134
rect 561568 362866 561888 362898
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 23968 345454 24288 345486
rect 23968 345218 24010 345454
rect 24246 345218 24288 345454
rect 23968 345134 24288 345218
rect 23968 344898 24010 345134
rect 24246 344898 24288 345134
rect 23968 344866 24288 344898
rect 54688 345454 55008 345486
rect 54688 345218 54730 345454
rect 54966 345218 55008 345454
rect 54688 345134 55008 345218
rect 54688 344898 54730 345134
rect 54966 344898 55008 345134
rect 54688 344866 55008 344898
rect 85408 345454 85728 345486
rect 85408 345218 85450 345454
rect 85686 345218 85728 345454
rect 85408 345134 85728 345218
rect 85408 344898 85450 345134
rect 85686 344898 85728 345134
rect 85408 344866 85728 344898
rect 116128 345454 116448 345486
rect 116128 345218 116170 345454
rect 116406 345218 116448 345454
rect 116128 345134 116448 345218
rect 116128 344898 116170 345134
rect 116406 344898 116448 345134
rect 116128 344866 116448 344898
rect 146848 345454 147168 345486
rect 146848 345218 146890 345454
rect 147126 345218 147168 345454
rect 146848 345134 147168 345218
rect 146848 344898 146890 345134
rect 147126 344898 147168 345134
rect 146848 344866 147168 344898
rect 177568 345454 177888 345486
rect 177568 345218 177610 345454
rect 177846 345218 177888 345454
rect 177568 345134 177888 345218
rect 177568 344898 177610 345134
rect 177846 344898 177888 345134
rect 177568 344866 177888 344898
rect 208288 345454 208608 345486
rect 208288 345218 208330 345454
rect 208566 345218 208608 345454
rect 208288 345134 208608 345218
rect 208288 344898 208330 345134
rect 208566 344898 208608 345134
rect 208288 344866 208608 344898
rect 239008 345454 239328 345486
rect 239008 345218 239050 345454
rect 239286 345218 239328 345454
rect 239008 345134 239328 345218
rect 239008 344898 239050 345134
rect 239286 344898 239328 345134
rect 239008 344866 239328 344898
rect 269728 345454 270048 345486
rect 269728 345218 269770 345454
rect 270006 345218 270048 345454
rect 269728 345134 270048 345218
rect 269728 344898 269770 345134
rect 270006 344898 270048 345134
rect 269728 344866 270048 344898
rect 300448 345454 300768 345486
rect 300448 345218 300490 345454
rect 300726 345218 300768 345454
rect 300448 345134 300768 345218
rect 300448 344898 300490 345134
rect 300726 344898 300768 345134
rect 300448 344866 300768 344898
rect 331168 345454 331488 345486
rect 331168 345218 331210 345454
rect 331446 345218 331488 345454
rect 331168 345134 331488 345218
rect 331168 344898 331210 345134
rect 331446 344898 331488 345134
rect 331168 344866 331488 344898
rect 361888 345454 362208 345486
rect 361888 345218 361930 345454
rect 362166 345218 362208 345454
rect 361888 345134 362208 345218
rect 361888 344898 361930 345134
rect 362166 344898 362208 345134
rect 361888 344866 362208 344898
rect 392608 345454 392928 345486
rect 392608 345218 392650 345454
rect 392886 345218 392928 345454
rect 392608 345134 392928 345218
rect 392608 344898 392650 345134
rect 392886 344898 392928 345134
rect 392608 344866 392928 344898
rect 423328 345454 423648 345486
rect 423328 345218 423370 345454
rect 423606 345218 423648 345454
rect 423328 345134 423648 345218
rect 423328 344898 423370 345134
rect 423606 344898 423648 345134
rect 423328 344866 423648 344898
rect 454048 345454 454368 345486
rect 454048 345218 454090 345454
rect 454326 345218 454368 345454
rect 454048 345134 454368 345218
rect 454048 344898 454090 345134
rect 454326 344898 454368 345134
rect 454048 344866 454368 344898
rect 484768 345454 485088 345486
rect 484768 345218 484810 345454
rect 485046 345218 485088 345454
rect 484768 345134 485088 345218
rect 484768 344898 484810 345134
rect 485046 344898 485088 345134
rect 484768 344866 485088 344898
rect 515488 345454 515808 345486
rect 515488 345218 515530 345454
rect 515766 345218 515808 345454
rect 515488 345134 515808 345218
rect 515488 344898 515530 345134
rect 515766 344898 515808 345134
rect 515488 344866 515808 344898
rect 546208 345454 546528 345486
rect 546208 345218 546250 345454
rect 546486 345218 546528 345454
rect 546208 345134 546528 345218
rect 546208 344898 546250 345134
rect 546486 344898 546528 345134
rect 546208 344866 546528 344898
rect 576928 345454 577248 345486
rect 576928 345218 576970 345454
rect 577206 345218 577248 345454
rect 576928 345134 577248 345218
rect 576928 344898 576970 345134
rect 577206 344898 577248 345134
rect 576928 344866 577248 344898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect 8608 327454 8928 327486
rect 8608 327218 8650 327454
rect 8886 327218 8928 327454
rect 8608 327134 8928 327218
rect 8608 326898 8650 327134
rect 8886 326898 8928 327134
rect 8608 326866 8928 326898
rect 39328 327454 39648 327486
rect 39328 327218 39370 327454
rect 39606 327218 39648 327454
rect 39328 327134 39648 327218
rect 39328 326898 39370 327134
rect 39606 326898 39648 327134
rect 39328 326866 39648 326898
rect 70048 327454 70368 327486
rect 70048 327218 70090 327454
rect 70326 327218 70368 327454
rect 70048 327134 70368 327218
rect 70048 326898 70090 327134
rect 70326 326898 70368 327134
rect 70048 326866 70368 326898
rect 100768 327454 101088 327486
rect 100768 327218 100810 327454
rect 101046 327218 101088 327454
rect 100768 327134 101088 327218
rect 100768 326898 100810 327134
rect 101046 326898 101088 327134
rect 100768 326866 101088 326898
rect 131488 327454 131808 327486
rect 131488 327218 131530 327454
rect 131766 327218 131808 327454
rect 131488 327134 131808 327218
rect 131488 326898 131530 327134
rect 131766 326898 131808 327134
rect 131488 326866 131808 326898
rect 162208 327454 162528 327486
rect 162208 327218 162250 327454
rect 162486 327218 162528 327454
rect 162208 327134 162528 327218
rect 162208 326898 162250 327134
rect 162486 326898 162528 327134
rect 162208 326866 162528 326898
rect 192928 327454 193248 327486
rect 192928 327218 192970 327454
rect 193206 327218 193248 327454
rect 192928 327134 193248 327218
rect 192928 326898 192970 327134
rect 193206 326898 193248 327134
rect 192928 326866 193248 326898
rect 223648 327454 223968 327486
rect 223648 327218 223690 327454
rect 223926 327218 223968 327454
rect 223648 327134 223968 327218
rect 223648 326898 223690 327134
rect 223926 326898 223968 327134
rect 223648 326866 223968 326898
rect 254368 327454 254688 327486
rect 254368 327218 254410 327454
rect 254646 327218 254688 327454
rect 254368 327134 254688 327218
rect 254368 326898 254410 327134
rect 254646 326898 254688 327134
rect 254368 326866 254688 326898
rect 285088 327454 285408 327486
rect 285088 327218 285130 327454
rect 285366 327218 285408 327454
rect 285088 327134 285408 327218
rect 285088 326898 285130 327134
rect 285366 326898 285408 327134
rect 285088 326866 285408 326898
rect 315808 327454 316128 327486
rect 315808 327218 315850 327454
rect 316086 327218 316128 327454
rect 315808 327134 316128 327218
rect 315808 326898 315850 327134
rect 316086 326898 316128 327134
rect 315808 326866 316128 326898
rect 346528 327454 346848 327486
rect 346528 327218 346570 327454
rect 346806 327218 346848 327454
rect 346528 327134 346848 327218
rect 346528 326898 346570 327134
rect 346806 326898 346848 327134
rect 346528 326866 346848 326898
rect 377248 327454 377568 327486
rect 377248 327218 377290 327454
rect 377526 327218 377568 327454
rect 377248 327134 377568 327218
rect 377248 326898 377290 327134
rect 377526 326898 377568 327134
rect 377248 326866 377568 326898
rect 407968 327454 408288 327486
rect 407968 327218 408010 327454
rect 408246 327218 408288 327454
rect 407968 327134 408288 327218
rect 407968 326898 408010 327134
rect 408246 326898 408288 327134
rect 407968 326866 408288 326898
rect 438688 327454 439008 327486
rect 438688 327218 438730 327454
rect 438966 327218 439008 327454
rect 438688 327134 439008 327218
rect 438688 326898 438730 327134
rect 438966 326898 439008 327134
rect 438688 326866 439008 326898
rect 469408 327454 469728 327486
rect 469408 327218 469450 327454
rect 469686 327218 469728 327454
rect 469408 327134 469728 327218
rect 469408 326898 469450 327134
rect 469686 326898 469728 327134
rect 469408 326866 469728 326898
rect 500128 327454 500448 327486
rect 500128 327218 500170 327454
rect 500406 327218 500448 327454
rect 500128 327134 500448 327218
rect 500128 326898 500170 327134
rect 500406 326898 500448 327134
rect 500128 326866 500448 326898
rect 530848 327454 531168 327486
rect 530848 327218 530890 327454
rect 531126 327218 531168 327454
rect 530848 327134 531168 327218
rect 530848 326898 530890 327134
rect 531126 326898 531168 327134
rect 530848 326866 531168 326898
rect 561568 327454 561888 327486
rect 561568 327218 561610 327454
rect 561846 327218 561888 327454
rect 561568 327134 561888 327218
rect 561568 326898 561610 327134
rect 561846 326898 561888 327134
rect 561568 326866 561888 326898
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 23968 309454 24288 309486
rect 23968 309218 24010 309454
rect 24246 309218 24288 309454
rect 23968 309134 24288 309218
rect 23968 308898 24010 309134
rect 24246 308898 24288 309134
rect 23968 308866 24288 308898
rect 54688 309454 55008 309486
rect 54688 309218 54730 309454
rect 54966 309218 55008 309454
rect 54688 309134 55008 309218
rect 54688 308898 54730 309134
rect 54966 308898 55008 309134
rect 54688 308866 55008 308898
rect 85408 309454 85728 309486
rect 85408 309218 85450 309454
rect 85686 309218 85728 309454
rect 85408 309134 85728 309218
rect 85408 308898 85450 309134
rect 85686 308898 85728 309134
rect 85408 308866 85728 308898
rect 116128 309454 116448 309486
rect 116128 309218 116170 309454
rect 116406 309218 116448 309454
rect 116128 309134 116448 309218
rect 116128 308898 116170 309134
rect 116406 308898 116448 309134
rect 116128 308866 116448 308898
rect 146848 309454 147168 309486
rect 146848 309218 146890 309454
rect 147126 309218 147168 309454
rect 146848 309134 147168 309218
rect 146848 308898 146890 309134
rect 147126 308898 147168 309134
rect 146848 308866 147168 308898
rect 177568 309454 177888 309486
rect 177568 309218 177610 309454
rect 177846 309218 177888 309454
rect 177568 309134 177888 309218
rect 177568 308898 177610 309134
rect 177846 308898 177888 309134
rect 177568 308866 177888 308898
rect 208288 309454 208608 309486
rect 208288 309218 208330 309454
rect 208566 309218 208608 309454
rect 208288 309134 208608 309218
rect 208288 308898 208330 309134
rect 208566 308898 208608 309134
rect 208288 308866 208608 308898
rect 239008 309454 239328 309486
rect 239008 309218 239050 309454
rect 239286 309218 239328 309454
rect 239008 309134 239328 309218
rect 239008 308898 239050 309134
rect 239286 308898 239328 309134
rect 239008 308866 239328 308898
rect 269728 309454 270048 309486
rect 269728 309218 269770 309454
rect 270006 309218 270048 309454
rect 269728 309134 270048 309218
rect 269728 308898 269770 309134
rect 270006 308898 270048 309134
rect 269728 308866 270048 308898
rect 300448 309454 300768 309486
rect 300448 309218 300490 309454
rect 300726 309218 300768 309454
rect 300448 309134 300768 309218
rect 300448 308898 300490 309134
rect 300726 308898 300768 309134
rect 300448 308866 300768 308898
rect 331168 309454 331488 309486
rect 331168 309218 331210 309454
rect 331446 309218 331488 309454
rect 331168 309134 331488 309218
rect 331168 308898 331210 309134
rect 331446 308898 331488 309134
rect 331168 308866 331488 308898
rect 361888 309454 362208 309486
rect 361888 309218 361930 309454
rect 362166 309218 362208 309454
rect 361888 309134 362208 309218
rect 361888 308898 361930 309134
rect 362166 308898 362208 309134
rect 361888 308866 362208 308898
rect 392608 309454 392928 309486
rect 392608 309218 392650 309454
rect 392886 309218 392928 309454
rect 392608 309134 392928 309218
rect 392608 308898 392650 309134
rect 392886 308898 392928 309134
rect 392608 308866 392928 308898
rect 423328 309454 423648 309486
rect 423328 309218 423370 309454
rect 423606 309218 423648 309454
rect 423328 309134 423648 309218
rect 423328 308898 423370 309134
rect 423606 308898 423648 309134
rect 423328 308866 423648 308898
rect 454048 309454 454368 309486
rect 454048 309218 454090 309454
rect 454326 309218 454368 309454
rect 454048 309134 454368 309218
rect 454048 308898 454090 309134
rect 454326 308898 454368 309134
rect 454048 308866 454368 308898
rect 484768 309454 485088 309486
rect 484768 309218 484810 309454
rect 485046 309218 485088 309454
rect 484768 309134 485088 309218
rect 484768 308898 484810 309134
rect 485046 308898 485088 309134
rect 484768 308866 485088 308898
rect 515488 309454 515808 309486
rect 515488 309218 515530 309454
rect 515766 309218 515808 309454
rect 515488 309134 515808 309218
rect 515488 308898 515530 309134
rect 515766 308898 515808 309134
rect 515488 308866 515808 308898
rect 546208 309454 546528 309486
rect 546208 309218 546250 309454
rect 546486 309218 546528 309454
rect 546208 309134 546528 309218
rect 546208 308898 546250 309134
rect 546486 308898 546528 309134
rect 546208 308866 546528 308898
rect 576928 309454 577248 309486
rect 576928 309218 576970 309454
rect 577206 309218 577248 309454
rect 576928 309134 577248 309218
rect 576928 308898 576970 309134
rect 577206 308898 577248 309134
rect 576928 308866 577248 308898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect 8608 291454 8928 291486
rect 8608 291218 8650 291454
rect 8886 291218 8928 291454
rect 8608 291134 8928 291218
rect 8608 290898 8650 291134
rect 8886 290898 8928 291134
rect 8608 290866 8928 290898
rect 39328 291454 39648 291486
rect 39328 291218 39370 291454
rect 39606 291218 39648 291454
rect 39328 291134 39648 291218
rect 39328 290898 39370 291134
rect 39606 290898 39648 291134
rect 39328 290866 39648 290898
rect 70048 291454 70368 291486
rect 70048 291218 70090 291454
rect 70326 291218 70368 291454
rect 70048 291134 70368 291218
rect 70048 290898 70090 291134
rect 70326 290898 70368 291134
rect 70048 290866 70368 290898
rect 100768 291454 101088 291486
rect 100768 291218 100810 291454
rect 101046 291218 101088 291454
rect 100768 291134 101088 291218
rect 100768 290898 100810 291134
rect 101046 290898 101088 291134
rect 100768 290866 101088 290898
rect 131488 291454 131808 291486
rect 131488 291218 131530 291454
rect 131766 291218 131808 291454
rect 131488 291134 131808 291218
rect 131488 290898 131530 291134
rect 131766 290898 131808 291134
rect 131488 290866 131808 290898
rect 162208 291454 162528 291486
rect 162208 291218 162250 291454
rect 162486 291218 162528 291454
rect 162208 291134 162528 291218
rect 162208 290898 162250 291134
rect 162486 290898 162528 291134
rect 162208 290866 162528 290898
rect 192928 291454 193248 291486
rect 192928 291218 192970 291454
rect 193206 291218 193248 291454
rect 192928 291134 193248 291218
rect 192928 290898 192970 291134
rect 193206 290898 193248 291134
rect 192928 290866 193248 290898
rect 223648 291454 223968 291486
rect 223648 291218 223690 291454
rect 223926 291218 223968 291454
rect 223648 291134 223968 291218
rect 223648 290898 223690 291134
rect 223926 290898 223968 291134
rect 223648 290866 223968 290898
rect 254368 291454 254688 291486
rect 254368 291218 254410 291454
rect 254646 291218 254688 291454
rect 254368 291134 254688 291218
rect 254368 290898 254410 291134
rect 254646 290898 254688 291134
rect 254368 290866 254688 290898
rect 285088 291454 285408 291486
rect 285088 291218 285130 291454
rect 285366 291218 285408 291454
rect 285088 291134 285408 291218
rect 285088 290898 285130 291134
rect 285366 290898 285408 291134
rect 285088 290866 285408 290898
rect 315808 291454 316128 291486
rect 315808 291218 315850 291454
rect 316086 291218 316128 291454
rect 315808 291134 316128 291218
rect 315808 290898 315850 291134
rect 316086 290898 316128 291134
rect 315808 290866 316128 290898
rect 346528 291454 346848 291486
rect 346528 291218 346570 291454
rect 346806 291218 346848 291454
rect 346528 291134 346848 291218
rect 346528 290898 346570 291134
rect 346806 290898 346848 291134
rect 346528 290866 346848 290898
rect 377248 291454 377568 291486
rect 377248 291218 377290 291454
rect 377526 291218 377568 291454
rect 377248 291134 377568 291218
rect 377248 290898 377290 291134
rect 377526 290898 377568 291134
rect 377248 290866 377568 290898
rect 407968 291454 408288 291486
rect 407968 291218 408010 291454
rect 408246 291218 408288 291454
rect 407968 291134 408288 291218
rect 407968 290898 408010 291134
rect 408246 290898 408288 291134
rect 407968 290866 408288 290898
rect 438688 291454 439008 291486
rect 438688 291218 438730 291454
rect 438966 291218 439008 291454
rect 438688 291134 439008 291218
rect 438688 290898 438730 291134
rect 438966 290898 439008 291134
rect 438688 290866 439008 290898
rect 469408 291454 469728 291486
rect 469408 291218 469450 291454
rect 469686 291218 469728 291454
rect 469408 291134 469728 291218
rect 469408 290898 469450 291134
rect 469686 290898 469728 291134
rect 469408 290866 469728 290898
rect 500128 291454 500448 291486
rect 500128 291218 500170 291454
rect 500406 291218 500448 291454
rect 500128 291134 500448 291218
rect 500128 290898 500170 291134
rect 500406 290898 500448 291134
rect 500128 290866 500448 290898
rect 530848 291454 531168 291486
rect 530848 291218 530890 291454
rect 531126 291218 531168 291454
rect 530848 291134 531168 291218
rect 530848 290898 530890 291134
rect 531126 290898 531168 291134
rect 530848 290866 531168 290898
rect 561568 291454 561888 291486
rect 561568 291218 561610 291454
rect 561846 291218 561888 291454
rect 561568 291134 561888 291218
rect 561568 290898 561610 291134
rect 561846 290898 561888 291134
rect 561568 290866 561888 290898
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 23968 273454 24288 273486
rect 23968 273218 24010 273454
rect 24246 273218 24288 273454
rect 23968 273134 24288 273218
rect 23968 272898 24010 273134
rect 24246 272898 24288 273134
rect 23968 272866 24288 272898
rect 54688 273454 55008 273486
rect 54688 273218 54730 273454
rect 54966 273218 55008 273454
rect 54688 273134 55008 273218
rect 54688 272898 54730 273134
rect 54966 272898 55008 273134
rect 54688 272866 55008 272898
rect 85408 273454 85728 273486
rect 85408 273218 85450 273454
rect 85686 273218 85728 273454
rect 85408 273134 85728 273218
rect 85408 272898 85450 273134
rect 85686 272898 85728 273134
rect 85408 272866 85728 272898
rect 116128 273454 116448 273486
rect 116128 273218 116170 273454
rect 116406 273218 116448 273454
rect 116128 273134 116448 273218
rect 116128 272898 116170 273134
rect 116406 272898 116448 273134
rect 116128 272866 116448 272898
rect 146848 273454 147168 273486
rect 146848 273218 146890 273454
rect 147126 273218 147168 273454
rect 146848 273134 147168 273218
rect 146848 272898 146890 273134
rect 147126 272898 147168 273134
rect 146848 272866 147168 272898
rect 177568 273454 177888 273486
rect 177568 273218 177610 273454
rect 177846 273218 177888 273454
rect 177568 273134 177888 273218
rect 177568 272898 177610 273134
rect 177846 272898 177888 273134
rect 177568 272866 177888 272898
rect 208288 273454 208608 273486
rect 208288 273218 208330 273454
rect 208566 273218 208608 273454
rect 208288 273134 208608 273218
rect 208288 272898 208330 273134
rect 208566 272898 208608 273134
rect 208288 272866 208608 272898
rect 239008 273454 239328 273486
rect 239008 273218 239050 273454
rect 239286 273218 239328 273454
rect 239008 273134 239328 273218
rect 239008 272898 239050 273134
rect 239286 272898 239328 273134
rect 239008 272866 239328 272898
rect 269728 273454 270048 273486
rect 269728 273218 269770 273454
rect 270006 273218 270048 273454
rect 269728 273134 270048 273218
rect 269728 272898 269770 273134
rect 270006 272898 270048 273134
rect 269728 272866 270048 272898
rect 300448 273454 300768 273486
rect 300448 273218 300490 273454
rect 300726 273218 300768 273454
rect 300448 273134 300768 273218
rect 300448 272898 300490 273134
rect 300726 272898 300768 273134
rect 300448 272866 300768 272898
rect 331168 273454 331488 273486
rect 331168 273218 331210 273454
rect 331446 273218 331488 273454
rect 331168 273134 331488 273218
rect 331168 272898 331210 273134
rect 331446 272898 331488 273134
rect 331168 272866 331488 272898
rect 361888 273454 362208 273486
rect 361888 273218 361930 273454
rect 362166 273218 362208 273454
rect 361888 273134 362208 273218
rect 361888 272898 361930 273134
rect 362166 272898 362208 273134
rect 361888 272866 362208 272898
rect 392608 273454 392928 273486
rect 392608 273218 392650 273454
rect 392886 273218 392928 273454
rect 392608 273134 392928 273218
rect 392608 272898 392650 273134
rect 392886 272898 392928 273134
rect 392608 272866 392928 272898
rect 423328 273454 423648 273486
rect 423328 273218 423370 273454
rect 423606 273218 423648 273454
rect 423328 273134 423648 273218
rect 423328 272898 423370 273134
rect 423606 272898 423648 273134
rect 423328 272866 423648 272898
rect 454048 273454 454368 273486
rect 454048 273218 454090 273454
rect 454326 273218 454368 273454
rect 454048 273134 454368 273218
rect 454048 272898 454090 273134
rect 454326 272898 454368 273134
rect 454048 272866 454368 272898
rect 484768 273454 485088 273486
rect 484768 273218 484810 273454
rect 485046 273218 485088 273454
rect 484768 273134 485088 273218
rect 484768 272898 484810 273134
rect 485046 272898 485088 273134
rect 484768 272866 485088 272898
rect 515488 273454 515808 273486
rect 515488 273218 515530 273454
rect 515766 273218 515808 273454
rect 515488 273134 515808 273218
rect 515488 272898 515530 273134
rect 515766 272898 515808 273134
rect 515488 272866 515808 272898
rect 546208 273454 546528 273486
rect 546208 273218 546250 273454
rect 546486 273218 546528 273454
rect 546208 273134 546528 273218
rect 546208 272898 546250 273134
rect 546486 272898 546528 273134
rect 546208 272866 546528 272898
rect 576928 273454 577248 273486
rect 576928 273218 576970 273454
rect 577206 273218 577248 273454
rect 576928 273134 577248 273218
rect 576928 272898 576970 273134
rect 577206 272898 577248 273134
rect 576928 272866 577248 272898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect 8608 255454 8928 255486
rect 8608 255218 8650 255454
rect 8886 255218 8928 255454
rect 8608 255134 8928 255218
rect 8608 254898 8650 255134
rect 8886 254898 8928 255134
rect 8608 254866 8928 254898
rect 39328 255454 39648 255486
rect 39328 255218 39370 255454
rect 39606 255218 39648 255454
rect 39328 255134 39648 255218
rect 39328 254898 39370 255134
rect 39606 254898 39648 255134
rect 39328 254866 39648 254898
rect 70048 255454 70368 255486
rect 70048 255218 70090 255454
rect 70326 255218 70368 255454
rect 70048 255134 70368 255218
rect 70048 254898 70090 255134
rect 70326 254898 70368 255134
rect 70048 254866 70368 254898
rect 100768 255454 101088 255486
rect 100768 255218 100810 255454
rect 101046 255218 101088 255454
rect 100768 255134 101088 255218
rect 100768 254898 100810 255134
rect 101046 254898 101088 255134
rect 100768 254866 101088 254898
rect 131488 255454 131808 255486
rect 131488 255218 131530 255454
rect 131766 255218 131808 255454
rect 131488 255134 131808 255218
rect 131488 254898 131530 255134
rect 131766 254898 131808 255134
rect 131488 254866 131808 254898
rect 162208 255454 162528 255486
rect 162208 255218 162250 255454
rect 162486 255218 162528 255454
rect 162208 255134 162528 255218
rect 162208 254898 162250 255134
rect 162486 254898 162528 255134
rect 162208 254866 162528 254898
rect 192928 255454 193248 255486
rect 192928 255218 192970 255454
rect 193206 255218 193248 255454
rect 192928 255134 193248 255218
rect 192928 254898 192970 255134
rect 193206 254898 193248 255134
rect 192928 254866 193248 254898
rect 223648 255454 223968 255486
rect 223648 255218 223690 255454
rect 223926 255218 223968 255454
rect 223648 255134 223968 255218
rect 223648 254898 223690 255134
rect 223926 254898 223968 255134
rect 223648 254866 223968 254898
rect 254368 255454 254688 255486
rect 254368 255218 254410 255454
rect 254646 255218 254688 255454
rect 254368 255134 254688 255218
rect 254368 254898 254410 255134
rect 254646 254898 254688 255134
rect 254368 254866 254688 254898
rect 285088 255454 285408 255486
rect 285088 255218 285130 255454
rect 285366 255218 285408 255454
rect 285088 255134 285408 255218
rect 285088 254898 285130 255134
rect 285366 254898 285408 255134
rect 285088 254866 285408 254898
rect 315808 255454 316128 255486
rect 315808 255218 315850 255454
rect 316086 255218 316128 255454
rect 315808 255134 316128 255218
rect 315808 254898 315850 255134
rect 316086 254898 316128 255134
rect 315808 254866 316128 254898
rect 346528 255454 346848 255486
rect 346528 255218 346570 255454
rect 346806 255218 346848 255454
rect 346528 255134 346848 255218
rect 346528 254898 346570 255134
rect 346806 254898 346848 255134
rect 346528 254866 346848 254898
rect 377248 255454 377568 255486
rect 377248 255218 377290 255454
rect 377526 255218 377568 255454
rect 377248 255134 377568 255218
rect 377248 254898 377290 255134
rect 377526 254898 377568 255134
rect 377248 254866 377568 254898
rect 407968 255454 408288 255486
rect 407968 255218 408010 255454
rect 408246 255218 408288 255454
rect 407968 255134 408288 255218
rect 407968 254898 408010 255134
rect 408246 254898 408288 255134
rect 407968 254866 408288 254898
rect 438688 255454 439008 255486
rect 438688 255218 438730 255454
rect 438966 255218 439008 255454
rect 438688 255134 439008 255218
rect 438688 254898 438730 255134
rect 438966 254898 439008 255134
rect 438688 254866 439008 254898
rect 469408 255454 469728 255486
rect 469408 255218 469450 255454
rect 469686 255218 469728 255454
rect 469408 255134 469728 255218
rect 469408 254898 469450 255134
rect 469686 254898 469728 255134
rect 469408 254866 469728 254898
rect 500128 255454 500448 255486
rect 500128 255218 500170 255454
rect 500406 255218 500448 255454
rect 500128 255134 500448 255218
rect 500128 254898 500170 255134
rect 500406 254898 500448 255134
rect 500128 254866 500448 254898
rect 530848 255454 531168 255486
rect 530848 255218 530890 255454
rect 531126 255218 531168 255454
rect 530848 255134 531168 255218
rect 530848 254898 530890 255134
rect 531126 254898 531168 255134
rect 530848 254866 531168 254898
rect 561568 255454 561888 255486
rect 561568 255218 561610 255454
rect 561846 255218 561888 255454
rect 561568 255134 561888 255218
rect 561568 254898 561610 255134
rect 561846 254898 561888 255134
rect 561568 254866 561888 254898
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 23968 237454 24288 237486
rect 23968 237218 24010 237454
rect 24246 237218 24288 237454
rect 23968 237134 24288 237218
rect 23968 236898 24010 237134
rect 24246 236898 24288 237134
rect 23968 236866 24288 236898
rect 54688 237454 55008 237486
rect 54688 237218 54730 237454
rect 54966 237218 55008 237454
rect 54688 237134 55008 237218
rect 54688 236898 54730 237134
rect 54966 236898 55008 237134
rect 54688 236866 55008 236898
rect 85408 237454 85728 237486
rect 85408 237218 85450 237454
rect 85686 237218 85728 237454
rect 85408 237134 85728 237218
rect 85408 236898 85450 237134
rect 85686 236898 85728 237134
rect 85408 236866 85728 236898
rect 116128 237454 116448 237486
rect 116128 237218 116170 237454
rect 116406 237218 116448 237454
rect 116128 237134 116448 237218
rect 116128 236898 116170 237134
rect 116406 236898 116448 237134
rect 116128 236866 116448 236898
rect 146848 237454 147168 237486
rect 146848 237218 146890 237454
rect 147126 237218 147168 237454
rect 146848 237134 147168 237218
rect 146848 236898 146890 237134
rect 147126 236898 147168 237134
rect 146848 236866 147168 236898
rect 177568 237454 177888 237486
rect 177568 237218 177610 237454
rect 177846 237218 177888 237454
rect 177568 237134 177888 237218
rect 177568 236898 177610 237134
rect 177846 236898 177888 237134
rect 177568 236866 177888 236898
rect 208288 237454 208608 237486
rect 208288 237218 208330 237454
rect 208566 237218 208608 237454
rect 208288 237134 208608 237218
rect 208288 236898 208330 237134
rect 208566 236898 208608 237134
rect 208288 236866 208608 236898
rect 239008 237454 239328 237486
rect 239008 237218 239050 237454
rect 239286 237218 239328 237454
rect 239008 237134 239328 237218
rect 239008 236898 239050 237134
rect 239286 236898 239328 237134
rect 239008 236866 239328 236898
rect 269728 237454 270048 237486
rect 269728 237218 269770 237454
rect 270006 237218 270048 237454
rect 269728 237134 270048 237218
rect 269728 236898 269770 237134
rect 270006 236898 270048 237134
rect 269728 236866 270048 236898
rect 300448 237454 300768 237486
rect 300448 237218 300490 237454
rect 300726 237218 300768 237454
rect 300448 237134 300768 237218
rect 300448 236898 300490 237134
rect 300726 236898 300768 237134
rect 300448 236866 300768 236898
rect 331168 237454 331488 237486
rect 331168 237218 331210 237454
rect 331446 237218 331488 237454
rect 331168 237134 331488 237218
rect 331168 236898 331210 237134
rect 331446 236898 331488 237134
rect 331168 236866 331488 236898
rect 361888 237454 362208 237486
rect 361888 237218 361930 237454
rect 362166 237218 362208 237454
rect 361888 237134 362208 237218
rect 361888 236898 361930 237134
rect 362166 236898 362208 237134
rect 361888 236866 362208 236898
rect 392608 237454 392928 237486
rect 392608 237218 392650 237454
rect 392886 237218 392928 237454
rect 392608 237134 392928 237218
rect 392608 236898 392650 237134
rect 392886 236898 392928 237134
rect 392608 236866 392928 236898
rect 423328 237454 423648 237486
rect 423328 237218 423370 237454
rect 423606 237218 423648 237454
rect 423328 237134 423648 237218
rect 423328 236898 423370 237134
rect 423606 236898 423648 237134
rect 423328 236866 423648 236898
rect 454048 237454 454368 237486
rect 454048 237218 454090 237454
rect 454326 237218 454368 237454
rect 454048 237134 454368 237218
rect 454048 236898 454090 237134
rect 454326 236898 454368 237134
rect 454048 236866 454368 236898
rect 484768 237454 485088 237486
rect 484768 237218 484810 237454
rect 485046 237218 485088 237454
rect 484768 237134 485088 237218
rect 484768 236898 484810 237134
rect 485046 236898 485088 237134
rect 484768 236866 485088 236898
rect 515488 237454 515808 237486
rect 515488 237218 515530 237454
rect 515766 237218 515808 237454
rect 515488 237134 515808 237218
rect 515488 236898 515530 237134
rect 515766 236898 515808 237134
rect 515488 236866 515808 236898
rect 546208 237454 546528 237486
rect 546208 237218 546250 237454
rect 546486 237218 546528 237454
rect 546208 237134 546528 237218
rect 546208 236898 546250 237134
rect 546486 236898 546528 237134
rect 546208 236866 546528 236898
rect 576928 237454 577248 237486
rect 576928 237218 576970 237454
rect 577206 237218 577248 237454
rect 576928 237134 577248 237218
rect 576928 236898 576970 237134
rect 577206 236898 577248 237134
rect 576928 236866 577248 236898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect 8608 219454 8928 219486
rect 8608 219218 8650 219454
rect 8886 219218 8928 219454
rect 8608 219134 8928 219218
rect 8608 218898 8650 219134
rect 8886 218898 8928 219134
rect 8608 218866 8928 218898
rect 39328 219454 39648 219486
rect 39328 219218 39370 219454
rect 39606 219218 39648 219454
rect 39328 219134 39648 219218
rect 39328 218898 39370 219134
rect 39606 218898 39648 219134
rect 39328 218866 39648 218898
rect 70048 219454 70368 219486
rect 70048 219218 70090 219454
rect 70326 219218 70368 219454
rect 70048 219134 70368 219218
rect 70048 218898 70090 219134
rect 70326 218898 70368 219134
rect 70048 218866 70368 218898
rect 100768 219454 101088 219486
rect 100768 219218 100810 219454
rect 101046 219218 101088 219454
rect 100768 219134 101088 219218
rect 100768 218898 100810 219134
rect 101046 218898 101088 219134
rect 100768 218866 101088 218898
rect 131488 219454 131808 219486
rect 131488 219218 131530 219454
rect 131766 219218 131808 219454
rect 131488 219134 131808 219218
rect 131488 218898 131530 219134
rect 131766 218898 131808 219134
rect 131488 218866 131808 218898
rect 162208 219454 162528 219486
rect 162208 219218 162250 219454
rect 162486 219218 162528 219454
rect 162208 219134 162528 219218
rect 162208 218898 162250 219134
rect 162486 218898 162528 219134
rect 162208 218866 162528 218898
rect 192928 219454 193248 219486
rect 192928 219218 192970 219454
rect 193206 219218 193248 219454
rect 192928 219134 193248 219218
rect 192928 218898 192970 219134
rect 193206 218898 193248 219134
rect 192928 218866 193248 218898
rect 223648 219454 223968 219486
rect 223648 219218 223690 219454
rect 223926 219218 223968 219454
rect 223648 219134 223968 219218
rect 223648 218898 223690 219134
rect 223926 218898 223968 219134
rect 223648 218866 223968 218898
rect 254368 219454 254688 219486
rect 254368 219218 254410 219454
rect 254646 219218 254688 219454
rect 254368 219134 254688 219218
rect 254368 218898 254410 219134
rect 254646 218898 254688 219134
rect 254368 218866 254688 218898
rect 285088 219454 285408 219486
rect 285088 219218 285130 219454
rect 285366 219218 285408 219454
rect 285088 219134 285408 219218
rect 285088 218898 285130 219134
rect 285366 218898 285408 219134
rect 285088 218866 285408 218898
rect 315808 219454 316128 219486
rect 315808 219218 315850 219454
rect 316086 219218 316128 219454
rect 315808 219134 316128 219218
rect 315808 218898 315850 219134
rect 316086 218898 316128 219134
rect 315808 218866 316128 218898
rect 346528 219454 346848 219486
rect 346528 219218 346570 219454
rect 346806 219218 346848 219454
rect 346528 219134 346848 219218
rect 346528 218898 346570 219134
rect 346806 218898 346848 219134
rect 346528 218866 346848 218898
rect 377248 219454 377568 219486
rect 377248 219218 377290 219454
rect 377526 219218 377568 219454
rect 377248 219134 377568 219218
rect 377248 218898 377290 219134
rect 377526 218898 377568 219134
rect 377248 218866 377568 218898
rect 407968 219454 408288 219486
rect 407968 219218 408010 219454
rect 408246 219218 408288 219454
rect 407968 219134 408288 219218
rect 407968 218898 408010 219134
rect 408246 218898 408288 219134
rect 407968 218866 408288 218898
rect 438688 219454 439008 219486
rect 438688 219218 438730 219454
rect 438966 219218 439008 219454
rect 438688 219134 439008 219218
rect 438688 218898 438730 219134
rect 438966 218898 439008 219134
rect 438688 218866 439008 218898
rect 469408 219454 469728 219486
rect 469408 219218 469450 219454
rect 469686 219218 469728 219454
rect 469408 219134 469728 219218
rect 469408 218898 469450 219134
rect 469686 218898 469728 219134
rect 469408 218866 469728 218898
rect 500128 219454 500448 219486
rect 500128 219218 500170 219454
rect 500406 219218 500448 219454
rect 500128 219134 500448 219218
rect 500128 218898 500170 219134
rect 500406 218898 500448 219134
rect 500128 218866 500448 218898
rect 530848 219454 531168 219486
rect 530848 219218 530890 219454
rect 531126 219218 531168 219454
rect 530848 219134 531168 219218
rect 530848 218898 530890 219134
rect 531126 218898 531168 219134
rect 530848 218866 531168 218898
rect 561568 219454 561888 219486
rect 561568 219218 561610 219454
rect 561846 219218 561888 219454
rect 561568 219134 561888 219218
rect 561568 218898 561610 219134
rect 561846 218898 561888 219134
rect 561568 218866 561888 218898
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 23968 201454 24288 201486
rect 23968 201218 24010 201454
rect 24246 201218 24288 201454
rect 23968 201134 24288 201218
rect 23968 200898 24010 201134
rect 24246 200898 24288 201134
rect 23968 200866 24288 200898
rect 54688 201454 55008 201486
rect 54688 201218 54730 201454
rect 54966 201218 55008 201454
rect 54688 201134 55008 201218
rect 54688 200898 54730 201134
rect 54966 200898 55008 201134
rect 54688 200866 55008 200898
rect 85408 201454 85728 201486
rect 85408 201218 85450 201454
rect 85686 201218 85728 201454
rect 85408 201134 85728 201218
rect 85408 200898 85450 201134
rect 85686 200898 85728 201134
rect 85408 200866 85728 200898
rect 116128 201454 116448 201486
rect 116128 201218 116170 201454
rect 116406 201218 116448 201454
rect 116128 201134 116448 201218
rect 116128 200898 116170 201134
rect 116406 200898 116448 201134
rect 116128 200866 116448 200898
rect 146848 201454 147168 201486
rect 146848 201218 146890 201454
rect 147126 201218 147168 201454
rect 146848 201134 147168 201218
rect 146848 200898 146890 201134
rect 147126 200898 147168 201134
rect 146848 200866 147168 200898
rect 177568 201454 177888 201486
rect 177568 201218 177610 201454
rect 177846 201218 177888 201454
rect 177568 201134 177888 201218
rect 177568 200898 177610 201134
rect 177846 200898 177888 201134
rect 177568 200866 177888 200898
rect 208288 201454 208608 201486
rect 208288 201218 208330 201454
rect 208566 201218 208608 201454
rect 208288 201134 208608 201218
rect 208288 200898 208330 201134
rect 208566 200898 208608 201134
rect 208288 200866 208608 200898
rect 239008 201454 239328 201486
rect 239008 201218 239050 201454
rect 239286 201218 239328 201454
rect 239008 201134 239328 201218
rect 239008 200898 239050 201134
rect 239286 200898 239328 201134
rect 239008 200866 239328 200898
rect 269728 201454 270048 201486
rect 269728 201218 269770 201454
rect 270006 201218 270048 201454
rect 269728 201134 270048 201218
rect 269728 200898 269770 201134
rect 270006 200898 270048 201134
rect 269728 200866 270048 200898
rect 300448 201454 300768 201486
rect 300448 201218 300490 201454
rect 300726 201218 300768 201454
rect 300448 201134 300768 201218
rect 300448 200898 300490 201134
rect 300726 200898 300768 201134
rect 300448 200866 300768 200898
rect 331168 201454 331488 201486
rect 331168 201218 331210 201454
rect 331446 201218 331488 201454
rect 331168 201134 331488 201218
rect 331168 200898 331210 201134
rect 331446 200898 331488 201134
rect 331168 200866 331488 200898
rect 361888 201454 362208 201486
rect 361888 201218 361930 201454
rect 362166 201218 362208 201454
rect 361888 201134 362208 201218
rect 361888 200898 361930 201134
rect 362166 200898 362208 201134
rect 361888 200866 362208 200898
rect 392608 201454 392928 201486
rect 392608 201218 392650 201454
rect 392886 201218 392928 201454
rect 392608 201134 392928 201218
rect 392608 200898 392650 201134
rect 392886 200898 392928 201134
rect 392608 200866 392928 200898
rect 423328 201454 423648 201486
rect 423328 201218 423370 201454
rect 423606 201218 423648 201454
rect 423328 201134 423648 201218
rect 423328 200898 423370 201134
rect 423606 200898 423648 201134
rect 423328 200866 423648 200898
rect 454048 201454 454368 201486
rect 454048 201218 454090 201454
rect 454326 201218 454368 201454
rect 454048 201134 454368 201218
rect 454048 200898 454090 201134
rect 454326 200898 454368 201134
rect 454048 200866 454368 200898
rect 484768 201454 485088 201486
rect 484768 201218 484810 201454
rect 485046 201218 485088 201454
rect 484768 201134 485088 201218
rect 484768 200898 484810 201134
rect 485046 200898 485088 201134
rect 484768 200866 485088 200898
rect 515488 201454 515808 201486
rect 515488 201218 515530 201454
rect 515766 201218 515808 201454
rect 515488 201134 515808 201218
rect 515488 200898 515530 201134
rect 515766 200898 515808 201134
rect 515488 200866 515808 200898
rect 546208 201454 546528 201486
rect 546208 201218 546250 201454
rect 546486 201218 546528 201454
rect 546208 201134 546528 201218
rect 546208 200898 546250 201134
rect 546486 200898 546528 201134
rect 546208 200866 546528 200898
rect 576928 201454 577248 201486
rect 576928 201218 576970 201454
rect 577206 201218 577248 201454
rect 576928 201134 577248 201218
rect 576928 200898 576970 201134
rect 577206 200898 577248 201134
rect 576928 200866 577248 200898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect 8608 183454 8928 183486
rect 8608 183218 8650 183454
rect 8886 183218 8928 183454
rect 8608 183134 8928 183218
rect 8608 182898 8650 183134
rect 8886 182898 8928 183134
rect 8608 182866 8928 182898
rect 39328 183454 39648 183486
rect 39328 183218 39370 183454
rect 39606 183218 39648 183454
rect 39328 183134 39648 183218
rect 39328 182898 39370 183134
rect 39606 182898 39648 183134
rect 39328 182866 39648 182898
rect 70048 183454 70368 183486
rect 70048 183218 70090 183454
rect 70326 183218 70368 183454
rect 70048 183134 70368 183218
rect 70048 182898 70090 183134
rect 70326 182898 70368 183134
rect 70048 182866 70368 182898
rect 100768 183454 101088 183486
rect 100768 183218 100810 183454
rect 101046 183218 101088 183454
rect 100768 183134 101088 183218
rect 100768 182898 100810 183134
rect 101046 182898 101088 183134
rect 100768 182866 101088 182898
rect 131488 183454 131808 183486
rect 131488 183218 131530 183454
rect 131766 183218 131808 183454
rect 131488 183134 131808 183218
rect 131488 182898 131530 183134
rect 131766 182898 131808 183134
rect 131488 182866 131808 182898
rect 162208 183454 162528 183486
rect 162208 183218 162250 183454
rect 162486 183218 162528 183454
rect 162208 183134 162528 183218
rect 162208 182898 162250 183134
rect 162486 182898 162528 183134
rect 162208 182866 162528 182898
rect 192928 183454 193248 183486
rect 192928 183218 192970 183454
rect 193206 183218 193248 183454
rect 192928 183134 193248 183218
rect 192928 182898 192970 183134
rect 193206 182898 193248 183134
rect 192928 182866 193248 182898
rect 223648 183454 223968 183486
rect 223648 183218 223690 183454
rect 223926 183218 223968 183454
rect 223648 183134 223968 183218
rect 223648 182898 223690 183134
rect 223926 182898 223968 183134
rect 223648 182866 223968 182898
rect 254368 183454 254688 183486
rect 254368 183218 254410 183454
rect 254646 183218 254688 183454
rect 254368 183134 254688 183218
rect 254368 182898 254410 183134
rect 254646 182898 254688 183134
rect 254368 182866 254688 182898
rect 285088 183454 285408 183486
rect 285088 183218 285130 183454
rect 285366 183218 285408 183454
rect 285088 183134 285408 183218
rect 285088 182898 285130 183134
rect 285366 182898 285408 183134
rect 285088 182866 285408 182898
rect 315808 183454 316128 183486
rect 315808 183218 315850 183454
rect 316086 183218 316128 183454
rect 315808 183134 316128 183218
rect 315808 182898 315850 183134
rect 316086 182898 316128 183134
rect 315808 182866 316128 182898
rect 346528 183454 346848 183486
rect 346528 183218 346570 183454
rect 346806 183218 346848 183454
rect 346528 183134 346848 183218
rect 346528 182898 346570 183134
rect 346806 182898 346848 183134
rect 346528 182866 346848 182898
rect 377248 183454 377568 183486
rect 377248 183218 377290 183454
rect 377526 183218 377568 183454
rect 377248 183134 377568 183218
rect 377248 182898 377290 183134
rect 377526 182898 377568 183134
rect 377248 182866 377568 182898
rect 407968 183454 408288 183486
rect 407968 183218 408010 183454
rect 408246 183218 408288 183454
rect 407968 183134 408288 183218
rect 407968 182898 408010 183134
rect 408246 182898 408288 183134
rect 407968 182866 408288 182898
rect 438688 183454 439008 183486
rect 438688 183218 438730 183454
rect 438966 183218 439008 183454
rect 438688 183134 439008 183218
rect 438688 182898 438730 183134
rect 438966 182898 439008 183134
rect 438688 182866 439008 182898
rect 469408 183454 469728 183486
rect 469408 183218 469450 183454
rect 469686 183218 469728 183454
rect 469408 183134 469728 183218
rect 469408 182898 469450 183134
rect 469686 182898 469728 183134
rect 469408 182866 469728 182898
rect 500128 183454 500448 183486
rect 500128 183218 500170 183454
rect 500406 183218 500448 183454
rect 500128 183134 500448 183218
rect 500128 182898 500170 183134
rect 500406 182898 500448 183134
rect 500128 182866 500448 182898
rect 530848 183454 531168 183486
rect 530848 183218 530890 183454
rect 531126 183218 531168 183454
rect 530848 183134 531168 183218
rect 530848 182898 530890 183134
rect 531126 182898 531168 183134
rect 530848 182866 531168 182898
rect 561568 183454 561888 183486
rect 561568 183218 561610 183454
rect 561846 183218 561888 183454
rect 561568 183134 561888 183218
rect 561568 182898 561610 183134
rect 561846 182898 561888 183134
rect 561568 182866 561888 182898
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 23968 165454 24288 165486
rect 23968 165218 24010 165454
rect 24246 165218 24288 165454
rect 23968 165134 24288 165218
rect 23968 164898 24010 165134
rect 24246 164898 24288 165134
rect 23968 164866 24288 164898
rect 54688 165454 55008 165486
rect 54688 165218 54730 165454
rect 54966 165218 55008 165454
rect 54688 165134 55008 165218
rect 54688 164898 54730 165134
rect 54966 164898 55008 165134
rect 54688 164866 55008 164898
rect 85408 165454 85728 165486
rect 85408 165218 85450 165454
rect 85686 165218 85728 165454
rect 85408 165134 85728 165218
rect 85408 164898 85450 165134
rect 85686 164898 85728 165134
rect 85408 164866 85728 164898
rect 116128 165454 116448 165486
rect 116128 165218 116170 165454
rect 116406 165218 116448 165454
rect 116128 165134 116448 165218
rect 116128 164898 116170 165134
rect 116406 164898 116448 165134
rect 116128 164866 116448 164898
rect 146848 165454 147168 165486
rect 146848 165218 146890 165454
rect 147126 165218 147168 165454
rect 146848 165134 147168 165218
rect 146848 164898 146890 165134
rect 147126 164898 147168 165134
rect 146848 164866 147168 164898
rect 177568 165454 177888 165486
rect 177568 165218 177610 165454
rect 177846 165218 177888 165454
rect 177568 165134 177888 165218
rect 177568 164898 177610 165134
rect 177846 164898 177888 165134
rect 177568 164866 177888 164898
rect 208288 165454 208608 165486
rect 208288 165218 208330 165454
rect 208566 165218 208608 165454
rect 208288 165134 208608 165218
rect 208288 164898 208330 165134
rect 208566 164898 208608 165134
rect 208288 164866 208608 164898
rect 239008 165454 239328 165486
rect 239008 165218 239050 165454
rect 239286 165218 239328 165454
rect 239008 165134 239328 165218
rect 239008 164898 239050 165134
rect 239286 164898 239328 165134
rect 239008 164866 239328 164898
rect 269728 165454 270048 165486
rect 269728 165218 269770 165454
rect 270006 165218 270048 165454
rect 269728 165134 270048 165218
rect 269728 164898 269770 165134
rect 270006 164898 270048 165134
rect 269728 164866 270048 164898
rect 300448 165454 300768 165486
rect 300448 165218 300490 165454
rect 300726 165218 300768 165454
rect 300448 165134 300768 165218
rect 300448 164898 300490 165134
rect 300726 164898 300768 165134
rect 300448 164866 300768 164898
rect 331168 165454 331488 165486
rect 331168 165218 331210 165454
rect 331446 165218 331488 165454
rect 331168 165134 331488 165218
rect 331168 164898 331210 165134
rect 331446 164898 331488 165134
rect 331168 164866 331488 164898
rect 361888 165454 362208 165486
rect 361888 165218 361930 165454
rect 362166 165218 362208 165454
rect 361888 165134 362208 165218
rect 361888 164898 361930 165134
rect 362166 164898 362208 165134
rect 361888 164866 362208 164898
rect 392608 165454 392928 165486
rect 392608 165218 392650 165454
rect 392886 165218 392928 165454
rect 392608 165134 392928 165218
rect 392608 164898 392650 165134
rect 392886 164898 392928 165134
rect 392608 164866 392928 164898
rect 423328 165454 423648 165486
rect 423328 165218 423370 165454
rect 423606 165218 423648 165454
rect 423328 165134 423648 165218
rect 423328 164898 423370 165134
rect 423606 164898 423648 165134
rect 423328 164866 423648 164898
rect 454048 165454 454368 165486
rect 454048 165218 454090 165454
rect 454326 165218 454368 165454
rect 454048 165134 454368 165218
rect 454048 164898 454090 165134
rect 454326 164898 454368 165134
rect 454048 164866 454368 164898
rect 484768 165454 485088 165486
rect 484768 165218 484810 165454
rect 485046 165218 485088 165454
rect 484768 165134 485088 165218
rect 484768 164898 484810 165134
rect 485046 164898 485088 165134
rect 484768 164866 485088 164898
rect 515488 165454 515808 165486
rect 515488 165218 515530 165454
rect 515766 165218 515808 165454
rect 515488 165134 515808 165218
rect 515488 164898 515530 165134
rect 515766 164898 515808 165134
rect 515488 164866 515808 164898
rect 546208 165454 546528 165486
rect 546208 165218 546250 165454
rect 546486 165218 546528 165454
rect 546208 165134 546528 165218
rect 546208 164898 546250 165134
rect 546486 164898 546528 165134
rect 546208 164866 546528 164898
rect 576928 165454 577248 165486
rect 576928 165218 576970 165454
rect 577206 165218 577248 165454
rect 576928 165134 577248 165218
rect 576928 164898 576970 165134
rect 577206 164898 577248 165134
rect 576928 164866 577248 164898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect 8608 147454 8928 147486
rect 8608 147218 8650 147454
rect 8886 147218 8928 147454
rect 8608 147134 8928 147218
rect 8608 146898 8650 147134
rect 8886 146898 8928 147134
rect 8608 146866 8928 146898
rect 39328 147454 39648 147486
rect 39328 147218 39370 147454
rect 39606 147218 39648 147454
rect 39328 147134 39648 147218
rect 39328 146898 39370 147134
rect 39606 146898 39648 147134
rect 39328 146866 39648 146898
rect 70048 147454 70368 147486
rect 70048 147218 70090 147454
rect 70326 147218 70368 147454
rect 70048 147134 70368 147218
rect 70048 146898 70090 147134
rect 70326 146898 70368 147134
rect 70048 146866 70368 146898
rect 100768 147454 101088 147486
rect 100768 147218 100810 147454
rect 101046 147218 101088 147454
rect 100768 147134 101088 147218
rect 100768 146898 100810 147134
rect 101046 146898 101088 147134
rect 100768 146866 101088 146898
rect 131488 147454 131808 147486
rect 131488 147218 131530 147454
rect 131766 147218 131808 147454
rect 131488 147134 131808 147218
rect 131488 146898 131530 147134
rect 131766 146898 131808 147134
rect 131488 146866 131808 146898
rect 162208 147454 162528 147486
rect 162208 147218 162250 147454
rect 162486 147218 162528 147454
rect 162208 147134 162528 147218
rect 162208 146898 162250 147134
rect 162486 146898 162528 147134
rect 162208 146866 162528 146898
rect 192928 147454 193248 147486
rect 192928 147218 192970 147454
rect 193206 147218 193248 147454
rect 192928 147134 193248 147218
rect 192928 146898 192970 147134
rect 193206 146898 193248 147134
rect 192928 146866 193248 146898
rect 223648 147454 223968 147486
rect 223648 147218 223690 147454
rect 223926 147218 223968 147454
rect 223648 147134 223968 147218
rect 223648 146898 223690 147134
rect 223926 146898 223968 147134
rect 223648 146866 223968 146898
rect 254368 147454 254688 147486
rect 254368 147218 254410 147454
rect 254646 147218 254688 147454
rect 254368 147134 254688 147218
rect 254368 146898 254410 147134
rect 254646 146898 254688 147134
rect 254368 146866 254688 146898
rect 285088 147454 285408 147486
rect 285088 147218 285130 147454
rect 285366 147218 285408 147454
rect 285088 147134 285408 147218
rect 285088 146898 285130 147134
rect 285366 146898 285408 147134
rect 285088 146866 285408 146898
rect 315808 147454 316128 147486
rect 315808 147218 315850 147454
rect 316086 147218 316128 147454
rect 315808 147134 316128 147218
rect 315808 146898 315850 147134
rect 316086 146898 316128 147134
rect 315808 146866 316128 146898
rect 346528 147454 346848 147486
rect 346528 147218 346570 147454
rect 346806 147218 346848 147454
rect 346528 147134 346848 147218
rect 346528 146898 346570 147134
rect 346806 146898 346848 147134
rect 346528 146866 346848 146898
rect 377248 147454 377568 147486
rect 377248 147218 377290 147454
rect 377526 147218 377568 147454
rect 377248 147134 377568 147218
rect 377248 146898 377290 147134
rect 377526 146898 377568 147134
rect 377248 146866 377568 146898
rect 407968 147454 408288 147486
rect 407968 147218 408010 147454
rect 408246 147218 408288 147454
rect 407968 147134 408288 147218
rect 407968 146898 408010 147134
rect 408246 146898 408288 147134
rect 407968 146866 408288 146898
rect 438688 147454 439008 147486
rect 438688 147218 438730 147454
rect 438966 147218 439008 147454
rect 438688 147134 439008 147218
rect 438688 146898 438730 147134
rect 438966 146898 439008 147134
rect 438688 146866 439008 146898
rect 469408 147454 469728 147486
rect 469408 147218 469450 147454
rect 469686 147218 469728 147454
rect 469408 147134 469728 147218
rect 469408 146898 469450 147134
rect 469686 146898 469728 147134
rect 469408 146866 469728 146898
rect 500128 147454 500448 147486
rect 500128 147218 500170 147454
rect 500406 147218 500448 147454
rect 500128 147134 500448 147218
rect 500128 146898 500170 147134
rect 500406 146898 500448 147134
rect 500128 146866 500448 146898
rect 530848 147454 531168 147486
rect 530848 147218 530890 147454
rect 531126 147218 531168 147454
rect 530848 147134 531168 147218
rect 530848 146898 530890 147134
rect 531126 146898 531168 147134
rect 530848 146866 531168 146898
rect 561568 147454 561888 147486
rect 561568 147218 561610 147454
rect 561846 147218 561888 147454
rect 561568 147134 561888 147218
rect 561568 146898 561610 147134
rect 561846 146898 561888 147134
rect 561568 146866 561888 146898
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 23968 129454 24288 129486
rect 23968 129218 24010 129454
rect 24246 129218 24288 129454
rect 23968 129134 24288 129218
rect 23968 128898 24010 129134
rect 24246 128898 24288 129134
rect 23968 128866 24288 128898
rect 54688 129454 55008 129486
rect 54688 129218 54730 129454
rect 54966 129218 55008 129454
rect 54688 129134 55008 129218
rect 54688 128898 54730 129134
rect 54966 128898 55008 129134
rect 54688 128866 55008 128898
rect 85408 129454 85728 129486
rect 85408 129218 85450 129454
rect 85686 129218 85728 129454
rect 85408 129134 85728 129218
rect 85408 128898 85450 129134
rect 85686 128898 85728 129134
rect 85408 128866 85728 128898
rect 116128 129454 116448 129486
rect 116128 129218 116170 129454
rect 116406 129218 116448 129454
rect 116128 129134 116448 129218
rect 116128 128898 116170 129134
rect 116406 128898 116448 129134
rect 116128 128866 116448 128898
rect 146848 129454 147168 129486
rect 146848 129218 146890 129454
rect 147126 129218 147168 129454
rect 146848 129134 147168 129218
rect 146848 128898 146890 129134
rect 147126 128898 147168 129134
rect 146848 128866 147168 128898
rect 177568 129454 177888 129486
rect 177568 129218 177610 129454
rect 177846 129218 177888 129454
rect 177568 129134 177888 129218
rect 177568 128898 177610 129134
rect 177846 128898 177888 129134
rect 177568 128866 177888 128898
rect 208288 129454 208608 129486
rect 208288 129218 208330 129454
rect 208566 129218 208608 129454
rect 208288 129134 208608 129218
rect 208288 128898 208330 129134
rect 208566 128898 208608 129134
rect 208288 128866 208608 128898
rect 239008 129454 239328 129486
rect 239008 129218 239050 129454
rect 239286 129218 239328 129454
rect 239008 129134 239328 129218
rect 239008 128898 239050 129134
rect 239286 128898 239328 129134
rect 239008 128866 239328 128898
rect 269728 129454 270048 129486
rect 269728 129218 269770 129454
rect 270006 129218 270048 129454
rect 269728 129134 270048 129218
rect 269728 128898 269770 129134
rect 270006 128898 270048 129134
rect 269728 128866 270048 128898
rect 300448 129454 300768 129486
rect 300448 129218 300490 129454
rect 300726 129218 300768 129454
rect 300448 129134 300768 129218
rect 300448 128898 300490 129134
rect 300726 128898 300768 129134
rect 300448 128866 300768 128898
rect 331168 129454 331488 129486
rect 331168 129218 331210 129454
rect 331446 129218 331488 129454
rect 331168 129134 331488 129218
rect 331168 128898 331210 129134
rect 331446 128898 331488 129134
rect 331168 128866 331488 128898
rect 361888 129454 362208 129486
rect 361888 129218 361930 129454
rect 362166 129218 362208 129454
rect 361888 129134 362208 129218
rect 361888 128898 361930 129134
rect 362166 128898 362208 129134
rect 361888 128866 362208 128898
rect 392608 129454 392928 129486
rect 392608 129218 392650 129454
rect 392886 129218 392928 129454
rect 392608 129134 392928 129218
rect 392608 128898 392650 129134
rect 392886 128898 392928 129134
rect 392608 128866 392928 128898
rect 423328 129454 423648 129486
rect 423328 129218 423370 129454
rect 423606 129218 423648 129454
rect 423328 129134 423648 129218
rect 423328 128898 423370 129134
rect 423606 128898 423648 129134
rect 423328 128866 423648 128898
rect 454048 129454 454368 129486
rect 454048 129218 454090 129454
rect 454326 129218 454368 129454
rect 454048 129134 454368 129218
rect 454048 128898 454090 129134
rect 454326 128898 454368 129134
rect 454048 128866 454368 128898
rect 484768 129454 485088 129486
rect 484768 129218 484810 129454
rect 485046 129218 485088 129454
rect 484768 129134 485088 129218
rect 484768 128898 484810 129134
rect 485046 128898 485088 129134
rect 484768 128866 485088 128898
rect 515488 129454 515808 129486
rect 515488 129218 515530 129454
rect 515766 129218 515808 129454
rect 515488 129134 515808 129218
rect 515488 128898 515530 129134
rect 515766 128898 515808 129134
rect 515488 128866 515808 128898
rect 546208 129454 546528 129486
rect 546208 129218 546250 129454
rect 546486 129218 546528 129454
rect 546208 129134 546528 129218
rect 546208 128898 546250 129134
rect 546486 128898 546528 129134
rect 546208 128866 546528 128898
rect 576928 129454 577248 129486
rect 576928 129218 576970 129454
rect 577206 129218 577248 129454
rect 576928 129134 577248 129218
rect 576928 128898 576970 129134
rect 577206 128898 577248 129134
rect 576928 128866 577248 128898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect 8608 111454 8928 111486
rect 8608 111218 8650 111454
rect 8886 111218 8928 111454
rect 8608 111134 8928 111218
rect 8608 110898 8650 111134
rect 8886 110898 8928 111134
rect 8608 110866 8928 110898
rect 39328 111454 39648 111486
rect 39328 111218 39370 111454
rect 39606 111218 39648 111454
rect 39328 111134 39648 111218
rect 39328 110898 39370 111134
rect 39606 110898 39648 111134
rect 39328 110866 39648 110898
rect 70048 111454 70368 111486
rect 70048 111218 70090 111454
rect 70326 111218 70368 111454
rect 70048 111134 70368 111218
rect 70048 110898 70090 111134
rect 70326 110898 70368 111134
rect 70048 110866 70368 110898
rect 100768 111454 101088 111486
rect 100768 111218 100810 111454
rect 101046 111218 101088 111454
rect 100768 111134 101088 111218
rect 100768 110898 100810 111134
rect 101046 110898 101088 111134
rect 100768 110866 101088 110898
rect 131488 111454 131808 111486
rect 131488 111218 131530 111454
rect 131766 111218 131808 111454
rect 131488 111134 131808 111218
rect 131488 110898 131530 111134
rect 131766 110898 131808 111134
rect 131488 110866 131808 110898
rect 162208 111454 162528 111486
rect 162208 111218 162250 111454
rect 162486 111218 162528 111454
rect 162208 111134 162528 111218
rect 162208 110898 162250 111134
rect 162486 110898 162528 111134
rect 162208 110866 162528 110898
rect 192928 111454 193248 111486
rect 192928 111218 192970 111454
rect 193206 111218 193248 111454
rect 192928 111134 193248 111218
rect 192928 110898 192970 111134
rect 193206 110898 193248 111134
rect 192928 110866 193248 110898
rect 223648 111454 223968 111486
rect 223648 111218 223690 111454
rect 223926 111218 223968 111454
rect 223648 111134 223968 111218
rect 223648 110898 223690 111134
rect 223926 110898 223968 111134
rect 223648 110866 223968 110898
rect 254368 111454 254688 111486
rect 254368 111218 254410 111454
rect 254646 111218 254688 111454
rect 254368 111134 254688 111218
rect 254368 110898 254410 111134
rect 254646 110898 254688 111134
rect 254368 110866 254688 110898
rect 285088 111454 285408 111486
rect 285088 111218 285130 111454
rect 285366 111218 285408 111454
rect 285088 111134 285408 111218
rect 285088 110898 285130 111134
rect 285366 110898 285408 111134
rect 285088 110866 285408 110898
rect 315808 111454 316128 111486
rect 315808 111218 315850 111454
rect 316086 111218 316128 111454
rect 315808 111134 316128 111218
rect 315808 110898 315850 111134
rect 316086 110898 316128 111134
rect 315808 110866 316128 110898
rect 346528 111454 346848 111486
rect 346528 111218 346570 111454
rect 346806 111218 346848 111454
rect 346528 111134 346848 111218
rect 346528 110898 346570 111134
rect 346806 110898 346848 111134
rect 346528 110866 346848 110898
rect 377248 111454 377568 111486
rect 377248 111218 377290 111454
rect 377526 111218 377568 111454
rect 377248 111134 377568 111218
rect 377248 110898 377290 111134
rect 377526 110898 377568 111134
rect 377248 110866 377568 110898
rect 407968 111454 408288 111486
rect 407968 111218 408010 111454
rect 408246 111218 408288 111454
rect 407968 111134 408288 111218
rect 407968 110898 408010 111134
rect 408246 110898 408288 111134
rect 407968 110866 408288 110898
rect 438688 111454 439008 111486
rect 438688 111218 438730 111454
rect 438966 111218 439008 111454
rect 438688 111134 439008 111218
rect 438688 110898 438730 111134
rect 438966 110898 439008 111134
rect 438688 110866 439008 110898
rect 469408 111454 469728 111486
rect 469408 111218 469450 111454
rect 469686 111218 469728 111454
rect 469408 111134 469728 111218
rect 469408 110898 469450 111134
rect 469686 110898 469728 111134
rect 469408 110866 469728 110898
rect 500128 111454 500448 111486
rect 500128 111218 500170 111454
rect 500406 111218 500448 111454
rect 500128 111134 500448 111218
rect 500128 110898 500170 111134
rect 500406 110898 500448 111134
rect 500128 110866 500448 110898
rect 530848 111454 531168 111486
rect 530848 111218 530890 111454
rect 531126 111218 531168 111454
rect 530848 111134 531168 111218
rect 530848 110898 530890 111134
rect 531126 110898 531168 111134
rect 530848 110866 531168 110898
rect 561568 111454 561888 111486
rect 561568 111218 561610 111454
rect 561846 111218 561888 111454
rect 561568 111134 561888 111218
rect 561568 110898 561610 111134
rect 561846 110898 561888 111134
rect 561568 110866 561888 110898
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 23968 93454 24288 93486
rect 23968 93218 24010 93454
rect 24246 93218 24288 93454
rect 23968 93134 24288 93218
rect 23968 92898 24010 93134
rect 24246 92898 24288 93134
rect 23968 92866 24288 92898
rect 54688 93454 55008 93486
rect 54688 93218 54730 93454
rect 54966 93218 55008 93454
rect 54688 93134 55008 93218
rect 54688 92898 54730 93134
rect 54966 92898 55008 93134
rect 54688 92866 55008 92898
rect 85408 93454 85728 93486
rect 85408 93218 85450 93454
rect 85686 93218 85728 93454
rect 85408 93134 85728 93218
rect 85408 92898 85450 93134
rect 85686 92898 85728 93134
rect 85408 92866 85728 92898
rect 116128 93454 116448 93486
rect 116128 93218 116170 93454
rect 116406 93218 116448 93454
rect 116128 93134 116448 93218
rect 116128 92898 116170 93134
rect 116406 92898 116448 93134
rect 116128 92866 116448 92898
rect 146848 93454 147168 93486
rect 146848 93218 146890 93454
rect 147126 93218 147168 93454
rect 146848 93134 147168 93218
rect 146848 92898 146890 93134
rect 147126 92898 147168 93134
rect 146848 92866 147168 92898
rect 177568 93454 177888 93486
rect 177568 93218 177610 93454
rect 177846 93218 177888 93454
rect 177568 93134 177888 93218
rect 177568 92898 177610 93134
rect 177846 92898 177888 93134
rect 177568 92866 177888 92898
rect 208288 93454 208608 93486
rect 208288 93218 208330 93454
rect 208566 93218 208608 93454
rect 208288 93134 208608 93218
rect 208288 92898 208330 93134
rect 208566 92898 208608 93134
rect 208288 92866 208608 92898
rect 239008 93454 239328 93486
rect 239008 93218 239050 93454
rect 239286 93218 239328 93454
rect 239008 93134 239328 93218
rect 239008 92898 239050 93134
rect 239286 92898 239328 93134
rect 239008 92866 239328 92898
rect 269728 93454 270048 93486
rect 269728 93218 269770 93454
rect 270006 93218 270048 93454
rect 269728 93134 270048 93218
rect 269728 92898 269770 93134
rect 270006 92898 270048 93134
rect 269728 92866 270048 92898
rect 300448 93454 300768 93486
rect 300448 93218 300490 93454
rect 300726 93218 300768 93454
rect 300448 93134 300768 93218
rect 300448 92898 300490 93134
rect 300726 92898 300768 93134
rect 300448 92866 300768 92898
rect 331168 93454 331488 93486
rect 331168 93218 331210 93454
rect 331446 93218 331488 93454
rect 331168 93134 331488 93218
rect 331168 92898 331210 93134
rect 331446 92898 331488 93134
rect 331168 92866 331488 92898
rect 361888 93454 362208 93486
rect 361888 93218 361930 93454
rect 362166 93218 362208 93454
rect 361888 93134 362208 93218
rect 361888 92898 361930 93134
rect 362166 92898 362208 93134
rect 361888 92866 362208 92898
rect 392608 93454 392928 93486
rect 392608 93218 392650 93454
rect 392886 93218 392928 93454
rect 392608 93134 392928 93218
rect 392608 92898 392650 93134
rect 392886 92898 392928 93134
rect 392608 92866 392928 92898
rect 423328 93454 423648 93486
rect 423328 93218 423370 93454
rect 423606 93218 423648 93454
rect 423328 93134 423648 93218
rect 423328 92898 423370 93134
rect 423606 92898 423648 93134
rect 423328 92866 423648 92898
rect 454048 93454 454368 93486
rect 454048 93218 454090 93454
rect 454326 93218 454368 93454
rect 454048 93134 454368 93218
rect 454048 92898 454090 93134
rect 454326 92898 454368 93134
rect 454048 92866 454368 92898
rect 484768 93454 485088 93486
rect 484768 93218 484810 93454
rect 485046 93218 485088 93454
rect 484768 93134 485088 93218
rect 484768 92898 484810 93134
rect 485046 92898 485088 93134
rect 484768 92866 485088 92898
rect 515488 93454 515808 93486
rect 515488 93218 515530 93454
rect 515766 93218 515808 93454
rect 515488 93134 515808 93218
rect 515488 92898 515530 93134
rect 515766 92898 515808 93134
rect 515488 92866 515808 92898
rect 546208 93454 546528 93486
rect 546208 93218 546250 93454
rect 546486 93218 546528 93454
rect 546208 93134 546528 93218
rect 546208 92898 546250 93134
rect 546486 92898 546528 93134
rect 546208 92866 546528 92898
rect 576928 93454 577248 93486
rect 576928 93218 576970 93454
rect 577206 93218 577248 93454
rect 576928 93134 577248 93218
rect 576928 92898 576970 93134
rect 577206 92898 577248 93134
rect 576928 92866 577248 92898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect 8608 75454 8928 75486
rect 8608 75218 8650 75454
rect 8886 75218 8928 75454
rect 8608 75134 8928 75218
rect 8608 74898 8650 75134
rect 8886 74898 8928 75134
rect 8608 74866 8928 74898
rect 39328 75454 39648 75486
rect 39328 75218 39370 75454
rect 39606 75218 39648 75454
rect 39328 75134 39648 75218
rect 39328 74898 39370 75134
rect 39606 74898 39648 75134
rect 39328 74866 39648 74898
rect 70048 75454 70368 75486
rect 70048 75218 70090 75454
rect 70326 75218 70368 75454
rect 70048 75134 70368 75218
rect 70048 74898 70090 75134
rect 70326 74898 70368 75134
rect 70048 74866 70368 74898
rect 100768 75454 101088 75486
rect 100768 75218 100810 75454
rect 101046 75218 101088 75454
rect 100768 75134 101088 75218
rect 100768 74898 100810 75134
rect 101046 74898 101088 75134
rect 100768 74866 101088 74898
rect 131488 75454 131808 75486
rect 131488 75218 131530 75454
rect 131766 75218 131808 75454
rect 131488 75134 131808 75218
rect 131488 74898 131530 75134
rect 131766 74898 131808 75134
rect 131488 74866 131808 74898
rect 162208 75454 162528 75486
rect 162208 75218 162250 75454
rect 162486 75218 162528 75454
rect 162208 75134 162528 75218
rect 162208 74898 162250 75134
rect 162486 74898 162528 75134
rect 162208 74866 162528 74898
rect 192928 75454 193248 75486
rect 192928 75218 192970 75454
rect 193206 75218 193248 75454
rect 192928 75134 193248 75218
rect 192928 74898 192970 75134
rect 193206 74898 193248 75134
rect 192928 74866 193248 74898
rect 223648 75454 223968 75486
rect 223648 75218 223690 75454
rect 223926 75218 223968 75454
rect 223648 75134 223968 75218
rect 223648 74898 223690 75134
rect 223926 74898 223968 75134
rect 223648 74866 223968 74898
rect 254368 75454 254688 75486
rect 254368 75218 254410 75454
rect 254646 75218 254688 75454
rect 254368 75134 254688 75218
rect 254368 74898 254410 75134
rect 254646 74898 254688 75134
rect 254368 74866 254688 74898
rect 285088 75454 285408 75486
rect 285088 75218 285130 75454
rect 285366 75218 285408 75454
rect 285088 75134 285408 75218
rect 285088 74898 285130 75134
rect 285366 74898 285408 75134
rect 285088 74866 285408 74898
rect 315808 75454 316128 75486
rect 315808 75218 315850 75454
rect 316086 75218 316128 75454
rect 315808 75134 316128 75218
rect 315808 74898 315850 75134
rect 316086 74898 316128 75134
rect 315808 74866 316128 74898
rect 346528 75454 346848 75486
rect 346528 75218 346570 75454
rect 346806 75218 346848 75454
rect 346528 75134 346848 75218
rect 346528 74898 346570 75134
rect 346806 74898 346848 75134
rect 346528 74866 346848 74898
rect 377248 75454 377568 75486
rect 377248 75218 377290 75454
rect 377526 75218 377568 75454
rect 377248 75134 377568 75218
rect 377248 74898 377290 75134
rect 377526 74898 377568 75134
rect 377248 74866 377568 74898
rect 407968 75454 408288 75486
rect 407968 75218 408010 75454
rect 408246 75218 408288 75454
rect 407968 75134 408288 75218
rect 407968 74898 408010 75134
rect 408246 74898 408288 75134
rect 407968 74866 408288 74898
rect 438688 75454 439008 75486
rect 438688 75218 438730 75454
rect 438966 75218 439008 75454
rect 438688 75134 439008 75218
rect 438688 74898 438730 75134
rect 438966 74898 439008 75134
rect 438688 74866 439008 74898
rect 469408 75454 469728 75486
rect 469408 75218 469450 75454
rect 469686 75218 469728 75454
rect 469408 75134 469728 75218
rect 469408 74898 469450 75134
rect 469686 74898 469728 75134
rect 469408 74866 469728 74898
rect 500128 75454 500448 75486
rect 500128 75218 500170 75454
rect 500406 75218 500448 75454
rect 500128 75134 500448 75218
rect 500128 74898 500170 75134
rect 500406 74898 500448 75134
rect 500128 74866 500448 74898
rect 530848 75454 531168 75486
rect 530848 75218 530890 75454
rect 531126 75218 531168 75454
rect 530848 75134 531168 75218
rect 530848 74898 530890 75134
rect 531126 74898 531168 75134
rect 530848 74866 531168 74898
rect 561568 75454 561888 75486
rect 561568 75218 561610 75454
rect 561846 75218 561888 75454
rect 561568 75134 561888 75218
rect 561568 74898 561610 75134
rect 561846 74898 561888 75134
rect 561568 74866 561888 74898
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 23968 57454 24288 57486
rect 23968 57218 24010 57454
rect 24246 57218 24288 57454
rect 23968 57134 24288 57218
rect 23968 56898 24010 57134
rect 24246 56898 24288 57134
rect 23968 56866 24288 56898
rect 54688 57454 55008 57486
rect 54688 57218 54730 57454
rect 54966 57218 55008 57454
rect 54688 57134 55008 57218
rect 54688 56898 54730 57134
rect 54966 56898 55008 57134
rect 54688 56866 55008 56898
rect 85408 57454 85728 57486
rect 85408 57218 85450 57454
rect 85686 57218 85728 57454
rect 85408 57134 85728 57218
rect 85408 56898 85450 57134
rect 85686 56898 85728 57134
rect 85408 56866 85728 56898
rect 116128 57454 116448 57486
rect 116128 57218 116170 57454
rect 116406 57218 116448 57454
rect 116128 57134 116448 57218
rect 116128 56898 116170 57134
rect 116406 56898 116448 57134
rect 116128 56866 116448 56898
rect 146848 57454 147168 57486
rect 146848 57218 146890 57454
rect 147126 57218 147168 57454
rect 146848 57134 147168 57218
rect 146848 56898 146890 57134
rect 147126 56898 147168 57134
rect 146848 56866 147168 56898
rect 177568 57454 177888 57486
rect 177568 57218 177610 57454
rect 177846 57218 177888 57454
rect 177568 57134 177888 57218
rect 177568 56898 177610 57134
rect 177846 56898 177888 57134
rect 177568 56866 177888 56898
rect 208288 57454 208608 57486
rect 208288 57218 208330 57454
rect 208566 57218 208608 57454
rect 208288 57134 208608 57218
rect 208288 56898 208330 57134
rect 208566 56898 208608 57134
rect 208288 56866 208608 56898
rect 239008 57454 239328 57486
rect 239008 57218 239050 57454
rect 239286 57218 239328 57454
rect 239008 57134 239328 57218
rect 239008 56898 239050 57134
rect 239286 56898 239328 57134
rect 239008 56866 239328 56898
rect 269728 57454 270048 57486
rect 269728 57218 269770 57454
rect 270006 57218 270048 57454
rect 269728 57134 270048 57218
rect 269728 56898 269770 57134
rect 270006 56898 270048 57134
rect 269728 56866 270048 56898
rect 300448 57454 300768 57486
rect 300448 57218 300490 57454
rect 300726 57218 300768 57454
rect 300448 57134 300768 57218
rect 300448 56898 300490 57134
rect 300726 56898 300768 57134
rect 300448 56866 300768 56898
rect 331168 57454 331488 57486
rect 331168 57218 331210 57454
rect 331446 57218 331488 57454
rect 331168 57134 331488 57218
rect 331168 56898 331210 57134
rect 331446 56898 331488 57134
rect 331168 56866 331488 56898
rect 361888 57454 362208 57486
rect 361888 57218 361930 57454
rect 362166 57218 362208 57454
rect 361888 57134 362208 57218
rect 361888 56898 361930 57134
rect 362166 56898 362208 57134
rect 361888 56866 362208 56898
rect 392608 57454 392928 57486
rect 392608 57218 392650 57454
rect 392886 57218 392928 57454
rect 392608 57134 392928 57218
rect 392608 56898 392650 57134
rect 392886 56898 392928 57134
rect 392608 56866 392928 56898
rect 423328 57454 423648 57486
rect 423328 57218 423370 57454
rect 423606 57218 423648 57454
rect 423328 57134 423648 57218
rect 423328 56898 423370 57134
rect 423606 56898 423648 57134
rect 423328 56866 423648 56898
rect 454048 57454 454368 57486
rect 454048 57218 454090 57454
rect 454326 57218 454368 57454
rect 454048 57134 454368 57218
rect 454048 56898 454090 57134
rect 454326 56898 454368 57134
rect 454048 56866 454368 56898
rect 484768 57454 485088 57486
rect 484768 57218 484810 57454
rect 485046 57218 485088 57454
rect 484768 57134 485088 57218
rect 484768 56898 484810 57134
rect 485046 56898 485088 57134
rect 484768 56866 485088 56898
rect 515488 57454 515808 57486
rect 515488 57218 515530 57454
rect 515766 57218 515808 57454
rect 515488 57134 515808 57218
rect 515488 56898 515530 57134
rect 515766 56898 515808 57134
rect 515488 56866 515808 56898
rect 546208 57454 546528 57486
rect 546208 57218 546250 57454
rect 546486 57218 546528 57454
rect 546208 57134 546528 57218
rect 546208 56898 546250 57134
rect 546486 56898 546528 57134
rect 546208 56866 546528 56898
rect 576928 57454 577248 57486
rect 576928 57218 576970 57454
rect 577206 57218 577248 57454
rect 576928 57134 577248 57218
rect 576928 56898 576970 57134
rect 577206 56898 577248 57134
rect 576928 56866 577248 56898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect 8608 39454 8928 39486
rect 8608 39218 8650 39454
rect 8886 39218 8928 39454
rect 8608 39134 8928 39218
rect 8608 38898 8650 39134
rect 8886 38898 8928 39134
rect 8608 38866 8928 38898
rect 39328 39454 39648 39486
rect 39328 39218 39370 39454
rect 39606 39218 39648 39454
rect 39328 39134 39648 39218
rect 39328 38898 39370 39134
rect 39606 38898 39648 39134
rect 39328 38866 39648 38898
rect 70048 39454 70368 39486
rect 70048 39218 70090 39454
rect 70326 39218 70368 39454
rect 70048 39134 70368 39218
rect 70048 38898 70090 39134
rect 70326 38898 70368 39134
rect 70048 38866 70368 38898
rect 100768 39454 101088 39486
rect 100768 39218 100810 39454
rect 101046 39218 101088 39454
rect 100768 39134 101088 39218
rect 100768 38898 100810 39134
rect 101046 38898 101088 39134
rect 100768 38866 101088 38898
rect 131488 39454 131808 39486
rect 131488 39218 131530 39454
rect 131766 39218 131808 39454
rect 131488 39134 131808 39218
rect 131488 38898 131530 39134
rect 131766 38898 131808 39134
rect 131488 38866 131808 38898
rect 162208 39454 162528 39486
rect 162208 39218 162250 39454
rect 162486 39218 162528 39454
rect 162208 39134 162528 39218
rect 162208 38898 162250 39134
rect 162486 38898 162528 39134
rect 162208 38866 162528 38898
rect 192928 39454 193248 39486
rect 192928 39218 192970 39454
rect 193206 39218 193248 39454
rect 192928 39134 193248 39218
rect 192928 38898 192970 39134
rect 193206 38898 193248 39134
rect 192928 38866 193248 38898
rect 223648 39454 223968 39486
rect 223648 39218 223690 39454
rect 223926 39218 223968 39454
rect 223648 39134 223968 39218
rect 223648 38898 223690 39134
rect 223926 38898 223968 39134
rect 223648 38866 223968 38898
rect 254368 39454 254688 39486
rect 254368 39218 254410 39454
rect 254646 39218 254688 39454
rect 254368 39134 254688 39218
rect 254368 38898 254410 39134
rect 254646 38898 254688 39134
rect 254368 38866 254688 38898
rect 285088 39454 285408 39486
rect 285088 39218 285130 39454
rect 285366 39218 285408 39454
rect 285088 39134 285408 39218
rect 285088 38898 285130 39134
rect 285366 38898 285408 39134
rect 285088 38866 285408 38898
rect 315808 39454 316128 39486
rect 315808 39218 315850 39454
rect 316086 39218 316128 39454
rect 315808 39134 316128 39218
rect 315808 38898 315850 39134
rect 316086 38898 316128 39134
rect 315808 38866 316128 38898
rect 346528 39454 346848 39486
rect 346528 39218 346570 39454
rect 346806 39218 346848 39454
rect 346528 39134 346848 39218
rect 346528 38898 346570 39134
rect 346806 38898 346848 39134
rect 346528 38866 346848 38898
rect 377248 39454 377568 39486
rect 377248 39218 377290 39454
rect 377526 39218 377568 39454
rect 377248 39134 377568 39218
rect 377248 38898 377290 39134
rect 377526 38898 377568 39134
rect 377248 38866 377568 38898
rect 407968 39454 408288 39486
rect 407968 39218 408010 39454
rect 408246 39218 408288 39454
rect 407968 39134 408288 39218
rect 407968 38898 408010 39134
rect 408246 38898 408288 39134
rect 407968 38866 408288 38898
rect 438688 39454 439008 39486
rect 438688 39218 438730 39454
rect 438966 39218 439008 39454
rect 438688 39134 439008 39218
rect 438688 38898 438730 39134
rect 438966 38898 439008 39134
rect 438688 38866 439008 38898
rect 469408 39454 469728 39486
rect 469408 39218 469450 39454
rect 469686 39218 469728 39454
rect 469408 39134 469728 39218
rect 469408 38898 469450 39134
rect 469686 38898 469728 39134
rect 469408 38866 469728 38898
rect 500128 39454 500448 39486
rect 500128 39218 500170 39454
rect 500406 39218 500448 39454
rect 500128 39134 500448 39218
rect 500128 38898 500170 39134
rect 500406 38898 500448 39134
rect 500128 38866 500448 38898
rect 530848 39454 531168 39486
rect 530848 39218 530890 39454
rect 531126 39218 531168 39454
rect 530848 39134 531168 39218
rect 530848 38898 530890 39134
rect 531126 38898 531168 39134
rect 530848 38866 531168 38898
rect 561568 39454 561888 39486
rect 561568 39218 561610 39454
rect 561846 39218 561888 39454
rect 561568 39134 561888 39218
rect 561568 38898 561610 39134
rect 561846 38898 561888 39134
rect 561568 38866 561888 38898
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 23968 21454 24288 21486
rect 23968 21218 24010 21454
rect 24246 21218 24288 21454
rect 23968 21134 24288 21218
rect 23968 20898 24010 21134
rect 24246 20898 24288 21134
rect 23968 20866 24288 20898
rect 54688 21454 55008 21486
rect 54688 21218 54730 21454
rect 54966 21218 55008 21454
rect 54688 21134 55008 21218
rect 54688 20898 54730 21134
rect 54966 20898 55008 21134
rect 54688 20866 55008 20898
rect 85408 21454 85728 21486
rect 85408 21218 85450 21454
rect 85686 21218 85728 21454
rect 85408 21134 85728 21218
rect 85408 20898 85450 21134
rect 85686 20898 85728 21134
rect 85408 20866 85728 20898
rect 116128 21454 116448 21486
rect 116128 21218 116170 21454
rect 116406 21218 116448 21454
rect 116128 21134 116448 21218
rect 116128 20898 116170 21134
rect 116406 20898 116448 21134
rect 116128 20866 116448 20898
rect 146848 21454 147168 21486
rect 146848 21218 146890 21454
rect 147126 21218 147168 21454
rect 146848 21134 147168 21218
rect 146848 20898 146890 21134
rect 147126 20898 147168 21134
rect 146848 20866 147168 20898
rect 177568 21454 177888 21486
rect 177568 21218 177610 21454
rect 177846 21218 177888 21454
rect 177568 21134 177888 21218
rect 177568 20898 177610 21134
rect 177846 20898 177888 21134
rect 177568 20866 177888 20898
rect 208288 21454 208608 21486
rect 208288 21218 208330 21454
rect 208566 21218 208608 21454
rect 208288 21134 208608 21218
rect 208288 20898 208330 21134
rect 208566 20898 208608 21134
rect 208288 20866 208608 20898
rect 239008 21454 239328 21486
rect 239008 21218 239050 21454
rect 239286 21218 239328 21454
rect 239008 21134 239328 21218
rect 239008 20898 239050 21134
rect 239286 20898 239328 21134
rect 239008 20866 239328 20898
rect 269728 21454 270048 21486
rect 269728 21218 269770 21454
rect 270006 21218 270048 21454
rect 269728 21134 270048 21218
rect 269728 20898 269770 21134
rect 270006 20898 270048 21134
rect 269728 20866 270048 20898
rect 300448 21454 300768 21486
rect 300448 21218 300490 21454
rect 300726 21218 300768 21454
rect 300448 21134 300768 21218
rect 300448 20898 300490 21134
rect 300726 20898 300768 21134
rect 300448 20866 300768 20898
rect 331168 21454 331488 21486
rect 331168 21218 331210 21454
rect 331446 21218 331488 21454
rect 331168 21134 331488 21218
rect 331168 20898 331210 21134
rect 331446 20898 331488 21134
rect 331168 20866 331488 20898
rect 361888 21454 362208 21486
rect 361888 21218 361930 21454
rect 362166 21218 362208 21454
rect 361888 21134 362208 21218
rect 361888 20898 361930 21134
rect 362166 20898 362208 21134
rect 361888 20866 362208 20898
rect 392608 21454 392928 21486
rect 392608 21218 392650 21454
rect 392886 21218 392928 21454
rect 392608 21134 392928 21218
rect 392608 20898 392650 21134
rect 392886 20898 392928 21134
rect 392608 20866 392928 20898
rect 423328 21454 423648 21486
rect 423328 21218 423370 21454
rect 423606 21218 423648 21454
rect 423328 21134 423648 21218
rect 423328 20898 423370 21134
rect 423606 20898 423648 21134
rect 423328 20866 423648 20898
rect 454048 21454 454368 21486
rect 454048 21218 454090 21454
rect 454326 21218 454368 21454
rect 454048 21134 454368 21218
rect 454048 20898 454090 21134
rect 454326 20898 454368 21134
rect 454048 20866 454368 20898
rect 484768 21454 485088 21486
rect 484768 21218 484810 21454
rect 485046 21218 485088 21454
rect 484768 21134 485088 21218
rect 484768 20898 484810 21134
rect 485046 20898 485088 21134
rect 484768 20866 485088 20898
rect 515488 21454 515808 21486
rect 515488 21218 515530 21454
rect 515766 21218 515808 21454
rect 515488 21134 515808 21218
rect 515488 20898 515530 21134
rect 515766 20898 515808 21134
rect 515488 20866 515808 20898
rect 546208 21454 546528 21486
rect 546208 21218 546250 21454
rect 546486 21218 546528 21454
rect 546208 21134 546528 21218
rect 546208 20898 546250 21134
rect 546486 20898 546528 21134
rect 546208 20866 546528 20898
rect 576928 21454 577248 21486
rect 576928 21218 576970 21454
rect 577206 21218 577248 21454
rect 576928 21134 577248 21218
rect 576928 20898 576970 21134
rect 577206 20898 577248 21134
rect 576928 20866 577248 20898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 -346 2414 2400
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 2400
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 2400
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 2400
rect 19794 -1306 20414 2400
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 -3226 24134 2400
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 2400
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 2400
rect 37794 -346 38414 2400
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 -2266 42134 2400
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 -4186 45854 2400
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 2400
rect 55794 -1306 56414 2400
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 -3226 60134 2400
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 2400
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 2400
rect 73794 -346 74414 2400
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 -2266 78134 2400
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 -4186 81854 2400
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 2400
rect 91794 -1306 92414 2400
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 -3226 96134 2400
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 2400
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 2400
rect 109794 -346 110414 2400
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 -2266 114134 2400
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 -4186 117854 2400
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 2400
rect 127794 -1306 128414 2400
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 -3226 132134 2400
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 2400
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 2400
rect 145794 -346 146414 2400
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 -2266 150134 2400
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 -4186 153854 2400
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 2400
rect 163794 -1306 164414 2400
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 2400
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 2400
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 2400
rect 181794 -346 182414 2400
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 -2266 186134 2400
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 2400
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 2400
rect 199794 -1306 200414 2400
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 -3226 204134 2400
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 2400
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 2400
rect 217794 -346 218414 2400
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 -2266 222134 2400
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 -4186 225854 2400
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 2400
rect 235794 -1306 236414 2400
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 -3226 240134 2400
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 2400
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 2400
rect 253794 -346 254414 2400
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 -2266 258134 2400
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 -4186 261854 2400
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 2400
rect 271794 -1306 272414 2400
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 -3226 276134 2400
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 2400
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 2400
rect 289794 -346 290414 2400
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 -2266 294134 2400
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 2400
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 2400
rect 307794 -1306 308414 2400
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 -3226 312134 2400
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 2400
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 2400
rect 325794 -346 326414 2400
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 -2266 330134 2400
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 -4186 333854 2400
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 2400
rect 343794 -1306 344414 2400
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 -3226 348134 2400
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 2400
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 2400
rect 361794 -346 362414 2400
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 -2266 366134 2400
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 2400
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 2400
rect 379794 -1306 380414 2400
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 -3226 384134 2400
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 2400
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 2400
rect 397794 -346 398414 2400
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 -2266 402134 2400
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 -4186 405854 2400
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 2400
rect 415794 -1306 416414 2400
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 -3226 420134 2400
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 2400
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 2400
rect 433794 -346 434414 2400
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 -2266 438134 2400
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 -4186 441854 2400
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 2400
rect 451794 -1306 452414 2400
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 -3226 456134 2400
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 2400
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 2400
rect 469794 -346 470414 2400
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 -2266 474134 2400
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 -4186 477854 2400
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 2400
rect 487794 -1306 488414 2400
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 -3226 492134 2400
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 2400
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 2400
rect 505794 -346 506414 2400
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 -2266 510134 2400
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 -4186 513854 2400
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 2400
rect 523794 -1306 524414 2400
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 -3226 528134 2400
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 2400
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 2400
rect 541794 -346 542414 2400
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 -2266 546134 2400
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 -4186 549854 2400
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 2400
rect 559794 -1306 560414 2400
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 -3226 564134 2400
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 -5146 567854 2400
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 2400
rect 577794 -346 578414 2400
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 -2266 582134 2400
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect 8650 687218 8886 687454
rect 8650 686898 8886 687134
rect 39370 687218 39606 687454
rect 39370 686898 39606 687134
rect 70090 687218 70326 687454
rect 70090 686898 70326 687134
rect 100810 687218 101046 687454
rect 100810 686898 101046 687134
rect 131530 687218 131766 687454
rect 131530 686898 131766 687134
rect 162250 687218 162486 687454
rect 162250 686898 162486 687134
rect 192970 687218 193206 687454
rect 192970 686898 193206 687134
rect 223690 687218 223926 687454
rect 223690 686898 223926 687134
rect 254410 687218 254646 687454
rect 254410 686898 254646 687134
rect 285130 687218 285366 687454
rect 285130 686898 285366 687134
rect 315850 687218 316086 687454
rect 315850 686898 316086 687134
rect 346570 687218 346806 687454
rect 346570 686898 346806 687134
rect 377290 687218 377526 687454
rect 377290 686898 377526 687134
rect 408010 687218 408246 687454
rect 408010 686898 408246 687134
rect 438730 687218 438966 687454
rect 438730 686898 438966 687134
rect 469450 687218 469686 687454
rect 469450 686898 469686 687134
rect 500170 687218 500406 687454
rect 500170 686898 500406 687134
rect 530890 687218 531126 687454
rect 530890 686898 531126 687134
rect 561610 687218 561846 687454
rect 561610 686898 561846 687134
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 24010 669218 24246 669454
rect 24010 668898 24246 669134
rect 54730 669218 54966 669454
rect 54730 668898 54966 669134
rect 85450 669218 85686 669454
rect 85450 668898 85686 669134
rect 116170 669218 116406 669454
rect 116170 668898 116406 669134
rect 146890 669218 147126 669454
rect 146890 668898 147126 669134
rect 177610 669218 177846 669454
rect 177610 668898 177846 669134
rect 208330 669218 208566 669454
rect 208330 668898 208566 669134
rect 239050 669218 239286 669454
rect 239050 668898 239286 669134
rect 269770 669218 270006 669454
rect 269770 668898 270006 669134
rect 300490 669218 300726 669454
rect 300490 668898 300726 669134
rect 331210 669218 331446 669454
rect 331210 668898 331446 669134
rect 361930 669218 362166 669454
rect 361930 668898 362166 669134
rect 392650 669218 392886 669454
rect 392650 668898 392886 669134
rect 423370 669218 423606 669454
rect 423370 668898 423606 669134
rect 454090 669218 454326 669454
rect 454090 668898 454326 669134
rect 484810 669218 485046 669454
rect 484810 668898 485046 669134
rect 515530 669218 515766 669454
rect 515530 668898 515766 669134
rect 546250 669218 546486 669454
rect 546250 668898 546486 669134
rect 576970 669218 577206 669454
rect 576970 668898 577206 669134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect 8650 651218 8886 651454
rect 8650 650898 8886 651134
rect 39370 651218 39606 651454
rect 39370 650898 39606 651134
rect 70090 651218 70326 651454
rect 70090 650898 70326 651134
rect 100810 651218 101046 651454
rect 100810 650898 101046 651134
rect 131530 651218 131766 651454
rect 131530 650898 131766 651134
rect 162250 651218 162486 651454
rect 162250 650898 162486 651134
rect 192970 651218 193206 651454
rect 192970 650898 193206 651134
rect 223690 651218 223926 651454
rect 223690 650898 223926 651134
rect 254410 651218 254646 651454
rect 254410 650898 254646 651134
rect 285130 651218 285366 651454
rect 285130 650898 285366 651134
rect 315850 651218 316086 651454
rect 315850 650898 316086 651134
rect 346570 651218 346806 651454
rect 346570 650898 346806 651134
rect 377290 651218 377526 651454
rect 377290 650898 377526 651134
rect 408010 651218 408246 651454
rect 408010 650898 408246 651134
rect 438730 651218 438966 651454
rect 438730 650898 438966 651134
rect 469450 651218 469686 651454
rect 469450 650898 469686 651134
rect 500170 651218 500406 651454
rect 500170 650898 500406 651134
rect 530890 651218 531126 651454
rect 530890 650898 531126 651134
rect 561610 651218 561846 651454
rect 561610 650898 561846 651134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 24010 633218 24246 633454
rect 24010 632898 24246 633134
rect 54730 633218 54966 633454
rect 54730 632898 54966 633134
rect 85450 633218 85686 633454
rect 85450 632898 85686 633134
rect 116170 633218 116406 633454
rect 116170 632898 116406 633134
rect 146890 633218 147126 633454
rect 146890 632898 147126 633134
rect 177610 633218 177846 633454
rect 177610 632898 177846 633134
rect 208330 633218 208566 633454
rect 208330 632898 208566 633134
rect 239050 633218 239286 633454
rect 239050 632898 239286 633134
rect 269770 633218 270006 633454
rect 269770 632898 270006 633134
rect 300490 633218 300726 633454
rect 300490 632898 300726 633134
rect 331210 633218 331446 633454
rect 331210 632898 331446 633134
rect 361930 633218 362166 633454
rect 361930 632898 362166 633134
rect 392650 633218 392886 633454
rect 392650 632898 392886 633134
rect 423370 633218 423606 633454
rect 423370 632898 423606 633134
rect 454090 633218 454326 633454
rect 454090 632898 454326 633134
rect 484810 633218 485046 633454
rect 484810 632898 485046 633134
rect 515530 633218 515766 633454
rect 515530 632898 515766 633134
rect 546250 633218 546486 633454
rect 546250 632898 546486 633134
rect 576970 633218 577206 633454
rect 576970 632898 577206 633134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect 8650 615218 8886 615454
rect 8650 614898 8886 615134
rect 39370 615218 39606 615454
rect 39370 614898 39606 615134
rect 70090 615218 70326 615454
rect 70090 614898 70326 615134
rect 100810 615218 101046 615454
rect 100810 614898 101046 615134
rect 131530 615218 131766 615454
rect 131530 614898 131766 615134
rect 162250 615218 162486 615454
rect 162250 614898 162486 615134
rect 192970 615218 193206 615454
rect 192970 614898 193206 615134
rect 223690 615218 223926 615454
rect 223690 614898 223926 615134
rect 254410 615218 254646 615454
rect 254410 614898 254646 615134
rect 285130 615218 285366 615454
rect 285130 614898 285366 615134
rect 315850 615218 316086 615454
rect 315850 614898 316086 615134
rect 346570 615218 346806 615454
rect 346570 614898 346806 615134
rect 377290 615218 377526 615454
rect 377290 614898 377526 615134
rect 408010 615218 408246 615454
rect 408010 614898 408246 615134
rect 438730 615218 438966 615454
rect 438730 614898 438966 615134
rect 469450 615218 469686 615454
rect 469450 614898 469686 615134
rect 500170 615218 500406 615454
rect 500170 614898 500406 615134
rect 530890 615218 531126 615454
rect 530890 614898 531126 615134
rect 561610 615218 561846 615454
rect 561610 614898 561846 615134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 24010 597218 24246 597454
rect 24010 596898 24246 597134
rect 54730 597218 54966 597454
rect 54730 596898 54966 597134
rect 85450 597218 85686 597454
rect 85450 596898 85686 597134
rect 116170 597218 116406 597454
rect 116170 596898 116406 597134
rect 146890 597218 147126 597454
rect 146890 596898 147126 597134
rect 177610 597218 177846 597454
rect 177610 596898 177846 597134
rect 208330 597218 208566 597454
rect 208330 596898 208566 597134
rect 239050 597218 239286 597454
rect 239050 596898 239286 597134
rect 269770 597218 270006 597454
rect 269770 596898 270006 597134
rect 300490 597218 300726 597454
rect 300490 596898 300726 597134
rect 331210 597218 331446 597454
rect 331210 596898 331446 597134
rect 361930 597218 362166 597454
rect 361930 596898 362166 597134
rect 392650 597218 392886 597454
rect 392650 596898 392886 597134
rect 423370 597218 423606 597454
rect 423370 596898 423606 597134
rect 454090 597218 454326 597454
rect 454090 596898 454326 597134
rect 484810 597218 485046 597454
rect 484810 596898 485046 597134
rect 515530 597218 515766 597454
rect 515530 596898 515766 597134
rect 546250 597218 546486 597454
rect 546250 596898 546486 597134
rect 576970 597218 577206 597454
rect 576970 596898 577206 597134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect 8650 579218 8886 579454
rect 8650 578898 8886 579134
rect 39370 579218 39606 579454
rect 39370 578898 39606 579134
rect 70090 579218 70326 579454
rect 70090 578898 70326 579134
rect 100810 579218 101046 579454
rect 100810 578898 101046 579134
rect 131530 579218 131766 579454
rect 131530 578898 131766 579134
rect 162250 579218 162486 579454
rect 162250 578898 162486 579134
rect 192970 579218 193206 579454
rect 192970 578898 193206 579134
rect 223690 579218 223926 579454
rect 223690 578898 223926 579134
rect 254410 579218 254646 579454
rect 254410 578898 254646 579134
rect 285130 579218 285366 579454
rect 285130 578898 285366 579134
rect 315850 579218 316086 579454
rect 315850 578898 316086 579134
rect 346570 579218 346806 579454
rect 346570 578898 346806 579134
rect 377290 579218 377526 579454
rect 377290 578898 377526 579134
rect 408010 579218 408246 579454
rect 408010 578898 408246 579134
rect 438730 579218 438966 579454
rect 438730 578898 438966 579134
rect 469450 579218 469686 579454
rect 469450 578898 469686 579134
rect 500170 579218 500406 579454
rect 500170 578898 500406 579134
rect 530890 579218 531126 579454
rect 530890 578898 531126 579134
rect 561610 579218 561846 579454
rect 561610 578898 561846 579134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 24010 561218 24246 561454
rect 24010 560898 24246 561134
rect 54730 561218 54966 561454
rect 54730 560898 54966 561134
rect 85450 561218 85686 561454
rect 85450 560898 85686 561134
rect 116170 561218 116406 561454
rect 116170 560898 116406 561134
rect 146890 561218 147126 561454
rect 146890 560898 147126 561134
rect 177610 561218 177846 561454
rect 177610 560898 177846 561134
rect 208330 561218 208566 561454
rect 208330 560898 208566 561134
rect 239050 561218 239286 561454
rect 239050 560898 239286 561134
rect 269770 561218 270006 561454
rect 269770 560898 270006 561134
rect 300490 561218 300726 561454
rect 300490 560898 300726 561134
rect 331210 561218 331446 561454
rect 331210 560898 331446 561134
rect 361930 561218 362166 561454
rect 361930 560898 362166 561134
rect 392650 561218 392886 561454
rect 392650 560898 392886 561134
rect 423370 561218 423606 561454
rect 423370 560898 423606 561134
rect 454090 561218 454326 561454
rect 454090 560898 454326 561134
rect 484810 561218 485046 561454
rect 484810 560898 485046 561134
rect 515530 561218 515766 561454
rect 515530 560898 515766 561134
rect 546250 561218 546486 561454
rect 546250 560898 546486 561134
rect 576970 561218 577206 561454
rect 576970 560898 577206 561134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect 8650 543218 8886 543454
rect 8650 542898 8886 543134
rect 39370 543218 39606 543454
rect 39370 542898 39606 543134
rect 70090 543218 70326 543454
rect 70090 542898 70326 543134
rect 100810 543218 101046 543454
rect 100810 542898 101046 543134
rect 131530 543218 131766 543454
rect 131530 542898 131766 543134
rect 162250 543218 162486 543454
rect 162250 542898 162486 543134
rect 192970 543218 193206 543454
rect 192970 542898 193206 543134
rect 223690 543218 223926 543454
rect 223690 542898 223926 543134
rect 254410 543218 254646 543454
rect 254410 542898 254646 543134
rect 285130 543218 285366 543454
rect 285130 542898 285366 543134
rect 315850 543218 316086 543454
rect 315850 542898 316086 543134
rect 346570 543218 346806 543454
rect 346570 542898 346806 543134
rect 377290 543218 377526 543454
rect 377290 542898 377526 543134
rect 408010 543218 408246 543454
rect 408010 542898 408246 543134
rect 438730 543218 438966 543454
rect 438730 542898 438966 543134
rect 469450 543218 469686 543454
rect 469450 542898 469686 543134
rect 500170 543218 500406 543454
rect 500170 542898 500406 543134
rect 530890 543218 531126 543454
rect 530890 542898 531126 543134
rect 561610 543218 561846 543454
rect 561610 542898 561846 543134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 24010 525218 24246 525454
rect 24010 524898 24246 525134
rect 54730 525218 54966 525454
rect 54730 524898 54966 525134
rect 85450 525218 85686 525454
rect 85450 524898 85686 525134
rect 116170 525218 116406 525454
rect 116170 524898 116406 525134
rect 146890 525218 147126 525454
rect 146890 524898 147126 525134
rect 177610 525218 177846 525454
rect 177610 524898 177846 525134
rect 208330 525218 208566 525454
rect 208330 524898 208566 525134
rect 239050 525218 239286 525454
rect 239050 524898 239286 525134
rect 269770 525218 270006 525454
rect 269770 524898 270006 525134
rect 300490 525218 300726 525454
rect 300490 524898 300726 525134
rect 331210 525218 331446 525454
rect 331210 524898 331446 525134
rect 361930 525218 362166 525454
rect 361930 524898 362166 525134
rect 392650 525218 392886 525454
rect 392650 524898 392886 525134
rect 423370 525218 423606 525454
rect 423370 524898 423606 525134
rect 454090 525218 454326 525454
rect 454090 524898 454326 525134
rect 484810 525218 485046 525454
rect 484810 524898 485046 525134
rect 515530 525218 515766 525454
rect 515530 524898 515766 525134
rect 546250 525218 546486 525454
rect 546250 524898 546486 525134
rect 576970 525218 577206 525454
rect 576970 524898 577206 525134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect 8650 507218 8886 507454
rect 8650 506898 8886 507134
rect 39370 507218 39606 507454
rect 39370 506898 39606 507134
rect 70090 507218 70326 507454
rect 70090 506898 70326 507134
rect 100810 507218 101046 507454
rect 100810 506898 101046 507134
rect 131530 507218 131766 507454
rect 131530 506898 131766 507134
rect 162250 507218 162486 507454
rect 162250 506898 162486 507134
rect 192970 507218 193206 507454
rect 192970 506898 193206 507134
rect 223690 507218 223926 507454
rect 223690 506898 223926 507134
rect 254410 507218 254646 507454
rect 254410 506898 254646 507134
rect 285130 507218 285366 507454
rect 285130 506898 285366 507134
rect 315850 507218 316086 507454
rect 315850 506898 316086 507134
rect 346570 507218 346806 507454
rect 346570 506898 346806 507134
rect 377290 507218 377526 507454
rect 377290 506898 377526 507134
rect 408010 507218 408246 507454
rect 408010 506898 408246 507134
rect 438730 507218 438966 507454
rect 438730 506898 438966 507134
rect 469450 507218 469686 507454
rect 469450 506898 469686 507134
rect 500170 507218 500406 507454
rect 500170 506898 500406 507134
rect 530890 507218 531126 507454
rect 530890 506898 531126 507134
rect 561610 507218 561846 507454
rect 561610 506898 561846 507134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 24010 489218 24246 489454
rect 24010 488898 24246 489134
rect 54730 489218 54966 489454
rect 54730 488898 54966 489134
rect 85450 489218 85686 489454
rect 85450 488898 85686 489134
rect 116170 489218 116406 489454
rect 116170 488898 116406 489134
rect 146890 489218 147126 489454
rect 146890 488898 147126 489134
rect 177610 489218 177846 489454
rect 177610 488898 177846 489134
rect 208330 489218 208566 489454
rect 208330 488898 208566 489134
rect 239050 489218 239286 489454
rect 239050 488898 239286 489134
rect 269770 489218 270006 489454
rect 269770 488898 270006 489134
rect 300490 489218 300726 489454
rect 300490 488898 300726 489134
rect 331210 489218 331446 489454
rect 331210 488898 331446 489134
rect 361930 489218 362166 489454
rect 361930 488898 362166 489134
rect 392650 489218 392886 489454
rect 392650 488898 392886 489134
rect 423370 489218 423606 489454
rect 423370 488898 423606 489134
rect 454090 489218 454326 489454
rect 454090 488898 454326 489134
rect 484810 489218 485046 489454
rect 484810 488898 485046 489134
rect 515530 489218 515766 489454
rect 515530 488898 515766 489134
rect 546250 489218 546486 489454
rect 546250 488898 546486 489134
rect 576970 489218 577206 489454
rect 576970 488898 577206 489134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect 8650 471218 8886 471454
rect 8650 470898 8886 471134
rect 39370 471218 39606 471454
rect 39370 470898 39606 471134
rect 70090 471218 70326 471454
rect 70090 470898 70326 471134
rect 100810 471218 101046 471454
rect 100810 470898 101046 471134
rect 131530 471218 131766 471454
rect 131530 470898 131766 471134
rect 162250 471218 162486 471454
rect 162250 470898 162486 471134
rect 192970 471218 193206 471454
rect 192970 470898 193206 471134
rect 223690 471218 223926 471454
rect 223690 470898 223926 471134
rect 254410 471218 254646 471454
rect 254410 470898 254646 471134
rect 285130 471218 285366 471454
rect 285130 470898 285366 471134
rect 315850 471218 316086 471454
rect 315850 470898 316086 471134
rect 346570 471218 346806 471454
rect 346570 470898 346806 471134
rect 377290 471218 377526 471454
rect 377290 470898 377526 471134
rect 408010 471218 408246 471454
rect 408010 470898 408246 471134
rect 438730 471218 438966 471454
rect 438730 470898 438966 471134
rect 469450 471218 469686 471454
rect 469450 470898 469686 471134
rect 500170 471218 500406 471454
rect 500170 470898 500406 471134
rect 530890 471218 531126 471454
rect 530890 470898 531126 471134
rect 561610 471218 561846 471454
rect 561610 470898 561846 471134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 24010 453218 24246 453454
rect 24010 452898 24246 453134
rect 54730 453218 54966 453454
rect 54730 452898 54966 453134
rect 85450 453218 85686 453454
rect 85450 452898 85686 453134
rect 116170 453218 116406 453454
rect 116170 452898 116406 453134
rect 146890 453218 147126 453454
rect 146890 452898 147126 453134
rect 177610 453218 177846 453454
rect 177610 452898 177846 453134
rect 208330 453218 208566 453454
rect 208330 452898 208566 453134
rect 239050 453218 239286 453454
rect 239050 452898 239286 453134
rect 269770 453218 270006 453454
rect 269770 452898 270006 453134
rect 300490 453218 300726 453454
rect 300490 452898 300726 453134
rect 331210 453218 331446 453454
rect 331210 452898 331446 453134
rect 361930 453218 362166 453454
rect 361930 452898 362166 453134
rect 392650 453218 392886 453454
rect 392650 452898 392886 453134
rect 423370 453218 423606 453454
rect 423370 452898 423606 453134
rect 454090 453218 454326 453454
rect 454090 452898 454326 453134
rect 484810 453218 485046 453454
rect 484810 452898 485046 453134
rect 515530 453218 515766 453454
rect 515530 452898 515766 453134
rect 546250 453218 546486 453454
rect 546250 452898 546486 453134
rect 576970 453218 577206 453454
rect 576970 452898 577206 453134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect 8650 435218 8886 435454
rect 8650 434898 8886 435134
rect 39370 435218 39606 435454
rect 39370 434898 39606 435134
rect 70090 435218 70326 435454
rect 70090 434898 70326 435134
rect 100810 435218 101046 435454
rect 100810 434898 101046 435134
rect 131530 435218 131766 435454
rect 131530 434898 131766 435134
rect 162250 435218 162486 435454
rect 162250 434898 162486 435134
rect 192970 435218 193206 435454
rect 192970 434898 193206 435134
rect 223690 435218 223926 435454
rect 223690 434898 223926 435134
rect 254410 435218 254646 435454
rect 254410 434898 254646 435134
rect 285130 435218 285366 435454
rect 285130 434898 285366 435134
rect 315850 435218 316086 435454
rect 315850 434898 316086 435134
rect 346570 435218 346806 435454
rect 346570 434898 346806 435134
rect 377290 435218 377526 435454
rect 377290 434898 377526 435134
rect 408010 435218 408246 435454
rect 408010 434898 408246 435134
rect 438730 435218 438966 435454
rect 438730 434898 438966 435134
rect 469450 435218 469686 435454
rect 469450 434898 469686 435134
rect 500170 435218 500406 435454
rect 500170 434898 500406 435134
rect 530890 435218 531126 435454
rect 530890 434898 531126 435134
rect 561610 435218 561846 435454
rect 561610 434898 561846 435134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 24010 417218 24246 417454
rect 24010 416898 24246 417134
rect 54730 417218 54966 417454
rect 54730 416898 54966 417134
rect 85450 417218 85686 417454
rect 85450 416898 85686 417134
rect 116170 417218 116406 417454
rect 116170 416898 116406 417134
rect 146890 417218 147126 417454
rect 146890 416898 147126 417134
rect 177610 417218 177846 417454
rect 177610 416898 177846 417134
rect 208330 417218 208566 417454
rect 208330 416898 208566 417134
rect 239050 417218 239286 417454
rect 239050 416898 239286 417134
rect 269770 417218 270006 417454
rect 269770 416898 270006 417134
rect 300490 417218 300726 417454
rect 300490 416898 300726 417134
rect 331210 417218 331446 417454
rect 331210 416898 331446 417134
rect 361930 417218 362166 417454
rect 361930 416898 362166 417134
rect 392650 417218 392886 417454
rect 392650 416898 392886 417134
rect 423370 417218 423606 417454
rect 423370 416898 423606 417134
rect 454090 417218 454326 417454
rect 454090 416898 454326 417134
rect 484810 417218 485046 417454
rect 484810 416898 485046 417134
rect 515530 417218 515766 417454
rect 515530 416898 515766 417134
rect 546250 417218 546486 417454
rect 546250 416898 546486 417134
rect 576970 417218 577206 417454
rect 576970 416898 577206 417134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect 8650 399218 8886 399454
rect 8650 398898 8886 399134
rect 39370 399218 39606 399454
rect 39370 398898 39606 399134
rect 70090 399218 70326 399454
rect 70090 398898 70326 399134
rect 100810 399218 101046 399454
rect 100810 398898 101046 399134
rect 131530 399218 131766 399454
rect 131530 398898 131766 399134
rect 162250 399218 162486 399454
rect 162250 398898 162486 399134
rect 192970 399218 193206 399454
rect 192970 398898 193206 399134
rect 223690 399218 223926 399454
rect 223690 398898 223926 399134
rect 254410 399218 254646 399454
rect 254410 398898 254646 399134
rect 285130 399218 285366 399454
rect 285130 398898 285366 399134
rect 315850 399218 316086 399454
rect 315850 398898 316086 399134
rect 346570 399218 346806 399454
rect 346570 398898 346806 399134
rect 377290 399218 377526 399454
rect 377290 398898 377526 399134
rect 408010 399218 408246 399454
rect 408010 398898 408246 399134
rect 438730 399218 438966 399454
rect 438730 398898 438966 399134
rect 469450 399218 469686 399454
rect 469450 398898 469686 399134
rect 500170 399218 500406 399454
rect 500170 398898 500406 399134
rect 530890 399218 531126 399454
rect 530890 398898 531126 399134
rect 561610 399218 561846 399454
rect 561610 398898 561846 399134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 24010 381218 24246 381454
rect 24010 380898 24246 381134
rect 54730 381218 54966 381454
rect 54730 380898 54966 381134
rect 85450 381218 85686 381454
rect 85450 380898 85686 381134
rect 116170 381218 116406 381454
rect 116170 380898 116406 381134
rect 146890 381218 147126 381454
rect 146890 380898 147126 381134
rect 177610 381218 177846 381454
rect 177610 380898 177846 381134
rect 208330 381218 208566 381454
rect 208330 380898 208566 381134
rect 239050 381218 239286 381454
rect 239050 380898 239286 381134
rect 269770 381218 270006 381454
rect 269770 380898 270006 381134
rect 300490 381218 300726 381454
rect 300490 380898 300726 381134
rect 331210 381218 331446 381454
rect 331210 380898 331446 381134
rect 361930 381218 362166 381454
rect 361930 380898 362166 381134
rect 392650 381218 392886 381454
rect 392650 380898 392886 381134
rect 423370 381218 423606 381454
rect 423370 380898 423606 381134
rect 454090 381218 454326 381454
rect 454090 380898 454326 381134
rect 484810 381218 485046 381454
rect 484810 380898 485046 381134
rect 515530 381218 515766 381454
rect 515530 380898 515766 381134
rect 546250 381218 546486 381454
rect 546250 380898 546486 381134
rect 576970 381218 577206 381454
rect 576970 380898 577206 381134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect 8650 363218 8886 363454
rect 8650 362898 8886 363134
rect 39370 363218 39606 363454
rect 39370 362898 39606 363134
rect 70090 363218 70326 363454
rect 70090 362898 70326 363134
rect 100810 363218 101046 363454
rect 100810 362898 101046 363134
rect 131530 363218 131766 363454
rect 131530 362898 131766 363134
rect 162250 363218 162486 363454
rect 162250 362898 162486 363134
rect 192970 363218 193206 363454
rect 192970 362898 193206 363134
rect 223690 363218 223926 363454
rect 223690 362898 223926 363134
rect 254410 363218 254646 363454
rect 254410 362898 254646 363134
rect 285130 363218 285366 363454
rect 285130 362898 285366 363134
rect 315850 363218 316086 363454
rect 315850 362898 316086 363134
rect 346570 363218 346806 363454
rect 346570 362898 346806 363134
rect 377290 363218 377526 363454
rect 377290 362898 377526 363134
rect 408010 363218 408246 363454
rect 408010 362898 408246 363134
rect 438730 363218 438966 363454
rect 438730 362898 438966 363134
rect 469450 363218 469686 363454
rect 469450 362898 469686 363134
rect 500170 363218 500406 363454
rect 500170 362898 500406 363134
rect 530890 363218 531126 363454
rect 530890 362898 531126 363134
rect 561610 363218 561846 363454
rect 561610 362898 561846 363134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 24010 345218 24246 345454
rect 24010 344898 24246 345134
rect 54730 345218 54966 345454
rect 54730 344898 54966 345134
rect 85450 345218 85686 345454
rect 85450 344898 85686 345134
rect 116170 345218 116406 345454
rect 116170 344898 116406 345134
rect 146890 345218 147126 345454
rect 146890 344898 147126 345134
rect 177610 345218 177846 345454
rect 177610 344898 177846 345134
rect 208330 345218 208566 345454
rect 208330 344898 208566 345134
rect 239050 345218 239286 345454
rect 239050 344898 239286 345134
rect 269770 345218 270006 345454
rect 269770 344898 270006 345134
rect 300490 345218 300726 345454
rect 300490 344898 300726 345134
rect 331210 345218 331446 345454
rect 331210 344898 331446 345134
rect 361930 345218 362166 345454
rect 361930 344898 362166 345134
rect 392650 345218 392886 345454
rect 392650 344898 392886 345134
rect 423370 345218 423606 345454
rect 423370 344898 423606 345134
rect 454090 345218 454326 345454
rect 454090 344898 454326 345134
rect 484810 345218 485046 345454
rect 484810 344898 485046 345134
rect 515530 345218 515766 345454
rect 515530 344898 515766 345134
rect 546250 345218 546486 345454
rect 546250 344898 546486 345134
rect 576970 345218 577206 345454
rect 576970 344898 577206 345134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect 8650 327218 8886 327454
rect 8650 326898 8886 327134
rect 39370 327218 39606 327454
rect 39370 326898 39606 327134
rect 70090 327218 70326 327454
rect 70090 326898 70326 327134
rect 100810 327218 101046 327454
rect 100810 326898 101046 327134
rect 131530 327218 131766 327454
rect 131530 326898 131766 327134
rect 162250 327218 162486 327454
rect 162250 326898 162486 327134
rect 192970 327218 193206 327454
rect 192970 326898 193206 327134
rect 223690 327218 223926 327454
rect 223690 326898 223926 327134
rect 254410 327218 254646 327454
rect 254410 326898 254646 327134
rect 285130 327218 285366 327454
rect 285130 326898 285366 327134
rect 315850 327218 316086 327454
rect 315850 326898 316086 327134
rect 346570 327218 346806 327454
rect 346570 326898 346806 327134
rect 377290 327218 377526 327454
rect 377290 326898 377526 327134
rect 408010 327218 408246 327454
rect 408010 326898 408246 327134
rect 438730 327218 438966 327454
rect 438730 326898 438966 327134
rect 469450 327218 469686 327454
rect 469450 326898 469686 327134
rect 500170 327218 500406 327454
rect 500170 326898 500406 327134
rect 530890 327218 531126 327454
rect 530890 326898 531126 327134
rect 561610 327218 561846 327454
rect 561610 326898 561846 327134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 24010 309218 24246 309454
rect 24010 308898 24246 309134
rect 54730 309218 54966 309454
rect 54730 308898 54966 309134
rect 85450 309218 85686 309454
rect 85450 308898 85686 309134
rect 116170 309218 116406 309454
rect 116170 308898 116406 309134
rect 146890 309218 147126 309454
rect 146890 308898 147126 309134
rect 177610 309218 177846 309454
rect 177610 308898 177846 309134
rect 208330 309218 208566 309454
rect 208330 308898 208566 309134
rect 239050 309218 239286 309454
rect 239050 308898 239286 309134
rect 269770 309218 270006 309454
rect 269770 308898 270006 309134
rect 300490 309218 300726 309454
rect 300490 308898 300726 309134
rect 331210 309218 331446 309454
rect 331210 308898 331446 309134
rect 361930 309218 362166 309454
rect 361930 308898 362166 309134
rect 392650 309218 392886 309454
rect 392650 308898 392886 309134
rect 423370 309218 423606 309454
rect 423370 308898 423606 309134
rect 454090 309218 454326 309454
rect 454090 308898 454326 309134
rect 484810 309218 485046 309454
rect 484810 308898 485046 309134
rect 515530 309218 515766 309454
rect 515530 308898 515766 309134
rect 546250 309218 546486 309454
rect 546250 308898 546486 309134
rect 576970 309218 577206 309454
rect 576970 308898 577206 309134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect 8650 291218 8886 291454
rect 8650 290898 8886 291134
rect 39370 291218 39606 291454
rect 39370 290898 39606 291134
rect 70090 291218 70326 291454
rect 70090 290898 70326 291134
rect 100810 291218 101046 291454
rect 100810 290898 101046 291134
rect 131530 291218 131766 291454
rect 131530 290898 131766 291134
rect 162250 291218 162486 291454
rect 162250 290898 162486 291134
rect 192970 291218 193206 291454
rect 192970 290898 193206 291134
rect 223690 291218 223926 291454
rect 223690 290898 223926 291134
rect 254410 291218 254646 291454
rect 254410 290898 254646 291134
rect 285130 291218 285366 291454
rect 285130 290898 285366 291134
rect 315850 291218 316086 291454
rect 315850 290898 316086 291134
rect 346570 291218 346806 291454
rect 346570 290898 346806 291134
rect 377290 291218 377526 291454
rect 377290 290898 377526 291134
rect 408010 291218 408246 291454
rect 408010 290898 408246 291134
rect 438730 291218 438966 291454
rect 438730 290898 438966 291134
rect 469450 291218 469686 291454
rect 469450 290898 469686 291134
rect 500170 291218 500406 291454
rect 500170 290898 500406 291134
rect 530890 291218 531126 291454
rect 530890 290898 531126 291134
rect 561610 291218 561846 291454
rect 561610 290898 561846 291134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 24010 273218 24246 273454
rect 24010 272898 24246 273134
rect 54730 273218 54966 273454
rect 54730 272898 54966 273134
rect 85450 273218 85686 273454
rect 85450 272898 85686 273134
rect 116170 273218 116406 273454
rect 116170 272898 116406 273134
rect 146890 273218 147126 273454
rect 146890 272898 147126 273134
rect 177610 273218 177846 273454
rect 177610 272898 177846 273134
rect 208330 273218 208566 273454
rect 208330 272898 208566 273134
rect 239050 273218 239286 273454
rect 239050 272898 239286 273134
rect 269770 273218 270006 273454
rect 269770 272898 270006 273134
rect 300490 273218 300726 273454
rect 300490 272898 300726 273134
rect 331210 273218 331446 273454
rect 331210 272898 331446 273134
rect 361930 273218 362166 273454
rect 361930 272898 362166 273134
rect 392650 273218 392886 273454
rect 392650 272898 392886 273134
rect 423370 273218 423606 273454
rect 423370 272898 423606 273134
rect 454090 273218 454326 273454
rect 454090 272898 454326 273134
rect 484810 273218 485046 273454
rect 484810 272898 485046 273134
rect 515530 273218 515766 273454
rect 515530 272898 515766 273134
rect 546250 273218 546486 273454
rect 546250 272898 546486 273134
rect 576970 273218 577206 273454
rect 576970 272898 577206 273134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect 8650 255218 8886 255454
rect 8650 254898 8886 255134
rect 39370 255218 39606 255454
rect 39370 254898 39606 255134
rect 70090 255218 70326 255454
rect 70090 254898 70326 255134
rect 100810 255218 101046 255454
rect 100810 254898 101046 255134
rect 131530 255218 131766 255454
rect 131530 254898 131766 255134
rect 162250 255218 162486 255454
rect 162250 254898 162486 255134
rect 192970 255218 193206 255454
rect 192970 254898 193206 255134
rect 223690 255218 223926 255454
rect 223690 254898 223926 255134
rect 254410 255218 254646 255454
rect 254410 254898 254646 255134
rect 285130 255218 285366 255454
rect 285130 254898 285366 255134
rect 315850 255218 316086 255454
rect 315850 254898 316086 255134
rect 346570 255218 346806 255454
rect 346570 254898 346806 255134
rect 377290 255218 377526 255454
rect 377290 254898 377526 255134
rect 408010 255218 408246 255454
rect 408010 254898 408246 255134
rect 438730 255218 438966 255454
rect 438730 254898 438966 255134
rect 469450 255218 469686 255454
rect 469450 254898 469686 255134
rect 500170 255218 500406 255454
rect 500170 254898 500406 255134
rect 530890 255218 531126 255454
rect 530890 254898 531126 255134
rect 561610 255218 561846 255454
rect 561610 254898 561846 255134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 24010 237218 24246 237454
rect 24010 236898 24246 237134
rect 54730 237218 54966 237454
rect 54730 236898 54966 237134
rect 85450 237218 85686 237454
rect 85450 236898 85686 237134
rect 116170 237218 116406 237454
rect 116170 236898 116406 237134
rect 146890 237218 147126 237454
rect 146890 236898 147126 237134
rect 177610 237218 177846 237454
rect 177610 236898 177846 237134
rect 208330 237218 208566 237454
rect 208330 236898 208566 237134
rect 239050 237218 239286 237454
rect 239050 236898 239286 237134
rect 269770 237218 270006 237454
rect 269770 236898 270006 237134
rect 300490 237218 300726 237454
rect 300490 236898 300726 237134
rect 331210 237218 331446 237454
rect 331210 236898 331446 237134
rect 361930 237218 362166 237454
rect 361930 236898 362166 237134
rect 392650 237218 392886 237454
rect 392650 236898 392886 237134
rect 423370 237218 423606 237454
rect 423370 236898 423606 237134
rect 454090 237218 454326 237454
rect 454090 236898 454326 237134
rect 484810 237218 485046 237454
rect 484810 236898 485046 237134
rect 515530 237218 515766 237454
rect 515530 236898 515766 237134
rect 546250 237218 546486 237454
rect 546250 236898 546486 237134
rect 576970 237218 577206 237454
rect 576970 236898 577206 237134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect 8650 219218 8886 219454
rect 8650 218898 8886 219134
rect 39370 219218 39606 219454
rect 39370 218898 39606 219134
rect 70090 219218 70326 219454
rect 70090 218898 70326 219134
rect 100810 219218 101046 219454
rect 100810 218898 101046 219134
rect 131530 219218 131766 219454
rect 131530 218898 131766 219134
rect 162250 219218 162486 219454
rect 162250 218898 162486 219134
rect 192970 219218 193206 219454
rect 192970 218898 193206 219134
rect 223690 219218 223926 219454
rect 223690 218898 223926 219134
rect 254410 219218 254646 219454
rect 254410 218898 254646 219134
rect 285130 219218 285366 219454
rect 285130 218898 285366 219134
rect 315850 219218 316086 219454
rect 315850 218898 316086 219134
rect 346570 219218 346806 219454
rect 346570 218898 346806 219134
rect 377290 219218 377526 219454
rect 377290 218898 377526 219134
rect 408010 219218 408246 219454
rect 408010 218898 408246 219134
rect 438730 219218 438966 219454
rect 438730 218898 438966 219134
rect 469450 219218 469686 219454
rect 469450 218898 469686 219134
rect 500170 219218 500406 219454
rect 500170 218898 500406 219134
rect 530890 219218 531126 219454
rect 530890 218898 531126 219134
rect 561610 219218 561846 219454
rect 561610 218898 561846 219134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 24010 201218 24246 201454
rect 24010 200898 24246 201134
rect 54730 201218 54966 201454
rect 54730 200898 54966 201134
rect 85450 201218 85686 201454
rect 85450 200898 85686 201134
rect 116170 201218 116406 201454
rect 116170 200898 116406 201134
rect 146890 201218 147126 201454
rect 146890 200898 147126 201134
rect 177610 201218 177846 201454
rect 177610 200898 177846 201134
rect 208330 201218 208566 201454
rect 208330 200898 208566 201134
rect 239050 201218 239286 201454
rect 239050 200898 239286 201134
rect 269770 201218 270006 201454
rect 269770 200898 270006 201134
rect 300490 201218 300726 201454
rect 300490 200898 300726 201134
rect 331210 201218 331446 201454
rect 331210 200898 331446 201134
rect 361930 201218 362166 201454
rect 361930 200898 362166 201134
rect 392650 201218 392886 201454
rect 392650 200898 392886 201134
rect 423370 201218 423606 201454
rect 423370 200898 423606 201134
rect 454090 201218 454326 201454
rect 454090 200898 454326 201134
rect 484810 201218 485046 201454
rect 484810 200898 485046 201134
rect 515530 201218 515766 201454
rect 515530 200898 515766 201134
rect 546250 201218 546486 201454
rect 546250 200898 546486 201134
rect 576970 201218 577206 201454
rect 576970 200898 577206 201134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect 8650 183218 8886 183454
rect 8650 182898 8886 183134
rect 39370 183218 39606 183454
rect 39370 182898 39606 183134
rect 70090 183218 70326 183454
rect 70090 182898 70326 183134
rect 100810 183218 101046 183454
rect 100810 182898 101046 183134
rect 131530 183218 131766 183454
rect 131530 182898 131766 183134
rect 162250 183218 162486 183454
rect 162250 182898 162486 183134
rect 192970 183218 193206 183454
rect 192970 182898 193206 183134
rect 223690 183218 223926 183454
rect 223690 182898 223926 183134
rect 254410 183218 254646 183454
rect 254410 182898 254646 183134
rect 285130 183218 285366 183454
rect 285130 182898 285366 183134
rect 315850 183218 316086 183454
rect 315850 182898 316086 183134
rect 346570 183218 346806 183454
rect 346570 182898 346806 183134
rect 377290 183218 377526 183454
rect 377290 182898 377526 183134
rect 408010 183218 408246 183454
rect 408010 182898 408246 183134
rect 438730 183218 438966 183454
rect 438730 182898 438966 183134
rect 469450 183218 469686 183454
rect 469450 182898 469686 183134
rect 500170 183218 500406 183454
rect 500170 182898 500406 183134
rect 530890 183218 531126 183454
rect 530890 182898 531126 183134
rect 561610 183218 561846 183454
rect 561610 182898 561846 183134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 24010 165218 24246 165454
rect 24010 164898 24246 165134
rect 54730 165218 54966 165454
rect 54730 164898 54966 165134
rect 85450 165218 85686 165454
rect 85450 164898 85686 165134
rect 116170 165218 116406 165454
rect 116170 164898 116406 165134
rect 146890 165218 147126 165454
rect 146890 164898 147126 165134
rect 177610 165218 177846 165454
rect 177610 164898 177846 165134
rect 208330 165218 208566 165454
rect 208330 164898 208566 165134
rect 239050 165218 239286 165454
rect 239050 164898 239286 165134
rect 269770 165218 270006 165454
rect 269770 164898 270006 165134
rect 300490 165218 300726 165454
rect 300490 164898 300726 165134
rect 331210 165218 331446 165454
rect 331210 164898 331446 165134
rect 361930 165218 362166 165454
rect 361930 164898 362166 165134
rect 392650 165218 392886 165454
rect 392650 164898 392886 165134
rect 423370 165218 423606 165454
rect 423370 164898 423606 165134
rect 454090 165218 454326 165454
rect 454090 164898 454326 165134
rect 484810 165218 485046 165454
rect 484810 164898 485046 165134
rect 515530 165218 515766 165454
rect 515530 164898 515766 165134
rect 546250 165218 546486 165454
rect 546250 164898 546486 165134
rect 576970 165218 577206 165454
rect 576970 164898 577206 165134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect 8650 147218 8886 147454
rect 8650 146898 8886 147134
rect 39370 147218 39606 147454
rect 39370 146898 39606 147134
rect 70090 147218 70326 147454
rect 70090 146898 70326 147134
rect 100810 147218 101046 147454
rect 100810 146898 101046 147134
rect 131530 147218 131766 147454
rect 131530 146898 131766 147134
rect 162250 147218 162486 147454
rect 162250 146898 162486 147134
rect 192970 147218 193206 147454
rect 192970 146898 193206 147134
rect 223690 147218 223926 147454
rect 223690 146898 223926 147134
rect 254410 147218 254646 147454
rect 254410 146898 254646 147134
rect 285130 147218 285366 147454
rect 285130 146898 285366 147134
rect 315850 147218 316086 147454
rect 315850 146898 316086 147134
rect 346570 147218 346806 147454
rect 346570 146898 346806 147134
rect 377290 147218 377526 147454
rect 377290 146898 377526 147134
rect 408010 147218 408246 147454
rect 408010 146898 408246 147134
rect 438730 147218 438966 147454
rect 438730 146898 438966 147134
rect 469450 147218 469686 147454
rect 469450 146898 469686 147134
rect 500170 147218 500406 147454
rect 500170 146898 500406 147134
rect 530890 147218 531126 147454
rect 530890 146898 531126 147134
rect 561610 147218 561846 147454
rect 561610 146898 561846 147134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 24010 129218 24246 129454
rect 24010 128898 24246 129134
rect 54730 129218 54966 129454
rect 54730 128898 54966 129134
rect 85450 129218 85686 129454
rect 85450 128898 85686 129134
rect 116170 129218 116406 129454
rect 116170 128898 116406 129134
rect 146890 129218 147126 129454
rect 146890 128898 147126 129134
rect 177610 129218 177846 129454
rect 177610 128898 177846 129134
rect 208330 129218 208566 129454
rect 208330 128898 208566 129134
rect 239050 129218 239286 129454
rect 239050 128898 239286 129134
rect 269770 129218 270006 129454
rect 269770 128898 270006 129134
rect 300490 129218 300726 129454
rect 300490 128898 300726 129134
rect 331210 129218 331446 129454
rect 331210 128898 331446 129134
rect 361930 129218 362166 129454
rect 361930 128898 362166 129134
rect 392650 129218 392886 129454
rect 392650 128898 392886 129134
rect 423370 129218 423606 129454
rect 423370 128898 423606 129134
rect 454090 129218 454326 129454
rect 454090 128898 454326 129134
rect 484810 129218 485046 129454
rect 484810 128898 485046 129134
rect 515530 129218 515766 129454
rect 515530 128898 515766 129134
rect 546250 129218 546486 129454
rect 546250 128898 546486 129134
rect 576970 129218 577206 129454
rect 576970 128898 577206 129134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect 8650 111218 8886 111454
rect 8650 110898 8886 111134
rect 39370 111218 39606 111454
rect 39370 110898 39606 111134
rect 70090 111218 70326 111454
rect 70090 110898 70326 111134
rect 100810 111218 101046 111454
rect 100810 110898 101046 111134
rect 131530 111218 131766 111454
rect 131530 110898 131766 111134
rect 162250 111218 162486 111454
rect 162250 110898 162486 111134
rect 192970 111218 193206 111454
rect 192970 110898 193206 111134
rect 223690 111218 223926 111454
rect 223690 110898 223926 111134
rect 254410 111218 254646 111454
rect 254410 110898 254646 111134
rect 285130 111218 285366 111454
rect 285130 110898 285366 111134
rect 315850 111218 316086 111454
rect 315850 110898 316086 111134
rect 346570 111218 346806 111454
rect 346570 110898 346806 111134
rect 377290 111218 377526 111454
rect 377290 110898 377526 111134
rect 408010 111218 408246 111454
rect 408010 110898 408246 111134
rect 438730 111218 438966 111454
rect 438730 110898 438966 111134
rect 469450 111218 469686 111454
rect 469450 110898 469686 111134
rect 500170 111218 500406 111454
rect 500170 110898 500406 111134
rect 530890 111218 531126 111454
rect 530890 110898 531126 111134
rect 561610 111218 561846 111454
rect 561610 110898 561846 111134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 24010 93218 24246 93454
rect 24010 92898 24246 93134
rect 54730 93218 54966 93454
rect 54730 92898 54966 93134
rect 85450 93218 85686 93454
rect 85450 92898 85686 93134
rect 116170 93218 116406 93454
rect 116170 92898 116406 93134
rect 146890 93218 147126 93454
rect 146890 92898 147126 93134
rect 177610 93218 177846 93454
rect 177610 92898 177846 93134
rect 208330 93218 208566 93454
rect 208330 92898 208566 93134
rect 239050 93218 239286 93454
rect 239050 92898 239286 93134
rect 269770 93218 270006 93454
rect 269770 92898 270006 93134
rect 300490 93218 300726 93454
rect 300490 92898 300726 93134
rect 331210 93218 331446 93454
rect 331210 92898 331446 93134
rect 361930 93218 362166 93454
rect 361930 92898 362166 93134
rect 392650 93218 392886 93454
rect 392650 92898 392886 93134
rect 423370 93218 423606 93454
rect 423370 92898 423606 93134
rect 454090 93218 454326 93454
rect 454090 92898 454326 93134
rect 484810 93218 485046 93454
rect 484810 92898 485046 93134
rect 515530 93218 515766 93454
rect 515530 92898 515766 93134
rect 546250 93218 546486 93454
rect 546250 92898 546486 93134
rect 576970 93218 577206 93454
rect 576970 92898 577206 93134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect 8650 75218 8886 75454
rect 8650 74898 8886 75134
rect 39370 75218 39606 75454
rect 39370 74898 39606 75134
rect 70090 75218 70326 75454
rect 70090 74898 70326 75134
rect 100810 75218 101046 75454
rect 100810 74898 101046 75134
rect 131530 75218 131766 75454
rect 131530 74898 131766 75134
rect 162250 75218 162486 75454
rect 162250 74898 162486 75134
rect 192970 75218 193206 75454
rect 192970 74898 193206 75134
rect 223690 75218 223926 75454
rect 223690 74898 223926 75134
rect 254410 75218 254646 75454
rect 254410 74898 254646 75134
rect 285130 75218 285366 75454
rect 285130 74898 285366 75134
rect 315850 75218 316086 75454
rect 315850 74898 316086 75134
rect 346570 75218 346806 75454
rect 346570 74898 346806 75134
rect 377290 75218 377526 75454
rect 377290 74898 377526 75134
rect 408010 75218 408246 75454
rect 408010 74898 408246 75134
rect 438730 75218 438966 75454
rect 438730 74898 438966 75134
rect 469450 75218 469686 75454
rect 469450 74898 469686 75134
rect 500170 75218 500406 75454
rect 500170 74898 500406 75134
rect 530890 75218 531126 75454
rect 530890 74898 531126 75134
rect 561610 75218 561846 75454
rect 561610 74898 561846 75134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 24010 57218 24246 57454
rect 24010 56898 24246 57134
rect 54730 57218 54966 57454
rect 54730 56898 54966 57134
rect 85450 57218 85686 57454
rect 85450 56898 85686 57134
rect 116170 57218 116406 57454
rect 116170 56898 116406 57134
rect 146890 57218 147126 57454
rect 146890 56898 147126 57134
rect 177610 57218 177846 57454
rect 177610 56898 177846 57134
rect 208330 57218 208566 57454
rect 208330 56898 208566 57134
rect 239050 57218 239286 57454
rect 239050 56898 239286 57134
rect 269770 57218 270006 57454
rect 269770 56898 270006 57134
rect 300490 57218 300726 57454
rect 300490 56898 300726 57134
rect 331210 57218 331446 57454
rect 331210 56898 331446 57134
rect 361930 57218 362166 57454
rect 361930 56898 362166 57134
rect 392650 57218 392886 57454
rect 392650 56898 392886 57134
rect 423370 57218 423606 57454
rect 423370 56898 423606 57134
rect 454090 57218 454326 57454
rect 454090 56898 454326 57134
rect 484810 57218 485046 57454
rect 484810 56898 485046 57134
rect 515530 57218 515766 57454
rect 515530 56898 515766 57134
rect 546250 57218 546486 57454
rect 546250 56898 546486 57134
rect 576970 57218 577206 57454
rect 576970 56898 577206 57134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect 8650 39218 8886 39454
rect 8650 38898 8886 39134
rect 39370 39218 39606 39454
rect 39370 38898 39606 39134
rect 70090 39218 70326 39454
rect 70090 38898 70326 39134
rect 100810 39218 101046 39454
rect 100810 38898 101046 39134
rect 131530 39218 131766 39454
rect 131530 38898 131766 39134
rect 162250 39218 162486 39454
rect 162250 38898 162486 39134
rect 192970 39218 193206 39454
rect 192970 38898 193206 39134
rect 223690 39218 223926 39454
rect 223690 38898 223926 39134
rect 254410 39218 254646 39454
rect 254410 38898 254646 39134
rect 285130 39218 285366 39454
rect 285130 38898 285366 39134
rect 315850 39218 316086 39454
rect 315850 38898 316086 39134
rect 346570 39218 346806 39454
rect 346570 38898 346806 39134
rect 377290 39218 377526 39454
rect 377290 38898 377526 39134
rect 408010 39218 408246 39454
rect 408010 38898 408246 39134
rect 438730 39218 438966 39454
rect 438730 38898 438966 39134
rect 469450 39218 469686 39454
rect 469450 38898 469686 39134
rect 500170 39218 500406 39454
rect 500170 38898 500406 39134
rect 530890 39218 531126 39454
rect 530890 38898 531126 39134
rect 561610 39218 561846 39454
rect 561610 38898 561846 39134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 24010 21218 24246 21454
rect 24010 20898 24246 21134
rect 54730 21218 54966 21454
rect 54730 20898 54966 21134
rect 85450 21218 85686 21454
rect 85450 20898 85686 21134
rect 116170 21218 116406 21454
rect 116170 20898 116406 21134
rect 146890 21218 147126 21454
rect 146890 20898 147126 21134
rect 177610 21218 177846 21454
rect 177610 20898 177846 21134
rect 208330 21218 208566 21454
rect 208330 20898 208566 21134
rect 239050 21218 239286 21454
rect 239050 20898 239286 21134
rect 269770 21218 270006 21454
rect 269770 20898 270006 21134
rect 300490 21218 300726 21454
rect 300490 20898 300726 21134
rect 331210 21218 331446 21454
rect 331210 20898 331446 21134
rect 361930 21218 362166 21454
rect 361930 20898 362166 21134
rect 392650 21218 392886 21454
rect 392650 20898 392886 21134
rect 423370 21218 423606 21454
rect 423370 20898 423606 21134
rect 454090 21218 454326 21454
rect 454090 20898 454326 21134
rect 484810 21218 485046 21454
rect 484810 20898 485046 21134
rect 515530 21218 515766 21454
rect 515530 20898 515766 21134
rect 546250 21218 546486 21454
rect 546250 20898 546486 21134
rect 576970 21218 577206 21454
rect 576970 20898 577206 21134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 8650 687454
rect 8886 687218 39370 687454
rect 39606 687218 70090 687454
rect 70326 687218 100810 687454
rect 101046 687218 131530 687454
rect 131766 687218 162250 687454
rect 162486 687218 192970 687454
rect 193206 687218 223690 687454
rect 223926 687218 254410 687454
rect 254646 687218 285130 687454
rect 285366 687218 315850 687454
rect 316086 687218 346570 687454
rect 346806 687218 377290 687454
rect 377526 687218 408010 687454
rect 408246 687218 438730 687454
rect 438966 687218 469450 687454
rect 469686 687218 500170 687454
rect 500406 687218 530890 687454
rect 531126 687218 561610 687454
rect 561846 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 8650 687134
rect 8886 686898 39370 687134
rect 39606 686898 70090 687134
rect 70326 686898 100810 687134
rect 101046 686898 131530 687134
rect 131766 686898 162250 687134
rect 162486 686898 192970 687134
rect 193206 686898 223690 687134
rect 223926 686898 254410 687134
rect 254646 686898 285130 687134
rect 285366 686898 315850 687134
rect 316086 686898 346570 687134
rect 346806 686898 377290 687134
rect 377526 686898 408010 687134
rect 408246 686898 438730 687134
rect 438966 686898 469450 687134
rect 469686 686898 500170 687134
rect 500406 686898 530890 687134
rect 531126 686898 561610 687134
rect 561846 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 24010 669454
rect 24246 669218 54730 669454
rect 54966 669218 85450 669454
rect 85686 669218 116170 669454
rect 116406 669218 146890 669454
rect 147126 669218 177610 669454
rect 177846 669218 208330 669454
rect 208566 669218 239050 669454
rect 239286 669218 269770 669454
rect 270006 669218 300490 669454
rect 300726 669218 331210 669454
rect 331446 669218 361930 669454
rect 362166 669218 392650 669454
rect 392886 669218 423370 669454
rect 423606 669218 454090 669454
rect 454326 669218 484810 669454
rect 485046 669218 515530 669454
rect 515766 669218 546250 669454
rect 546486 669218 576970 669454
rect 577206 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 24010 669134
rect 24246 668898 54730 669134
rect 54966 668898 85450 669134
rect 85686 668898 116170 669134
rect 116406 668898 146890 669134
rect 147126 668898 177610 669134
rect 177846 668898 208330 669134
rect 208566 668898 239050 669134
rect 239286 668898 269770 669134
rect 270006 668898 300490 669134
rect 300726 668898 331210 669134
rect 331446 668898 361930 669134
rect 362166 668898 392650 669134
rect 392886 668898 423370 669134
rect 423606 668898 454090 669134
rect 454326 668898 484810 669134
rect 485046 668898 515530 669134
rect 515766 668898 546250 669134
rect 546486 668898 576970 669134
rect 577206 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 8650 651454
rect 8886 651218 39370 651454
rect 39606 651218 70090 651454
rect 70326 651218 100810 651454
rect 101046 651218 131530 651454
rect 131766 651218 162250 651454
rect 162486 651218 192970 651454
rect 193206 651218 223690 651454
rect 223926 651218 254410 651454
rect 254646 651218 285130 651454
rect 285366 651218 315850 651454
rect 316086 651218 346570 651454
rect 346806 651218 377290 651454
rect 377526 651218 408010 651454
rect 408246 651218 438730 651454
rect 438966 651218 469450 651454
rect 469686 651218 500170 651454
rect 500406 651218 530890 651454
rect 531126 651218 561610 651454
rect 561846 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 8650 651134
rect 8886 650898 39370 651134
rect 39606 650898 70090 651134
rect 70326 650898 100810 651134
rect 101046 650898 131530 651134
rect 131766 650898 162250 651134
rect 162486 650898 192970 651134
rect 193206 650898 223690 651134
rect 223926 650898 254410 651134
rect 254646 650898 285130 651134
rect 285366 650898 315850 651134
rect 316086 650898 346570 651134
rect 346806 650898 377290 651134
rect 377526 650898 408010 651134
rect 408246 650898 438730 651134
rect 438966 650898 469450 651134
rect 469686 650898 500170 651134
rect 500406 650898 530890 651134
rect 531126 650898 561610 651134
rect 561846 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 24010 633454
rect 24246 633218 54730 633454
rect 54966 633218 85450 633454
rect 85686 633218 116170 633454
rect 116406 633218 146890 633454
rect 147126 633218 177610 633454
rect 177846 633218 208330 633454
rect 208566 633218 239050 633454
rect 239286 633218 269770 633454
rect 270006 633218 300490 633454
rect 300726 633218 331210 633454
rect 331446 633218 361930 633454
rect 362166 633218 392650 633454
rect 392886 633218 423370 633454
rect 423606 633218 454090 633454
rect 454326 633218 484810 633454
rect 485046 633218 515530 633454
rect 515766 633218 546250 633454
rect 546486 633218 576970 633454
rect 577206 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 24010 633134
rect 24246 632898 54730 633134
rect 54966 632898 85450 633134
rect 85686 632898 116170 633134
rect 116406 632898 146890 633134
rect 147126 632898 177610 633134
rect 177846 632898 208330 633134
rect 208566 632898 239050 633134
rect 239286 632898 269770 633134
rect 270006 632898 300490 633134
rect 300726 632898 331210 633134
rect 331446 632898 361930 633134
rect 362166 632898 392650 633134
rect 392886 632898 423370 633134
rect 423606 632898 454090 633134
rect 454326 632898 484810 633134
rect 485046 632898 515530 633134
rect 515766 632898 546250 633134
rect 546486 632898 576970 633134
rect 577206 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 8650 615454
rect 8886 615218 39370 615454
rect 39606 615218 70090 615454
rect 70326 615218 100810 615454
rect 101046 615218 131530 615454
rect 131766 615218 162250 615454
rect 162486 615218 192970 615454
rect 193206 615218 223690 615454
rect 223926 615218 254410 615454
rect 254646 615218 285130 615454
rect 285366 615218 315850 615454
rect 316086 615218 346570 615454
rect 346806 615218 377290 615454
rect 377526 615218 408010 615454
rect 408246 615218 438730 615454
rect 438966 615218 469450 615454
rect 469686 615218 500170 615454
rect 500406 615218 530890 615454
rect 531126 615218 561610 615454
rect 561846 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 8650 615134
rect 8886 614898 39370 615134
rect 39606 614898 70090 615134
rect 70326 614898 100810 615134
rect 101046 614898 131530 615134
rect 131766 614898 162250 615134
rect 162486 614898 192970 615134
rect 193206 614898 223690 615134
rect 223926 614898 254410 615134
rect 254646 614898 285130 615134
rect 285366 614898 315850 615134
rect 316086 614898 346570 615134
rect 346806 614898 377290 615134
rect 377526 614898 408010 615134
rect 408246 614898 438730 615134
rect 438966 614898 469450 615134
rect 469686 614898 500170 615134
rect 500406 614898 530890 615134
rect 531126 614898 561610 615134
rect 561846 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 24010 597454
rect 24246 597218 54730 597454
rect 54966 597218 85450 597454
rect 85686 597218 116170 597454
rect 116406 597218 146890 597454
rect 147126 597218 177610 597454
rect 177846 597218 208330 597454
rect 208566 597218 239050 597454
rect 239286 597218 269770 597454
rect 270006 597218 300490 597454
rect 300726 597218 331210 597454
rect 331446 597218 361930 597454
rect 362166 597218 392650 597454
rect 392886 597218 423370 597454
rect 423606 597218 454090 597454
rect 454326 597218 484810 597454
rect 485046 597218 515530 597454
rect 515766 597218 546250 597454
rect 546486 597218 576970 597454
rect 577206 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 24010 597134
rect 24246 596898 54730 597134
rect 54966 596898 85450 597134
rect 85686 596898 116170 597134
rect 116406 596898 146890 597134
rect 147126 596898 177610 597134
rect 177846 596898 208330 597134
rect 208566 596898 239050 597134
rect 239286 596898 269770 597134
rect 270006 596898 300490 597134
rect 300726 596898 331210 597134
rect 331446 596898 361930 597134
rect 362166 596898 392650 597134
rect 392886 596898 423370 597134
rect 423606 596898 454090 597134
rect 454326 596898 484810 597134
rect 485046 596898 515530 597134
rect 515766 596898 546250 597134
rect 546486 596898 576970 597134
rect 577206 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 8650 579454
rect 8886 579218 39370 579454
rect 39606 579218 70090 579454
rect 70326 579218 100810 579454
rect 101046 579218 131530 579454
rect 131766 579218 162250 579454
rect 162486 579218 192970 579454
rect 193206 579218 223690 579454
rect 223926 579218 254410 579454
rect 254646 579218 285130 579454
rect 285366 579218 315850 579454
rect 316086 579218 346570 579454
rect 346806 579218 377290 579454
rect 377526 579218 408010 579454
rect 408246 579218 438730 579454
rect 438966 579218 469450 579454
rect 469686 579218 500170 579454
rect 500406 579218 530890 579454
rect 531126 579218 561610 579454
rect 561846 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 8650 579134
rect 8886 578898 39370 579134
rect 39606 578898 70090 579134
rect 70326 578898 100810 579134
rect 101046 578898 131530 579134
rect 131766 578898 162250 579134
rect 162486 578898 192970 579134
rect 193206 578898 223690 579134
rect 223926 578898 254410 579134
rect 254646 578898 285130 579134
rect 285366 578898 315850 579134
rect 316086 578898 346570 579134
rect 346806 578898 377290 579134
rect 377526 578898 408010 579134
rect 408246 578898 438730 579134
rect 438966 578898 469450 579134
rect 469686 578898 500170 579134
rect 500406 578898 530890 579134
rect 531126 578898 561610 579134
rect 561846 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 24010 561454
rect 24246 561218 54730 561454
rect 54966 561218 85450 561454
rect 85686 561218 116170 561454
rect 116406 561218 146890 561454
rect 147126 561218 177610 561454
rect 177846 561218 208330 561454
rect 208566 561218 239050 561454
rect 239286 561218 269770 561454
rect 270006 561218 300490 561454
rect 300726 561218 331210 561454
rect 331446 561218 361930 561454
rect 362166 561218 392650 561454
rect 392886 561218 423370 561454
rect 423606 561218 454090 561454
rect 454326 561218 484810 561454
rect 485046 561218 515530 561454
rect 515766 561218 546250 561454
rect 546486 561218 576970 561454
rect 577206 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 24010 561134
rect 24246 560898 54730 561134
rect 54966 560898 85450 561134
rect 85686 560898 116170 561134
rect 116406 560898 146890 561134
rect 147126 560898 177610 561134
rect 177846 560898 208330 561134
rect 208566 560898 239050 561134
rect 239286 560898 269770 561134
rect 270006 560898 300490 561134
rect 300726 560898 331210 561134
rect 331446 560898 361930 561134
rect 362166 560898 392650 561134
rect 392886 560898 423370 561134
rect 423606 560898 454090 561134
rect 454326 560898 484810 561134
rect 485046 560898 515530 561134
rect 515766 560898 546250 561134
rect 546486 560898 576970 561134
rect 577206 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 8650 543454
rect 8886 543218 39370 543454
rect 39606 543218 70090 543454
rect 70326 543218 100810 543454
rect 101046 543218 131530 543454
rect 131766 543218 162250 543454
rect 162486 543218 192970 543454
rect 193206 543218 223690 543454
rect 223926 543218 254410 543454
rect 254646 543218 285130 543454
rect 285366 543218 315850 543454
rect 316086 543218 346570 543454
rect 346806 543218 377290 543454
rect 377526 543218 408010 543454
rect 408246 543218 438730 543454
rect 438966 543218 469450 543454
rect 469686 543218 500170 543454
rect 500406 543218 530890 543454
rect 531126 543218 561610 543454
rect 561846 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 8650 543134
rect 8886 542898 39370 543134
rect 39606 542898 70090 543134
rect 70326 542898 100810 543134
rect 101046 542898 131530 543134
rect 131766 542898 162250 543134
rect 162486 542898 192970 543134
rect 193206 542898 223690 543134
rect 223926 542898 254410 543134
rect 254646 542898 285130 543134
rect 285366 542898 315850 543134
rect 316086 542898 346570 543134
rect 346806 542898 377290 543134
rect 377526 542898 408010 543134
rect 408246 542898 438730 543134
rect 438966 542898 469450 543134
rect 469686 542898 500170 543134
rect 500406 542898 530890 543134
rect 531126 542898 561610 543134
rect 561846 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 24010 525454
rect 24246 525218 54730 525454
rect 54966 525218 85450 525454
rect 85686 525218 116170 525454
rect 116406 525218 146890 525454
rect 147126 525218 177610 525454
rect 177846 525218 208330 525454
rect 208566 525218 239050 525454
rect 239286 525218 269770 525454
rect 270006 525218 300490 525454
rect 300726 525218 331210 525454
rect 331446 525218 361930 525454
rect 362166 525218 392650 525454
rect 392886 525218 423370 525454
rect 423606 525218 454090 525454
rect 454326 525218 484810 525454
rect 485046 525218 515530 525454
rect 515766 525218 546250 525454
rect 546486 525218 576970 525454
rect 577206 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 24010 525134
rect 24246 524898 54730 525134
rect 54966 524898 85450 525134
rect 85686 524898 116170 525134
rect 116406 524898 146890 525134
rect 147126 524898 177610 525134
rect 177846 524898 208330 525134
rect 208566 524898 239050 525134
rect 239286 524898 269770 525134
rect 270006 524898 300490 525134
rect 300726 524898 331210 525134
rect 331446 524898 361930 525134
rect 362166 524898 392650 525134
rect 392886 524898 423370 525134
rect 423606 524898 454090 525134
rect 454326 524898 484810 525134
rect 485046 524898 515530 525134
rect 515766 524898 546250 525134
rect 546486 524898 576970 525134
rect 577206 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 8650 507454
rect 8886 507218 39370 507454
rect 39606 507218 70090 507454
rect 70326 507218 100810 507454
rect 101046 507218 131530 507454
rect 131766 507218 162250 507454
rect 162486 507218 192970 507454
rect 193206 507218 223690 507454
rect 223926 507218 254410 507454
rect 254646 507218 285130 507454
rect 285366 507218 315850 507454
rect 316086 507218 346570 507454
rect 346806 507218 377290 507454
rect 377526 507218 408010 507454
rect 408246 507218 438730 507454
rect 438966 507218 469450 507454
rect 469686 507218 500170 507454
rect 500406 507218 530890 507454
rect 531126 507218 561610 507454
rect 561846 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 8650 507134
rect 8886 506898 39370 507134
rect 39606 506898 70090 507134
rect 70326 506898 100810 507134
rect 101046 506898 131530 507134
rect 131766 506898 162250 507134
rect 162486 506898 192970 507134
rect 193206 506898 223690 507134
rect 223926 506898 254410 507134
rect 254646 506898 285130 507134
rect 285366 506898 315850 507134
rect 316086 506898 346570 507134
rect 346806 506898 377290 507134
rect 377526 506898 408010 507134
rect 408246 506898 438730 507134
rect 438966 506898 469450 507134
rect 469686 506898 500170 507134
rect 500406 506898 530890 507134
rect 531126 506898 561610 507134
rect 561846 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 24010 489454
rect 24246 489218 54730 489454
rect 54966 489218 85450 489454
rect 85686 489218 116170 489454
rect 116406 489218 146890 489454
rect 147126 489218 177610 489454
rect 177846 489218 208330 489454
rect 208566 489218 239050 489454
rect 239286 489218 269770 489454
rect 270006 489218 300490 489454
rect 300726 489218 331210 489454
rect 331446 489218 361930 489454
rect 362166 489218 392650 489454
rect 392886 489218 423370 489454
rect 423606 489218 454090 489454
rect 454326 489218 484810 489454
rect 485046 489218 515530 489454
rect 515766 489218 546250 489454
rect 546486 489218 576970 489454
rect 577206 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 24010 489134
rect 24246 488898 54730 489134
rect 54966 488898 85450 489134
rect 85686 488898 116170 489134
rect 116406 488898 146890 489134
rect 147126 488898 177610 489134
rect 177846 488898 208330 489134
rect 208566 488898 239050 489134
rect 239286 488898 269770 489134
rect 270006 488898 300490 489134
rect 300726 488898 331210 489134
rect 331446 488898 361930 489134
rect 362166 488898 392650 489134
rect 392886 488898 423370 489134
rect 423606 488898 454090 489134
rect 454326 488898 484810 489134
rect 485046 488898 515530 489134
rect 515766 488898 546250 489134
rect 546486 488898 576970 489134
rect 577206 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 8650 471454
rect 8886 471218 39370 471454
rect 39606 471218 70090 471454
rect 70326 471218 100810 471454
rect 101046 471218 131530 471454
rect 131766 471218 162250 471454
rect 162486 471218 192970 471454
rect 193206 471218 223690 471454
rect 223926 471218 254410 471454
rect 254646 471218 285130 471454
rect 285366 471218 315850 471454
rect 316086 471218 346570 471454
rect 346806 471218 377290 471454
rect 377526 471218 408010 471454
rect 408246 471218 438730 471454
rect 438966 471218 469450 471454
rect 469686 471218 500170 471454
rect 500406 471218 530890 471454
rect 531126 471218 561610 471454
rect 561846 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 8650 471134
rect 8886 470898 39370 471134
rect 39606 470898 70090 471134
rect 70326 470898 100810 471134
rect 101046 470898 131530 471134
rect 131766 470898 162250 471134
rect 162486 470898 192970 471134
rect 193206 470898 223690 471134
rect 223926 470898 254410 471134
rect 254646 470898 285130 471134
rect 285366 470898 315850 471134
rect 316086 470898 346570 471134
rect 346806 470898 377290 471134
rect 377526 470898 408010 471134
rect 408246 470898 438730 471134
rect 438966 470898 469450 471134
rect 469686 470898 500170 471134
rect 500406 470898 530890 471134
rect 531126 470898 561610 471134
rect 561846 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 24010 453454
rect 24246 453218 54730 453454
rect 54966 453218 85450 453454
rect 85686 453218 116170 453454
rect 116406 453218 146890 453454
rect 147126 453218 177610 453454
rect 177846 453218 208330 453454
rect 208566 453218 239050 453454
rect 239286 453218 269770 453454
rect 270006 453218 300490 453454
rect 300726 453218 331210 453454
rect 331446 453218 361930 453454
rect 362166 453218 392650 453454
rect 392886 453218 423370 453454
rect 423606 453218 454090 453454
rect 454326 453218 484810 453454
rect 485046 453218 515530 453454
rect 515766 453218 546250 453454
rect 546486 453218 576970 453454
rect 577206 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 24010 453134
rect 24246 452898 54730 453134
rect 54966 452898 85450 453134
rect 85686 452898 116170 453134
rect 116406 452898 146890 453134
rect 147126 452898 177610 453134
rect 177846 452898 208330 453134
rect 208566 452898 239050 453134
rect 239286 452898 269770 453134
rect 270006 452898 300490 453134
rect 300726 452898 331210 453134
rect 331446 452898 361930 453134
rect 362166 452898 392650 453134
rect 392886 452898 423370 453134
rect 423606 452898 454090 453134
rect 454326 452898 484810 453134
rect 485046 452898 515530 453134
rect 515766 452898 546250 453134
rect 546486 452898 576970 453134
rect 577206 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 8650 435454
rect 8886 435218 39370 435454
rect 39606 435218 70090 435454
rect 70326 435218 100810 435454
rect 101046 435218 131530 435454
rect 131766 435218 162250 435454
rect 162486 435218 192970 435454
rect 193206 435218 223690 435454
rect 223926 435218 254410 435454
rect 254646 435218 285130 435454
rect 285366 435218 315850 435454
rect 316086 435218 346570 435454
rect 346806 435218 377290 435454
rect 377526 435218 408010 435454
rect 408246 435218 438730 435454
rect 438966 435218 469450 435454
rect 469686 435218 500170 435454
rect 500406 435218 530890 435454
rect 531126 435218 561610 435454
rect 561846 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 8650 435134
rect 8886 434898 39370 435134
rect 39606 434898 70090 435134
rect 70326 434898 100810 435134
rect 101046 434898 131530 435134
rect 131766 434898 162250 435134
rect 162486 434898 192970 435134
rect 193206 434898 223690 435134
rect 223926 434898 254410 435134
rect 254646 434898 285130 435134
rect 285366 434898 315850 435134
rect 316086 434898 346570 435134
rect 346806 434898 377290 435134
rect 377526 434898 408010 435134
rect 408246 434898 438730 435134
rect 438966 434898 469450 435134
rect 469686 434898 500170 435134
rect 500406 434898 530890 435134
rect 531126 434898 561610 435134
rect 561846 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 24010 417454
rect 24246 417218 54730 417454
rect 54966 417218 85450 417454
rect 85686 417218 116170 417454
rect 116406 417218 146890 417454
rect 147126 417218 177610 417454
rect 177846 417218 208330 417454
rect 208566 417218 239050 417454
rect 239286 417218 269770 417454
rect 270006 417218 300490 417454
rect 300726 417218 331210 417454
rect 331446 417218 361930 417454
rect 362166 417218 392650 417454
rect 392886 417218 423370 417454
rect 423606 417218 454090 417454
rect 454326 417218 484810 417454
rect 485046 417218 515530 417454
rect 515766 417218 546250 417454
rect 546486 417218 576970 417454
rect 577206 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 24010 417134
rect 24246 416898 54730 417134
rect 54966 416898 85450 417134
rect 85686 416898 116170 417134
rect 116406 416898 146890 417134
rect 147126 416898 177610 417134
rect 177846 416898 208330 417134
rect 208566 416898 239050 417134
rect 239286 416898 269770 417134
rect 270006 416898 300490 417134
rect 300726 416898 331210 417134
rect 331446 416898 361930 417134
rect 362166 416898 392650 417134
rect 392886 416898 423370 417134
rect 423606 416898 454090 417134
rect 454326 416898 484810 417134
rect 485046 416898 515530 417134
rect 515766 416898 546250 417134
rect 546486 416898 576970 417134
rect 577206 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 8650 399454
rect 8886 399218 39370 399454
rect 39606 399218 70090 399454
rect 70326 399218 100810 399454
rect 101046 399218 131530 399454
rect 131766 399218 162250 399454
rect 162486 399218 192970 399454
rect 193206 399218 223690 399454
rect 223926 399218 254410 399454
rect 254646 399218 285130 399454
rect 285366 399218 315850 399454
rect 316086 399218 346570 399454
rect 346806 399218 377290 399454
rect 377526 399218 408010 399454
rect 408246 399218 438730 399454
rect 438966 399218 469450 399454
rect 469686 399218 500170 399454
rect 500406 399218 530890 399454
rect 531126 399218 561610 399454
rect 561846 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 8650 399134
rect 8886 398898 39370 399134
rect 39606 398898 70090 399134
rect 70326 398898 100810 399134
rect 101046 398898 131530 399134
rect 131766 398898 162250 399134
rect 162486 398898 192970 399134
rect 193206 398898 223690 399134
rect 223926 398898 254410 399134
rect 254646 398898 285130 399134
rect 285366 398898 315850 399134
rect 316086 398898 346570 399134
rect 346806 398898 377290 399134
rect 377526 398898 408010 399134
rect 408246 398898 438730 399134
rect 438966 398898 469450 399134
rect 469686 398898 500170 399134
rect 500406 398898 530890 399134
rect 531126 398898 561610 399134
rect 561846 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 24010 381454
rect 24246 381218 54730 381454
rect 54966 381218 85450 381454
rect 85686 381218 116170 381454
rect 116406 381218 146890 381454
rect 147126 381218 177610 381454
rect 177846 381218 208330 381454
rect 208566 381218 239050 381454
rect 239286 381218 269770 381454
rect 270006 381218 300490 381454
rect 300726 381218 331210 381454
rect 331446 381218 361930 381454
rect 362166 381218 392650 381454
rect 392886 381218 423370 381454
rect 423606 381218 454090 381454
rect 454326 381218 484810 381454
rect 485046 381218 515530 381454
rect 515766 381218 546250 381454
rect 546486 381218 576970 381454
rect 577206 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 24010 381134
rect 24246 380898 54730 381134
rect 54966 380898 85450 381134
rect 85686 380898 116170 381134
rect 116406 380898 146890 381134
rect 147126 380898 177610 381134
rect 177846 380898 208330 381134
rect 208566 380898 239050 381134
rect 239286 380898 269770 381134
rect 270006 380898 300490 381134
rect 300726 380898 331210 381134
rect 331446 380898 361930 381134
rect 362166 380898 392650 381134
rect 392886 380898 423370 381134
rect 423606 380898 454090 381134
rect 454326 380898 484810 381134
rect 485046 380898 515530 381134
rect 515766 380898 546250 381134
rect 546486 380898 576970 381134
rect 577206 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 8650 363454
rect 8886 363218 39370 363454
rect 39606 363218 70090 363454
rect 70326 363218 100810 363454
rect 101046 363218 131530 363454
rect 131766 363218 162250 363454
rect 162486 363218 192970 363454
rect 193206 363218 223690 363454
rect 223926 363218 254410 363454
rect 254646 363218 285130 363454
rect 285366 363218 315850 363454
rect 316086 363218 346570 363454
rect 346806 363218 377290 363454
rect 377526 363218 408010 363454
rect 408246 363218 438730 363454
rect 438966 363218 469450 363454
rect 469686 363218 500170 363454
rect 500406 363218 530890 363454
rect 531126 363218 561610 363454
rect 561846 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 8650 363134
rect 8886 362898 39370 363134
rect 39606 362898 70090 363134
rect 70326 362898 100810 363134
rect 101046 362898 131530 363134
rect 131766 362898 162250 363134
rect 162486 362898 192970 363134
rect 193206 362898 223690 363134
rect 223926 362898 254410 363134
rect 254646 362898 285130 363134
rect 285366 362898 315850 363134
rect 316086 362898 346570 363134
rect 346806 362898 377290 363134
rect 377526 362898 408010 363134
rect 408246 362898 438730 363134
rect 438966 362898 469450 363134
rect 469686 362898 500170 363134
rect 500406 362898 530890 363134
rect 531126 362898 561610 363134
rect 561846 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 24010 345454
rect 24246 345218 54730 345454
rect 54966 345218 85450 345454
rect 85686 345218 116170 345454
rect 116406 345218 146890 345454
rect 147126 345218 177610 345454
rect 177846 345218 208330 345454
rect 208566 345218 239050 345454
rect 239286 345218 269770 345454
rect 270006 345218 300490 345454
rect 300726 345218 331210 345454
rect 331446 345218 361930 345454
rect 362166 345218 392650 345454
rect 392886 345218 423370 345454
rect 423606 345218 454090 345454
rect 454326 345218 484810 345454
rect 485046 345218 515530 345454
rect 515766 345218 546250 345454
rect 546486 345218 576970 345454
rect 577206 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 24010 345134
rect 24246 344898 54730 345134
rect 54966 344898 85450 345134
rect 85686 344898 116170 345134
rect 116406 344898 146890 345134
rect 147126 344898 177610 345134
rect 177846 344898 208330 345134
rect 208566 344898 239050 345134
rect 239286 344898 269770 345134
rect 270006 344898 300490 345134
rect 300726 344898 331210 345134
rect 331446 344898 361930 345134
rect 362166 344898 392650 345134
rect 392886 344898 423370 345134
rect 423606 344898 454090 345134
rect 454326 344898 484810 345134
rect 485046 344898 515530 345134
rect 515766 344898 546250 345134
rect 546486 344898 576970 345134
rect 577206 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 8650 327454
rect 8886 327218 39370 327454
rect 39606 327218 70090 327454
rect 70326 327218 100810 327454
rect 101046 327218 131530 327454
rect 131766 327218 162250 327454
rect 162486 327218 192970 327454
rect 193206 327218 223690 327454
rect 223926 327218 254410 327454
rect 254646 327218 285130 327454
rect 285366 327218 315850 327454
rect 316086 327218 346570 327454
rect 346806 327218 377290 327454
rect 377526 327218 408010 327454
rect 408246 327218 438730 327454
rect 438966 327218 469450 327454
rect 469686 327218 500170 327454
rect 500406 327218 530890 327454
rect 531126 327218 561610 327454
rect 561846 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 8650 327134
rect 8886 326898 39370 327134
rect 39606 326898 70090 327134
rect 70326 326898 100810 327134
rect 101046 326898 131530 327134
rect 131766 326898 162250 327134
rect 162486 326898 192970 327134
rect 193206 326898 223690 327134
rect 223926 326898 254410 327134
rect 254646 326898 285130 327134
rect 285366 326898 315850 327134
rect 316086 326898 346570 327134
rect 346806 326898 377290 327134
rect 377526 326898 408010 327134
rect 408246 326898 438730 327134
rect 438966 326898 469450 327134
rect 469686 326898 500170 327134
rect 500406 326898 530890 327134
rect 531126 326898 561610 327134
rect 561846 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 24010 309454
rect 24246 309218 54730 309454
rect 54966 309218 85450 309454
rect 85686 309218 116170 309454
rect 116406 309218 146890 309454
rect 147126 309218 177610 309454
rect 177846 309218 208330 309454
rect 208566 309218 239050 309454
rect 239286 309218 269770 309454
rect 270006 309218 300490 309454
rect 300726 309218 331210 309454
rect 331446 309218 361930 309454
rect 362166 309218 392650 309454
rect 392886 309218 423370 309454
rect 423606 309218 454090 309454
rect 454326 309218 484810 309454
rect 485046 309218 515530 309454
rect 515766 309218 546250 309454
rect 546486 309218 576970 309454
rect 577206 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 24010 309134
rect 24246 308898 54730 309134
rect 54966 308898 85450 309134
rect 85686 308898 116170 309134
rect 116406 308898 146890 309134
rect 147126 308898 177610 309134
rect 177846 308898 208330 309134
rect 208566 308898 239050 309134
rect 239286 308898 269770 309134
rect 270006 308898 300490 309134
rect 300726 308898 331210 309134
rect 331446 308898 361930 309134
rect 362166 308898 392650 309134
rect 392886 308898 423370 309134
rect 423606 308898 454090 309134
rect 454326 308898 484810 309134
rect 485046 308898 515530 309134
rect 515766 308898 546250 309134
rect 546486 308898 576970 309134
rect 577206 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 8650 291454
rect 8886 291218 39370 291454
rect 39606 291218 70090 291454
rect 70326 291218 100810 291454
rect 101046 291218 131530 291454
rect 131766 291218 162250 291454
rect 162486 291218 192970 291454
rect 193206 291218 223690 291454
rect 223926 291218 254410 291454
rect 254646 291218 285130 291454
rect 285366 291218 315850 291454
rect 316086 291218 346570 291454
rect 346806 291218 377290 291454
rect 377526 291218 408010 291454
rect 408246 291218 438730 291454
rect 438966 291218 469450 291454
rect 469686 291218 500170 291454
rect 500406 291218 530890 291454
rect 531126 291218 561610 291454
rect 561846 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 8650 291134
rect 8886 290898 39370 291134
rect 39606 290898 70090 291134
rect 70326 290898 100810 291134
rect 101046 290898 131530 291134
rect 131766 290898 162250 291134
rect 162486 290898 192970 291134
rect 193206 290898 223690 291134
rect 223926 290898 254410 291134
rect 254646 290898 285130 291134
rect 285366 290898 315850 291134
rect 316086 290898 346570 291134
rect 346806 290898 377290 291134
rect 377526 290898 408010 291134
rect 408246 290898 438730 291134
rect 438966 290898 469450 291134
rect 469686 290898 500170 291134
rect 500406 290898 530890 291134
rect 531126 290898 561610 291134
rect 561846 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 24010 273454
rect 24246 273218 54730 273454
rect 54966 273218 85450 273454
rect 85686 273218 116170 273454
rect 116406 273218 146890 273454
rect 147126 273218 177610 273454
rect 177846 273218 208330 273454
rect 208566 273218 239050 273454
rect 239286 273218 269770 273454
rect 270006 273218 300490 273454
rect 300726 273218 331210 273454
rect 331446 273218 361930 273454
rect 362166 273218 392650 273454
rect 392886 273218 423370 273454
rect 423606 273218 454090 273454
rect 454326 273218 484810 273454
rect 485046 273218 515530 273454
rect 515766 273218 546250 273454
rect 546486 273218 576970 273454
rect 577206 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 24010 273134
rect 24246 272898 54730 273134
rect 54966 272898 85450 273134
rect 85686 272898 116170 273134
rect 116406 272898 146890 273134
rect 147126 272898 177610 273134
rect 177846 272898 208330 273134
rect 208566 272898 239050 273134
rect 239286 272898 269770 273134
rect 270006 272898 300490 273134
rect 300726 272898 331210 273134
rect 331446 272898 361930 273134
rect 362166 272898 392650 273134
rect 392886 272898 423370 273134
rect 423606 272898 454090 273134
rect 454326 272898 484810 273134
rect 485046 272898 515530 273134
rect 515766 272898 546250 273134
rect 546486 272898 576970 273134
rect 577206 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 8650 255454
rect 8886 255218 39370 255454
rect 39606 255218 70090 255454
rect 70326 255218 100810 255454
rect 101046 255218 131530 255454
rect 131766 255218 162250 255454
rect 162486 255218 192970 255454
rect 193206 255218 223690 255454
rect 223926 255218 254410 255454
rect 254646 255218 285130 255454
rect 285366 255218 315850 255454
rect 316086 255218 346570 255454
rect 346806 255218 377290 255454
rect 377526 255218 408010 255454
rect 408246 255218 438730 255454
rect 438966 255218 469450 255454
rect 469686 255218 500170 255454
rect 500406 255218 530890 255454
rect 531126 255218 561610 255454
rect 561846 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 8650 255134
rect 8886 254898 39370 255134
rect 39606 254898 70090 255134
rect 70326 254898 100810 255134
rect 101046 254898 131530 255134
rect 131766 254898 162250 255134
rect 162486 254898 192970 255134
rect 193206 254898 223690 255134
rect 223926 254898 254410 255134
rect 254646 254898 285130 255134
rect 285366 254898 315850 255134
rect 316086 254898 346570 255134
rect 346806 254898 377290 255134
rect 377526 254898 408010 255134
rect 408246 254898 438730 255134
rect 438966 254898 469450 255134
rect 469686 254898 500170 255134
rect 500406 254898 530890 255134
rect 531126 254898 561610 255134
rect 561846 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 24010 237454
rect 24246 237218 54730 237454
rect 54966 237218 85450 237454
rect 85686 237218 116170 237454
rect 116406 237218 146890 237454
rect 147126 237218 177610 237454
rect 177846 237218 208330 237454
rect 208566 237218 239050 237454
rect 239286 237218 269770 237454
rect 270006 237218 300490 237454
rect 300726 237218 331210 237454
rect 331446 237218 361930 237454
rect 362166 237218 392650 237454
rect 392886 237218 423370 237454
rect 423606 237218 454090 237454
rect 454326 237218 484810 237454
rect 485046 237218 515530 237454
rect 515766 237218 546250 237454
rect 546486 237218 576970 237454
rect 577206 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 24010 237134
rect 24246 236898 54730 237134
rect 54966 236898 85450 237134
rect 85686 236898 116170 237134
rect 116406 236898 146890 237134
rect 147126 236898 177610 237134
rect 177846 236898 208330 237134
rect 208566 236898 239050 237134
rect 239286 236898 269770 237134
rect 270006 236898 300490 237134
rect 300726 236898 331210 237134
rect 331446 236898 361930 237134
rect 362166 236898 392650 237134
rect 392886 236898 423370 237134
rect 423606 236898 454090 237134
rect 454326 236898 484810 237134
rect 485046 236898 515530 237134
rect 515766 236898 546250 237134
rect 546486 236898 576970 237134
rect 577206 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 8650 219454
rect 8886 219218 39370 219454
rect 39606 219218 70090 219454
rect 70326 219218 100810 219454
rect 101046 219218 131530 219454
rect 131766 219218 162250 219454
rect 162486 219218 192970 219454
rect 193206 219218 223690 219454
rect 223926 219218 254410 219454
rect 254646 219218 285130 219454
rect 285366 219218 315850 219454
rect 316086 219218 346570 219454
rect 346806 219218 377290 219454
rect 377526 219218 408010 219454
rect 408246 219218 438730 219454
rect 438966 219218 469450 219454
rect 469686 219218 500170 219454
rect 500406 219218 530890 219454
rect 531126 219218 561610 219454
rect 561846 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 8650 219134
rect 8886 218898 39370 219134
rect 39606 218898 70090 219134
rect 70326 218898 100810 219134
rect 101046 218898 131530 219134
rect 131766 218898 162250 219134
rect 162486 218898 192970 219134
rect 193206 218898 223690 219134
rect 223926 218898 254410 219134
rect 254646 218898 285130 219134
rect 285366 218898 315850 219134
rect 316086 218898 346570 219134
rect 346806 218898 377290 219134
rect 377526 218898 408010 219134
rect 408246 218898 438730 219134
rect 438966 218898 469450 219134
rect 469686 218898 500170 219134
rect 500406 218898 530890 219134
rect 531126 218898 561610 219134
rect 561846 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 24010 201454
rect 24246 201218 54730 201454
rect 54966 201218 85450 201454
rect 85686 201218 116170 201454
rect 116406 201218 146890 201454
rect 147126 201218 177610 201454
rect 177846 201218 208330 201454
rect 208566 201218 239050 201454
rect 239286 201218 269770 201454
rect 270006 201218 300490 201454
rect 300726 201218 331210 201454
rect 331446 201218 361930 201454
rect 362166 201218 392650 201454
rect 392886 201218 423370 201454
rect 423606 201218 454090 201454
rect 454326 201218 484810 201454
rect 485046 201218 515530 201454
rect 515766 201218 546250 201454
rect 546486 201218 576970 201454
rect 577206 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 24010 201134
rect 24246 200898 54730 201134
rect 54966 200898 85450 201134
rect 85686 200898 116170 201134
rect 116406 200898 146890 201134
rect 147126 200898 177610 201134
rect 177846 200898 208330 201134
rect 208566 200898 239050 201134
rect 239286 200898 269770 201134
rect 270006 200898 300490 201134
rect 300726 200898 331210 201134
rect 331446 200898 361930 201134
rect 362166 200898 392650 201134
rect 392886 200898 423370 201134
rect 423606 200898 454090 201134
rect 454326 200898 484810 201134
rect 485046 200898 515530 201134
rect 515766 200898 546250 201134
rect 546486 200898 576970 201134
rect 577206 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 8650 183454
rect 8886 183218 39370 183454
rect 39606 183218 70090 183454
rect 70326 183218 100810 183454
rect 101046 183218 131530 183454
rect 131766 183218 162250 183454
rect 162486 183218 192970 183454
rect 193206 183218 223690 183454
rect 223926 183218 254410 183454
rect 254646 183218 285130 183454
rect 285366 183218 315850 183454
rect 316086 183218 346570 183454
rect 346806 183218 377290 183454
rect 377526 183218 408010 183454
rect 408246 183218 438730 183454
rect 438966 183218 469450 183454
rect 469686 183218 500170 183454
rect 500406 183218 530890 183454
rect 531126 183218 561610 183454
rect 561846 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 8650 183134
rect 8886 182898 39370 183134
rect 39606 182898 70090 183134
rect 70326 182898 100810 183134
rect 101046 182898 131530 183134
rect 131766 182898 162250 183134
rect 162486 182898 192970 183134
rect 193206 182898 223690 183134
rect 223926 182898 254410 183134
rect 254646 182898 285130 183134
rect 285366 182898 315850 183134
rect 316086 182898 346570 183134
rect 346806 182898 377290 183134
rect 377526 182898 408010 183134
rect 408246 182898 438730 183134
rect 438966 182898 469450 183134
rect 469686 182898 500170 183134
rect 500406 182898 530890 183134
rect 531126 182898 561610 183134
rect 561846 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 24010 165454
rect 24246 165218 54730 165454
rect 54966 165218 85450 165454
rect 85686 165218 116170 165454
rect 116406 165218 146890 165454
rect 147126 165218 177610 165454
rect 177846 165218 208330 165454
rect 208566 165218 239050 165454
rect 239286 165218 269770 165454
rect 270006 165218 300490 165454
rect 300726 165218 331210 165454
rect 331446 165218 361930 165454
rect 362166 165218 392650 165454
rect 392886 165218 423370 165454
rect 423606 165218 454090 165454
rect 454326 165218 484810 165454
rect 485046 165218 515530 165454
rect 515766 165218 546250 165454
rect 546486 165218 576970 165454
rect 577206 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 24010 165134
rect 24246 164898 54730 165134
rect 54966 164898 85450 165134
rect 85686 164898 116170 165134
rect 116406 164898 146890 165134
rect 147126 164898 177610 165134
rect 177846 164898 208330 165134
rect 208566 164898 239050 165134
rect 239286 164898 269770 165134
rect 270006 164898 300490 165134
rect 300726 164898 331210 165134
rect 331446 164898 361930 165134
rect 362166 164898 392650 165134
rect 392886 164898 423370 165134
rect 423606 164898 454090 165134
rect 454326 164898 484810 165134
rect 485046 164898 515530 165134
rect 515766 164898 546250 165134
rect 546486 164898 576970 165134
rect 577206 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 8650 147454
rect 8886 147218 39370 147454
rect 39606 147218 70090 147454
rect 70326 147218 100810 147454
rect 101046 147218 131530 147454
rect 131766 147218 162250 147454
rect 162486 147218 192970 147454
rect 193206 147218 223690 147454
rect 223926 147218 254410 147454
rect 254646 147218 285130 147454
rect 285366 147218 315850 147454
rect 316086 147218 346570 147454
rect 346806 147218 377290 147454
rect 377526 147218 408010 147454
rect 408246 147218 438730 147454
rect 438966 147218 469450 147454
rect 469686 147218 500170 147454
rect 500406 147218 530890 147454
rect 531126 147218 561610 147454
rect 561846 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 8650 147134
rect 8886 146898 39370 147134
rect 39606 146898 70090 147134
rect 70326 146898 100810 147134
rect 101046 146898 131530 147134
rect 131766 146898 162250 147134
rect 162486 146898 192970 147134
rect 193206 146898 223690 147134
rect 223926 146898 254410 147134
rect 254646 146898 285130 147134
rect 285366 146898 315850 147134
rect 316086 146898 346570 147134
rect 346806 146898 377290 147134
rect 377526 146898 408010 147134
rect 408246 146898 438730 147134
rect 438966 146898 469450 147134
rect 469686 146898 500170 147134
rect 500406 146898 530890 147134
rect 531126 146898 561610 147134
rect 561846 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 24010 129454
rect 24246 129218 54730 129454
rect 54966 129218 85450 129454
rect 85686 129218 116170 129454
rect 116406 129218 146890 129454
rect 147126 129218 177610 129454
rect 177846 129218 208330 129454
rect 208566 129218 239050 129454
rect 239286 129218 269770 129454
rect 270006 129218 300490 129454
rect 300726 129218 331210 129454
rect 331446 129218 361930 129454
rect 362166 129218 392650 129454
rect 392886 129218 423370 129454
rect 423606 129218 454090 129454
rect 454326 129218 484810 129454
rect 485046 129218 515530 129454
rect 515766 129218 546250 129454
rect 546486 129218 576970 129454
rect 577206 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 24010 129134
rect 24246 128898 54730 129134
rect 54966 128898 85450 129134
rect 85686 128898 116170 129134
rect 116406 128898 146890 129134
rect 147126 128898 177610 129134
rect 177846 128898 208330 129134
rect 208566 128898 239050 129134
rect 239286 128898 269770 129134
rect 270006 128898 300490 129134
rect 300726 128898 331210 129134
rect 331446 128898 361930 129134
rect 362166 128898 392650 129134
rect 392886 128898 423370 129134
rect 423606 128898 454090 129134
rect 454326 128898 484810 129134
rect 485046 128898 515530 129134
rect 515766 128898 546250 129134
rect 546486 128898 576970 129134
rect 577206 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 8650 111454
rect 8886 111218 39370 111454
rect 39606 111218 70090 111454
rect 70326 111218 100810 111454
rect 101046 111218 131530 111454
rect 131766 111218 162250 111454
rect 162486 111218 192970 111454
rect 193206 111218 223690 111454
rect 223926 111218 254410 111454
rect 254646 111218 285130 111454
rect 285366 111218 315850 111454
rect 316086 111218 346570 111454
rect 346806 111218 377290 111454
rect 377526 111218 408010 111454
rect 408246 111218 438730 111454
rect 438966 111218 469450 111454
rect 469686 111218 500170 111454
rect 500406 111218 530890 111454
rect 531126 111218 561610 111454
rect 561846 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 8650 111134
rect 8886 110898 39370 111134
rect 39606 110898 70090 111134
rect 70326 110898 100810 111134
rect 101046 110898 131530 111134
rect 131766 110898 162250 111134
rect 162486 110898 192970 111134
rect 193206 110898 223690 111134
rect 223926 110898 254410 111134
rect 254646 110898 285130 111134
rect 285366 110898 315850 111134
rect 316086 110898 346570 111134
rect 346806 110898 377290 111134
rect 377526 110898 408010 111134
rect 408246 110898 438730 111134
rect 438966 110898 469450 111134
rect 469686 110898 500170 111134
rect 500406 110898 530890 111134
rect 531126 110898 561610 111134
rect 561846 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 24010 93454
rect 24246 93218 54730 93454
rect 54966 93218 85450 93454
rect 85686 93218 116170 93454
rect 116406 93218 146890 93454
rect 147126 93218 177610 93454
rect 177846 93218 208330 93454
rect 208566 93218 239050 93454
rect 239286 93218 269770 93454
rect 270006 93218 300490 93454
rect 300726 93218 331210 93454
rect 331446 93218 361930 93454
rect 362166 93218 392650 93454
rect 392886 93218 423370 93454
rect 423606 93218 454090 93454
rect 454326 93218 484810 93454
rect 485046 93218 515530 93454
rect 515766 93218 546250 93454
rect 546486 93218 576970 93454
rect 577206 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 24010 93134
rect 24246 92898 54730 93134
rect 54966 92898 85450 93134
rect 85686 92898 116170 93134
rect 116406 92898 146890 93134
rect 147126 92898 177610 93134
rect 177846 92898 208330 93134
rect 208566 92898 239050 93134
rect 239286 92898 269770 93134
rect 270006 92898 300490 93134
rect 300726 92898 331210 93134
rect 331446 92898 361930 93134
rect 362166 92898 392650 93134
rect 392886 92898 423370 93134
rect 423606 92898 454090 93134
rect 454326 92898 484810 93134
rect 485046 92898 515530 93134
rect 515766 92898 546250 93134
rect 546486 92898 576970 93134
rect 577206 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 8650 75454
rect 8886 75218 39370 75454
rect 39606 75218 70090 75454
rect 70326 75218 100810 75454
rect 101046 75218 131530 75454
rect 131766 75218 162250 75454
rect 162486 75218 192970 75454
rect 193206 75218 223690 75454
rect 223926 75218 254410 75454
rect 254646 75218 285130 75454
rect 285366 75218 315850 75454
rect 316086 75218 346570 75454
rect 346806 75218 377290 75454
rect 377526 75218 408010 75454
rect 408246 75218 438730 75454
rect 438966 75218 469450 75454
rect 469686 75218 500170 75454
rect 500406 75218 530890 75454
rect 531126 75218 561610 75454
rect 561846 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 8650 75134
rect 8886 74898 39370 75134
rect 39606 74898 70090 75134
rect 70326 74898 100810 75134
rect 101046 74898 131530 75134
rect 131766 74898 162250 75134
rect 162486 74898 192970 75134
rect 193206 74898 223690 75134
rect 223926 74898 254410 75134
rect 254646 74898 285130 75134
rect 285366 74898 315850 75134
rect 316086 74898 346570 75134
rect 346806 74898 377290 75134
rect 377526 74898 408010 75134
rect 408246 74898 438730 75134
rect 438966 74898 469450 75134
rect 469686 74898 500170 75134
rect 500406 74898 530890 75134
rect 531126 74898 561610 75134
rect 561846 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 24010 57454
rect 24246 57218 54730 57454
rect 54966 57218 85450 57454
rect 85686 57218 116170 57454
rect 116406 57218 146890 57454
rect 147126 57218 177610 57454
rect 177846 57218 208330 57454
rect 208566 57218 239050 57454
rect 239286 57218 269770 57454
rect 270006 57218 300490 57454
rect 300726 57218 331210 57454
rect 331446 57218 361930 57454
rect 362166 57218 392650 57454
rect 392886 57218 423370 57454
rect 423606 57218 454090 57454
rect 454326 57218 484810 57454
rect 485046 57218 515530 57454
rect 515766 57218 546250 57454
rect 546486 57218 576970 57454
rect 577206 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 24010 57134
rect 24246 56898 54730 57134
rect 54966 56898 85450 57134
rect 85686 56898 116170 57134
rect 116406 56898 146890 57134
rect 147126 56898 177610 57134
rect 177846 56898 208330 57134
rect 208566 56898 239050 57134
rect 239286 56898 269770 57134
rect 270006 56898 300490 57134
rect 300726 56898 331210 57134
rect 331446 56898 361930 57134
rect 362166 56898 392650 57134
rect 392886 56898 423370 57134
rect 423606 56898 454090 57134
rect 454326 56898 484810 57134
rect 485046 56898 515530 57134
rect 515766 56898 546250 57134
rect 546486 56898 576970 57134
rect 577206 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 8650 39454
rect 8886 39218 39370 39454
rect 39606 39218 70090 39454
rect 70326 39218 100810 39454
rect 101046 39218 131530 39454
rect 131766 39218 162250 39454
rect 162486 39218 192970 39454
rect 193206 39218 223690 39454
rect 223926 39218 254410 39454
rect 254646 39218 285130 39454
rect 285366 39218 315850 39454
rect 316086 39218 346570 39454
rect 346806 39218 377290 39454
rect 377526 39218 408010 39454
rect 408246 39218 438730 39454
rect 438966 39218 469450 39454
rect 469686 39218 500170 39454
rect 500406 39218 530890 39454
rect 531126 39218 561610 39454
rect 561846 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 8650 39134
rect 8886 38898 39370 39134
rect 39606 38898 70090 39134
rect 70326 38898 100810 39134
rect 101046 38898 131530 39134
rect 131766 38898 162250 39134
rect 162486 38898 192970 39134
rect 193206 38898 223690 39134
rect 223926 38898 254410 39134
rect 254646 38898 285130 39134
rect 285366 38898 315850 39134
rect 316086 38898 346570 39134
rect 346806 38898 377290 39134
rect 377526 38898 408010 39134
rect 408246 38898 438730 39134
rect 438966 38898 469450 39134
rect 469686 38898 500170 39134
rect 500406 38898 530890 39134
rect 531126 38898 561610 39134
rect 561846 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 24010 21454
rect 24246 21218 54730 21454
rect 54966 21218 85450 21454
rect 85686 21218 116170 21454
rect 116406 21218 146890 21454
rect 147126 21218 177610 21454
rect 177846 21218 208330 21454
rect 208566 21218 239050 21454
rect 239286 21218 269770 21454
rect 270006 21218 300490 21454
rect 300726 21218 331210 21454
rect 331446 21218 361930 21454
rect 362166 21218 392650 21454
rect 392886 21218 423370 21454
rect 423606 21218 454090 21454
rect 454326 21218 484810 21454
rect 485046 21218 515530 21454
rect 515766 21218 546250 21454
rect 546486 21218 576970 21454
rect 577206 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 24010 21134
rect 24246 20898 54730 21134
rect 54966 20898 85450 21134
rect 85686 20898 116170 21134
rect 116406 20898 146890 21134
rect 147126 20898 177610 21134
rect 177846 20898 208330 21134
rect 208566 20898 239050 21134
rect 239286 20898 269770 21134
rect 270006 20898 300490 21134
rect 300726 20898 331210 21134
rect 331446 20898 361930 21134
rect 362166 20898 392650 21134
rect 392886 20898 423370 21134
rect 423606 20898 454090 21134
rect 454326 20898 484810 21134
rect 485046 20898 515530 21134
rect 515766 20898 546250 21134
rect 546486 20898 576970 21134
rect 577206 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1635585791
transform 1 0 4400 0 1 4400
box 566 0 574618 695200
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 2400 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 701600 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 701600 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 701600 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 701600 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 701600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 701600 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 701600 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 701600 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 701600 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 701600 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 701600 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 701600 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 701600 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 701600 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 701600 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 701600 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 701600 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 2400 8 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 701600 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 701600 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 701600 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 701600 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 701600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 701600 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 701600 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 701600 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 701600 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 701600 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 701600 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 701600 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 701600 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 701600 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 701600 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 701600 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 701600 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 2400 8 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 701600 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 701600 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 701600 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 701600 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 701600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 701600 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 701600 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 701600 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 701600 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 701600 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 701600 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 701600 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 701600 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 701600 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 701600 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 701600 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 2400 8 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 701600 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 701600 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 701600 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 701600 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 701600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 701600 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 701600 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 701600 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 701600 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 701600 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 701600 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 701600 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 701600 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 701600 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 701600 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 701600 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 2400 8 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 701600 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 701600 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 701600 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 701600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 701600 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 701600 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 701600 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 701600 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 701600 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 701600 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 701600 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 701600 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 701600 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 701600 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 701600 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 701600 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 2400 8 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 701600 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 701600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 701600 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 701600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 701600 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 701600 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 701600 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 701600 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 701600 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 701600 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 701600 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 701600 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 701600 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 701600 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 701600 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 701600 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 2400 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 701600 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 701600 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 701600 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 701600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 701600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 701600 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 701600 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 701600 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 701600 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 701600 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 701600 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 701600 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 701600 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 701600 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 701600 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 701600 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 2400 8 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 701600 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 701600 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 701600 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 701600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 701600 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 701600 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 701600 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 701600 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 701600 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 701600 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 701600 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 701600 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 701600 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 701600 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 701600 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 701600 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
