magic
tech sky130A
magscale 1 2
timestamp 1636617456
<< locali >>
rect 435097 564519 435131 564689
rect 456073 136391 456107 136561
rect 195253 136051 195287 136289
rect 185593 135779 185627 136017
rect 190377 135779 190411 135949
rect 267197 135915 267231 136221
rect 422987 136017 423137 136051
rect 200681 135643 200715 135745
rect 220001 135711 220035 135881
rect 199945 135507 199979 135609
rect 222301 135507 222335 135881
rect 427093 135847 427127 136357
rect 461225 136323 461259 136425
rect 475393 136187 475427 136289
rect 480361 135371 480395 135745
rect 480453 135439 480487 135813
rect 496829 135439 496863 136561
rect 427001 4743 427035 5049
rect 514033 4743 514067 4913
rect 85497 3451 85531 4165
rect 90281 3519 90315 4165
rect 95525 3791 95559 3893
rect 95617 3723 95651 3893
rect 95375 3689 95651 3723
rect 106841 3383 106875 4165
rect 384681 4165 384899 4199
rect 384681 4131 384715 4165
rect 108313 3383 108347 3961
rect 53849 3111 53883 3281
rect 123401 3247 123435 4029
rect 146953 3587 146987 3893
rect 134073 3247 134107 3417
rect 146861 3247 146895 3553
rect 147045 3519 147079 3893
rect 193321 3587 193355 3825
rect 214573 3587 214607 3757
rect 384681 3655 384715 3825
rect 384773 3791 384807 4097
rect 384865 3995 384899 4165
rect 387533 3655 387567 3825
rect 324605 3519 324639 3621
rect 390385 3587 390419 3825
rect 394709 3689 394893 3723
rect 394709 3655 394743 3689
rect 352941 3247 352975 3349
rect 355885 3281 356161 3315
rect 355885 3111 355919 3281
rect 355977 3111 356011 3213
rect 213745 2975 213779 3077
rect 542829 3043 542863 3213
<< viali >>
rect 435097 564689 435131 564723
rect 435097 564485 435131 564519
rect 456073 136561 456107 136595
rect 496829 136561 496863 136595
rect 427093 136357 427127 136391
rect 456073 136357 456107 136391
rect 461225 136425 461259 136459
rect 195253 136289 195287 136323
rect 185593 136017 185627 136051
rect 195253 136017 195287 136051
rect 267197 136221 267231 136255
rect 185593 135745 185627 135779
rect 190377 135949 190411 135983
rect 422953 136017 422987 136051
rect 423137 136017 423171 136051
rect 220001 135881 220035 135915
rect 190377 135745 190411 135779
rect 200681 135745 200715 135779
rect 220001 135677 220035 135711
rect 222301 135881 222335 135915
rect 267197 135881 267231 135915
rect 199945 135609 199979 135643
rect 200681 135609 200715 135643
rect 199945 135473 199979 135507
rect 461225 136289 461259 136323
rect 475393 136289 475427 136323
rect 475393 136153 475427 136187
rect 427093 135813 427127 135847
rect 480453 135813 480487 135847
rect 222301 135473 222335 135507
rect 480361 135745 480395 135779
rect 480453 135405 480487 135439
rect 496829 135405 496863 135439
rect 480361 135337 480395 135371
rect 427001 5049 427035 5083
rect 427001 4709 427035 4743
rect 514033 4913 514067 4947
rect 514033 4709 514067 4743
rect 85497 4165 85531 4199
rect 90281 4165 90315 4199
rect 106841 4165 106875 4199
rect 95525 3893 95559 3927
rect 95525 3757 95559 3791
rect 95617 3893 95651 3927
rect 95341 3689 95375 3723
rect 90281 3485 90315 3519
rect 85497 3417 85531 3451
rect 384681 4097 384715 4131
rect 384773 4097 384807 4131
rect 123401 4029 123435 4063
rect 106841 3349 106875 3383
rect 108313 3961 108347 3995
rect 108313 3349 108347 3383
rect 53849 3281 53883 3315
rect 146953 3893 146987 3927
rect 146861 3553 146895 3587
rect 146953 3553 146987 3587
rect 147045 3893 147079 3927
rect 123401 3213 123435 3247
rect 134073 3417 134107 3451
rect 134073 3213 134107 3247
rect 193321 3825 193355 3859
rect 384681 3825 384715 3859
rect 193321 3553 193355 3587
rect 214573 3757 214607 3791
rect 384865 3961 384899 3995
rect 384773 3757 384807 3791
rect 387533 3825 387567 3859
rect 214573 3553 214607 3587
rect 324605 3621 324639 3655
rect 384681 3621 384715 3655
rect 387533 3621 387567 3655
rect 390385 3825 390419 3859
rect 147045 3485 147079 3519
rect 394893 3689 394927 3723
rect 394709 3621 394743 3655
rect 390385 3553 390419 3587
rect 324605 3485 324639 3519
rect 146861 3213 146895 3247
rect 352941 3349 352975 3383
rect 352941 3213 352975 3247
rect 356161 3281 356195 3315
rect 53849 3077 53883 3111
rect 213745 3077 213779 3111
rect 355885 3077 355919 3111
rect 355977 3213 356011 3247
rect 355977 3077 356011 3111
rect 542829 3213 542863 3247
rect 542829 3009 542863 3043
rect 213745 2941 213779 2975
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 322934 700992 322940 701004
rect 154172 700964 322940 700992
rect 154172 700952 154178 700964
rect 322934 700952 322940 700964
rect 322992 700952 322998 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 318794 700924 318800 700936
rect 137888 700896 318800 700924
rect 137888 700884 137894 700896
rect 318794 700884 318800 700896
rect 318852 700884 318858 700936
rect 264882 700816 264888 700868
rect 264940 700856 264946 700868
rect 462314 700856 462320 700868
rect 264940 700828 462320 700856
rect 264940 700816 264946 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 269022 700748 269028 700800
rect 269080 700788 269086 700800
rect 478506 700788 478512 700800
rect 269080 700760 478512 700788
rect 269080 700748 269086 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 333974 700720 333980 700732
rect 89220 700692 333980 700720
rect 89220 700680 89226 700692
rect 333974 700680 333980 700692
rect 334032 700680 334038 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 329834 700652 329840 700664
rect 73028 700624 329840 700652
rect 73028 700612 73034 700624
rect 329834 700612 329840 700624
rect 329892 700612 329898 700664
rect 253842 700544 253848 700596
rect 253900 700584 253906 700596
rect 527174 700584 527180 700596
rect 253900 700556 527180 700584
rect 253900 700544 253906 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 256602 700476 256608 700528
rect 256660 700516 256666 700528
rect 543458 700516 543464 700528
rect 256660 700488 543464 700516
rect 256660 700476 256666 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 338114 700448 338120 700460
rect 40552 700420 338120 700448
rect 40552 700408 40558 700420
rect 338114 700408 338120 700420
rect 338172 700408 338178 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 345014 700380 345020 700392
rect 24360 700352 345020 700380
rect 24360 700340 24366 700352
rect 345014 700340 345020 700352
rect 345072 700340 345078 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 342254 700312 342260 700324
rect 8168 700284 342260 700312
rect 8168 700272 8174 700284
rect 342254 700272 342260 700284
rect 342312 700272 342318 700324
rect 280062 700204 280068 700256
rect 280120 700244 280126 700256
rect 413646 700244 413652 700256
rect 280120 700216 413652 700244
rect 280120 700204 280126 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 275922 700136 275928 700188
rect 275980 700176 275986 700188
rect 397454 700176 397460 700188
rect 275980 700148 397460 700176
rect 275980 700136 275986 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 307754 700108 307760 700120
rect 202840 700080 307760 700108
rect 202840 700068 202846 700080
rect 307754 700068 307760 700080
rect 307812 700068 307818 700120
rect 218974 700000 218980 700052
rect 219032 700040 219038 700052
rect 311894 700040 311900 700052
rect 219032 700012 311900 700040
rect 219032 700000 219038 700012
rect 311894 700000 311900 700012
rect 311952 700000 311958 700052
rect 291102 699932 291108 699984
rect 291160 699972 291166 699984
rect 348786 699972 348792 699984
rect 291160 699944 348792 699972
rect 291160 699932 291166 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 286962 699864 286968 699916
rect 287020 699904 287026 699916
rect 332502 699904 332508 699916
rect 287020 699876 332508 699904
rect 287020 699864 287026 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 296714 699836 296720 699848
rect 267700 699808 296720 699836
rect 267700 699796 267706 699808
rect 296714 699796 296720 699808
rect 296772 699796 296778 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 300854 699768 300860 699780
rect 283892 699740 300860 699768
rect 283892 699728 283898 699740
rect 300854 699728 300860 699740
rect 300912 699728 300918 699780
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 242802 696940 242808 696992
rect 242860 696980 242866 696992
rect 580166 696980 580172 696992
rect 242860 696952 580172 696980
rect 242860 696940 242866 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 245562 683204 245568 683256
rect 245620 683244 245626 683256
rect 580166 683244 580172 683256
rect 245620 683216 580172 683244
rect 245620 683204 245626 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 349154 683176 349160 683188
rect 3476 683148 349160 683176
rect 3476 683136 3482 683148
rect 349154 683136 349160 683148
rect 349212 683136 349218 683188
rect 238662 670760 238668 670812
rect 238720 670800 238726 670812
rect 580166 670800 580172 670812
rect 238720 670772 580172 670800
rect 238720 670760 238726 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 356054 670732 356060 670744
rect 3568 670704 356060 670732
rect 3568 670692 3574 670704
rect 356054 670692 356060 670704
rect 356112 670692 356118 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 353294 656928 353300 656940
rect 3476 656900 353300 656928
rect 3476 656888 3482 656900
rect 353294 656888 353300 656900
rect 353352 656888 353358 656940
rect 231762 643084 231768 643136
rect 231820 643124 231826 643136
rect 580166 643124 580172 643136
rect 231820 643096 580172 643124
rect 231820 643084 231826 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 360194 632108 360200 632120
rect 3476 632080 360200 632108
rect 3476 632068 3482 632080
rect 360194 632068 360200 632080
rect 360252 632068 360258 632120
rect 234522 630640 234528 630692
rect 234580 630680 234586 630692
rect 580166 630680 580172 630692
rect 234580 630652 580172 630680
rect 234580 630640 234586 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 367094 618304 367100 618316
rect 3200 618276 367100 618304
rect 3200 618264 3206 618276
rect 367094 618264 367100 618276
rect 367152 618264 367158 618316
rect 227622 616836 227628 616888
rect 227680 616876 227686 616888
rect 580166 616876 580172 616888
rect 227680 616848 580172 616876
rect 227680 616836 227686 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 364426 605860 364432 605872
rect 3292 605832 364432 605860
rect 3292 605820 3298 605832
rect 364426 605820 364432 605832
rect 364484 605820 364490 605872
rect 219342 590656 219348 590708
rect 219400 590696 219406 590708
rect 579798 590696 579804 590708
rect 219400 590668 579804 590696
rect 219400 590656 219406 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 371234 579680 371240 579692
rect 3384 579652 371240 579680
rect 3384 579640 3390 579652
rect 371234 579640 371240 579652
rect 371292 579640 371298 579692
rect 223482 576852 223488 576904
rect 223540 576892 223546 576904
rect 580166 576892 580172 576904
rect 223540 576864 580172 576892
rect 223540 576852 223546 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 175090 569032 175096 569084
rect 175148 569072 175154 569084
rect 556798 569072 556804 569084
rect 175148 569044 556804 569072
rect 175148 569032 175154 569044
rect 556798 569032 556804 569044
rect 556856 569032 556862 569084
rect 152734 568964 152740 569016
rect 152792 569004 152798 569016
rect 547138 569004 547144 569016
rect 152792 568976 547144 569004
rect 152792 568964 152798 568976
rect 547138 568964 547144 568976
rect 547196 568964 547202 569016
rect 130378 568896 130384 568948
rect 130436 568936 130442 568948
rect 542998 568936 543004 568948
rect 130436 568908 543004 568936
rect 130436 568896 130442 568908
rect 542998 568896 543004 568908
rect 543056 568896 543062 568948
rect 7558 568828 7564 568880
rect 7616 568868 7622 568880
rect 423950 568868 423956 568880
rect 7616 568840 423956 568868
rect 7616 568828 7622 568840
rect 423950 568828 423956 568840
rect 424008 568828 424014 568880
rect 119154 568760 119160 568812
rect 119212 568800 119218 568812
rect 540238 568800 540244 568812
rect 119212 568772 540244 568800
rect 119212 568760 119218 568772
rect 540238 568760 540244 568772
rect 540296 568760 540302 568812
rect 111702 568692 111708 568744
rect 111760 568732 111766 568744
rect 560938 568732 560944 568744
rect 111760 568704 560944 568732
rect 111760 568692 111766 568704
rect 560938 568692 560944 568704
rect 560996 568692 561002 568744
rect 100570 568624 100576 568676
rect 100628 568664 100634 568676
rect 558178 568664 558184 568676
rect 100628 568636 558184 568664
rect 100628 568624 100634 568636
rect 558178 568624 558184 568636
rect 558236 568624 558242 568676
rect 14458 568556 14464 568608
rect 14516 568596 14522 568608
rect 502426 568596 502432 568608
rect 14516 568568 502432 568596
rect 14516 568556 14522 568568
rect 502426 568556 502432 568568
rect 502484 568556 502490 568608
rect 227162 568488 227168 568540
rect 227220 568528 227226 568540
rect 227622 568528 227628 568540
rect 227220 568500 227628 568528
rect 227220 568488 227226 568500
rect 227622 568488 227628 568500
rect 227680 568488 227686 568540
rect 230934 568488 230940 568540
rect 230992 568528 230998 568540
rect 231762 568528 231768 568540
rect 230992 568500 231768 568528
rect 230992 568488 230998 568500
rect 231762 568488 231768 568500
rect 231820 568488 231826 568540
rect 242066 568488 242072 568540
rect 242124 568528 242130 568540
rect 242802 568528 242808 568540
rect 242124 568500 242808 568528
rect 242124 568488 242130 568500
rect 242802 568488 242808 568500
rect 242860 568488 242866 568540
rect 253290 568488 253296 568540
rect 253348 568528 253354 568540
rect 253842 568528 253848 568540
rect 253348 568500 253848 568528
rect 253348 568488 253354 568500
rect 253842 568488 253848 568500
rect 253900 568488 253906 568540
rect 264422 568488 264428 568540
rect 264480 568528 264486 568540
rect 264882 568528 264888 568540
rect 264480 568500 264888 568528
rect 264480 568488 264486 568500
rect 264882 568488 264888 568500
rect 264940 568488 264946 568540
rect 268194 568488 268200 568540
rect 268252 568528 268258 568540
rect 269022 568528 269028 568540
rect 268252 568500 269028 568528
rect 268252 568488 268258 568500
rect 269022 568488 269028 568500
rect 269080 568488 269086 568540
rect 279326 568488 279332 568540
rect 279384 568528 279390 568540
rect 280062 568528 280068 568540
rect 279384 568500 280068 568528
rect 279384 568488 279390 568500
rect 280062 568488 280068 568500
rect 280120 568488 280126 568540
rect 290550 568488 290556 568540
rect 290608 568528 290614 568540
rect 291102 568528 291108 568540
rect 290608 568500 291108 568528
rect 290608 568488 290614 568500
rect 291102 568488 291108 568500
rect 291160 568488 291166 568540
rect 293862 568488 293868 568540
rect 293920 568528 293926 568540
rect 299474 568528 299480 568540
rect 293920 568500 299480 568528
rect 293920 568488 293926 568500
rect 299474 568488 299480 568500
rect 299532 568488 299538 568540
rect 235902 568420 235908 568472
rect 235960 568460 235966 568472
rect 304994 568460 305000 568472
rect 235960 568432 305000 568460
rect 235960 568420 235966 568432
rect 304994 568420 305000 568432
rect 305052 568420 305058 568472
rect 282822 568352 282828 568404
rect 282880 568392 282886 568404
rect 364334 568392 364340 568404
rect 282880 568364 364340 568392
rect 282880 568352 282886 568364
rect 364334 568352 364340 568364
rect 364392 568352 364398 568404
rect 171042 568284 171048 568336
rect 171100 568324 171106 568336
rect 316034 568324 316040 568336
rect 171100 568296 316040 568324
rect 171100 568284 171106 568296
rect 316034 568284 316040 568296
rect 316092 568284 316098 568336
rect 271782 568216 271788 568268
rect 271840 568256 271846 568268
rect 429194 568256 429200 568268
rect 271840 568228 429200 568256
rect 271840 568216 271846 568228
rect 429194 568216 429200 568228
rect 429252 568216 429258 568268
rect 106182 568148 106188 568200
rect 106240 568188 106246 568200
rect 327074 568188 327080 568200
rect 106240 568160 327080 568188
rect 106240 568148 106246 568160
rect 327074 568148 327080 568160
rect 327132 568148 327138 568200
rect 260558 568080 260564 568132
rect 260616 568120 260622 568132
rect 494054 568120 494060 568132
rect 260616 568092 494060 568120
rect 260616 568080 260622 568092
rect 494054 568080 494060 568092
rect 494112 568080 494118 568132
rect 249518 568012 249524 568064
rect 249576 568052 249582 568064
rect 558914 568052 558920 568064
rect 249576 568024 558920 568052
rect 249576 568012 249582 568024
rect 558914 568012 558920 568024
rect 558972 568012 558978 568064
rect 61378 567944 61384 567996
rect 61436 567984 61442 567996
rect 386690 567984 386696 567996
rect 61436 567956 386696 567984
rect 61436 567944 61442 567956
rect 386690 567944 386696 567956
rect 386748 567944 386754 567996
rect 189902 567876 189908 567928
rect 189960 567916 189966 567928
rect 525058 567916 525064 567928
rect 189960 567888 525064 567916
rect 189960 567876 189966 567888
rect 525058 567876 525064 567888
rect 525116 567876 525122 567928
rect 178770 567808 178776 567860
rect 178828 567848 178834 567860
rect 522298 567848 522304 567860
rect 178828 567820 522304 567848
rect 178828 567808 178834 567820
rect 522298 567808 522304 567820
rect 522356 567808 522362 567860
rect 57238 567740 57244 567792
rect 57296 567780 57302 567792
rect 409046 567780 409052 567792
rect 57296 567752 409052 567780
rect 57296 567740 57302 567752
rect 409046 567740 409052 567752
rect 409104 567740 409110 567792
rect 167638 567672 167644 567724
rect 167696 567712 167702 567724
rect 520918 567712 520924 567724
rect 167696 567684 520924 567712
rect 167696 567672 167702 567684
rect 520918 567672 520924 567684
rect 520976 567672 520982 567724
rect 156414 567604 156420 567656
rect 156472 567644 156478 567656
rect 519538 567644 519544 567656
rect 156472 567616 519544 567644
rect 156472 567604 156478 567616
rect 519538 567604 519544 567616
rect 519596 567604 519602 567656
rect 145282 567536 145288 567588
rect 145340 567576 145346 567588
rect 518158 567576 518164 567588
rect 145340 567548 518164 567576
rect 145340 567536 145346 567548
rect 518158 567536 518164 567548
rect 518216 567536 518222 567588
rect 51718 567468 51724 567520
rect 51776 567508 51782 567520
rect 431402 567508 431408 567520
rect 51776 567480 431408 567508
rect 51776 567468 51782 567480
rect 431402 567468 431408 567480
rect 431460 567468 431466 567520
rect 133782 567400 133788 567452
rect 133840 567440 133846 567452
rect 515398 567440 515404 567452
rect 133840 567412 515404 567440
rect 133840 567400 133846 567412
rect 515398 567400 515404 567412
rect 515456 567400 515462 567452
rect 4890 567332 4896 567384
rect 4948 567372 4954 567384
rect 446306 567372 446312 567384
rect 4948 567344 446312 567372
rect 4948 567332 4954 567344
rect 446306 567332 446312 567344
rect 446364 567332 446370 567384
rect 17218 567264 17224 567316
rect 17276 567304 17282 567316
rect 468662 567304 468668 567316
rect 17276 567276 468668 567304
rect 17276 567264 17282 567276
rect 468662 567264 468668 567276
rect 468720 567264 468726 567316
rect 4798 567196 4804 567248
rect 4856 567236 4862 567248
rect 457438 567236 457444 567248
rect 4856 567208 457444 567236
rect 4856 567196 4862 567208
rect 457438 567196 457444 567208
rect 457496 567196 457502 567248
rect 204806 567060 204812 567112
rect 204864 567100 204870 567112
rect 507118 567100 507124 567112
rect 204864 567072 507124 567100
rect 204864 567060 204870 567072
rect 507118 567060 507124 567072
rect 507176 567060 507182 567112
rect 193674 566992 193680 567044
rect 193732 567032 193738 567044
rect 505738 567032 505744 567044
rect 193732 567004 505744 567032
rect 193732 566992 193738 567004
rect 505738 566992 505744 567004
rect 505796 566992 505802 567044
rect 79318 566924 79324 566976
rect 79376 566964 79382 566976
rect 405274 566964 405280 566976
rect 79376 566936 405280 566964
rect 79376 566924 79382 566936
rect 405274 566924 405280 566936
rect 405332 566924 405338 566976
rect 65518 566856 65524 566908
rect 65576 566896 65582 566908
rect 394142 566896 394148 566908
rect 65576 566868 394148 566896
rect 65576 566856 65582 566868
rect 394142 566856 394148 566868
rect 394200 566856 394206 566908
rect 43438 566788 43444 566840
rect 43496 566828 43502 566840
rect 383010 566828 383016 566840
rect 43496 566800 383016 566828
rect 43496 566788 43502 566800
rect 383010 566788 383016 566800
rect 383068 566788 383074 566840
rect 75178 566720 75184 566772
rect 75236 566760 75242 566772
rect 416774 566760 416780 566772
rect 75236 566732 416780 566760
rect 75236 566720 75242 566732
rect 416774 566720 416780 566732
rect 416832 566720 416838 566772
rect 53098 566652 53104 566704
rect 53156 566692 53162 566704
rect 397914 566692 397920 566704
rect 53156 566664 397920 566692
rect 53156 566652 53162 566664
rect 397914 566652 397920 566664
rect 397972 566652 397978 566704
rect 197262 566584 197268 566636
rect 197320 566624 197326 566636
rect 548518 566624 548524 566636
rect 197320 566596 548524 566624
rect 197320 566584 197326 566596
rect 548518 566584 548524 566596
rect 548576 566584 548582 566636
rect 76558 566516 76564 566568
rect 76616 566556 76622 566568
rect 438854 566556 438860 566568
rect 76616 566528 438860 566556
rect 76616 566516 76622 566528
rect 438854 566516 438860 566528
rect 438912 566516 438918 566568
rect 170950 566448 170956 566500
rect 171008 566488 171014 566500
rect 533338 566488 533344 566500
rect 171008 566460 533344 566488
rect 171008 566448 171014 566460
rect 533338 566448 533344 566460
rect 533396 566448 533402 566500
rect 54478 566380 54484 566432
rect 54536 566420 54542 566432
rect 420178 566420 420184 566432
rect 54536 566392 420184 566420
rect 54536 566380 54542 566392
rect 420178 566380 420184 566392
rect 420236 566380 420242 566432
rect 3418 566312 3424 566364
rect 3476 566352 3482 566364
rect 379514 566352 379520 566364
rect 3476 566324 379520 566352
rect 3476 566312 3482 566324
rect 379514 566312 379520 566324
rect 379572 566312 379578 566364
rect 68278 566244 68284 566296
rect 68336 566284 68342 566296
rect 461210 566284 461216 566296
rect 68336 566256 461216 566284
rect 68336 566244 68342 566256
rect 461210 566244 461216 566256
rect 461268 566244 461274 566296
rect 126606 566176 126612 566228
rect 126664 566216 126670 566228
rect 526438 566216 526444 566228
rect 126664 566188 526444 566216
rect 126664 566176 126670 566188
rect 526438 566176 526444 566188
rect 526496 566176 526502 566228
rect 148962 566108 148968 566160
rect 149020 566148 149026 566160
rect 551278 566148 551284 566160
rect 149020 566120 551284 566148
rect 149020 566108 149026 566120
rect 551278 566108 551284 566120
rect 551336 566108 551342 566160
rect 104250 566040 104256 566092
rect 104308 566080 104314 566092
rect 508498 566080 508504 566092
rect 104308 566052 508504 566080
rect 104308 566040 104314 566052
rect 508498 566040 508504 566052
rect 508556 566040 508562 566092
rect 58618 565972 58624 566024
rect 58676 566012 58682 566024
rect 472342 566012 472348 566024
rect 58676 565984 472348 566012
rect 58676 565972 58682 565984
rect 472342 565972 472348 565984
rect 472400 565972 472406 566024
rect 32398 565904 32404 565956
rect 32456 565944 32462 565956
rect 454034 565944 454040 565956
rect 32456 565916 454040 565944
rect 32456 565904 32462 565916
rect 454034 565904 454040 565916
rect 454092 565904 454098 565956
rect 50338 565836 50344 565888
rect 50396 565876 50402 565888
rect 494698 565876 494704 565888
rect 50396 565848 494704 565876
rect 50396 565836 50402 565848
rect 494698 565836 494704 565848
rect 494756 565836 494762 565888
rect 71038 565632 71044 565684
rect 71096 565672 71102 565684
rect 375558 565672 375564 565684
rect 71096 565644 375564 565672
rect 71096 565632 71102 565644
rect 375558 565632 375564 565644
rect 375616 565632 375622 565684
rect 208210 565564 208216 565616
rect 208268 565604 208274 565616
rect 537478 565604 537484 565616
rect 208268 565576 537484 565604
rect 208268 565564 208274 565576
rect 537478 565564 537484 565576
rect 537536 565564 537542 565616
rect 77938 565496 77944 565548
rect 77996 565536 78002 565548
rect 427952 565536 427958 565548
rect 77996 565508 427958 565536
rect 77996 565496 78002 565508
rect 427952 565496 427958 565508
rect 428010 565496 428016 565548
rect 182220 565428 182226 565480
rect 182278 565468 182284 565480
rect 536098 565468 536104 565480
rect 182278 565440 536104 565468
rect 182278 565428 182284 565440
rect 536098 565428 536104 565440
rect 536156 565428 536162 565480
rect 211936 565360 211942 565412
rect 211994 565400 212000 565412
rect 580442 565400 580448 565412
rect 211994 565372 580448 565400
rect 211994 565360 212000 565372
rect 580442 565360 580448 565372
rect 580500 565360 580506 565412
rect 160002 565292 160008 565344
rect 160060 565332 160066 565344
rect 530578 565332 530584 565344
rect 160060 565304 530584 565332
rect 160060 565292 160066 565304
rect 530578 565292 530584 565304
rect 530636 565292 530642 565344
rect 72418 565224 72424 565276
rect 72476 565264 72482 565276
rect 449986 565264 449992 565276
rect 72476 565236 449992 565264
rect 72476 565224 72482 565236
rect 449986 565224 449992 565236
rect 450044 565224 450050 565276
rect 201126 565156 201132 565208
rect 201184 565196 201190 565208
rect 580350 565196 580356 565208
rect 201184 565168 580356 565196
rect 201184 565156 201190 565168
rect 580350 565156 580356 565168
rect 580408 565156 580414 565208
rect 3786 565088 3792 565140
rect 3844 565128 3850 565140
rect 390554 565128 390560 565140
rect 3844 565100 390560 565128
rect 3844 565088 3850 565100
rect 390554 565088 390560 565100
rect 390612 565088 390618 565140
rect 137830 565020 137836 565072
rect 137888 565060 137894 565072
rect 529198 565060 529204 565072
rect 137888 565032 529204 565060
rect 137888 565020 137894 565032
rect 529198 565020 529204 565032
rect 529256 565020 529262 565072
rect 47578 564952 47584 565004
rect 47636 564992 47642 565004
rect 442534 564992 442540 565004
rect 47636 564964 442540 564992
rect 47636 564952 47642 564964
rect 442534 564952 442540 564964
rect 442592 564952 442598 565004
rect 186222 564884 186228 564936
rect 186280 564924 186286 564936
rect 580258 564924 580264 564936
rect 186280 564896 580264 564924
rect 186280 564884 186286 564896
rect 580258 564884 580264 564896
rect 580316 564884 580322 564936
rect 115474 564816 115480 564868
rect 115532 564856 115538 564868
rect 511258 564856 511264 564868
rect 115532 564828 511264 564856
rect 115532 564816 115538 564828
rect 511258 564816 511264 564828
rect 511316 564816 511322 564868
rect 3694 564748 3700 564800
rect 3752 564788 3758 564800
rect 401594 564788 401600 564800
rect 3752 564760 401600 564788
rect 3752 564748 3758 564760
rect 401594 564748 401600 564760
rect 401652 564748 401658 564800
rect 3602 564680 3608 564732
rect 3660 564720 3666 564732
rect 412818 564720 412824 564732
rect 3660 564692 412824 564720
rect 3660 564680 3666 564692
rect 412818 564680 412824 564692
rect 412876 564680 412882 564732
rect 435082 564720 435088 564732
rect 435043 564692 435088 564720
rect 435082 564680 435088 564692
rect 435140 564680 435146 564732
rect 489886 564692 499574 564720
rect 69658 564612 69664 564664
rect 69716 564652 69722 564664
rect 483566 564652 483572 564664
rect 69716 564624 483572 564652
rect 69716 564612 69722 564624
rect 483566 564612 483572 564624
rect 483624 564612 483630 564664
rect 108022 564544 108028 564596
rect 108080 564584 108086 564596
rect 489886 564584 489914 564692
rect 108080 564556 489914 564584
rect 108080 564544 108086 564556
rect 491202 564544 491208 564596
rect 491260 564544 491266 564596
rect 499546 564584 499574 564692
rect 538858 564584 538864 564596
rect 499546 564556 538864 564584
rect 538858 564544 538864 564556
rect 538916 564544 538922 564596
rect 3510 564476 3516 564528
rect 3568 564516 3574 564528
rect 435085 564519 435143 564525
rect 435085 564516 435097 564519
rect 3568 564488 435097 564516
rect 3568 564476 3574 564488
rect 435085 564485 435097 564488
rect 435131 564485 435143 564519
rect 435085 564479 435143 564485
rect 3418 564408 3424 564460
rect 3476 564448 3482 564460
rect 491220 564448 491248 564544
rect 3476 564420 491248 564448
rect 3476 564408 3482 564420
rect 3326 554684 3332 554736
rect 3384 554724 3390 554736
rect 71038 554724 71044 554736
rect 3384 554696 71044 554724
rect 3384 554684 3390 554696
rect 71038 554684 71044 554696
rect 71096 554684 71102 554736
rect 537478 538160 537484 538212
rect 537536 538200 537542 538212
rect 580166 538200 580172 538212
rect 537536 538172 580172 538200
rect 537536 538160 537542 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 3234 528504 3240 528556
rect 3292 528544 3298 528556
rect 43438 528544 43444 528556
rect 3292 528516 43444 528544
rect 3292 528504 3298 528516
rect 43438 528504 43444 528516
rect 43496 528504 43502 528556
rect 507118 511912 507124 511964
rect 507176 511952 507182 511964
rect 580166 511952 580172 511964
rect 507176 511924 580172 511952
rect 507176 511912 507182 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 3234 502256 3240 502308
rect 3292 502296 3298 502308
rect 61378 502296 61384 502308
rect 3292 502268 61384 502296
rect 3292 502256 3298 502268
rect 61378 502256 61384 502268
rect 61436 502256 61442 502308
rect 548518 485732 548524 485784
rect 548576 485772 548582 485784
rect 580166 485772 580172 485784
rect 548576 485744 580172 485772
rect 548576 485732 548582 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 3326 476008 3332 476060
rect 3384 476048 3390 476060
rect 65518 476048 65524 476060
rect 3384 476020 65524 476048
rect 3384 476008 3390 476020
rect 65518 476008 65524 476020
rect 65576 476008 65582 476060
rect 505738 458124 505744 458176
rect 505796 458164 505802 458176
rect 580166 458164 580172 458176
rect 505796 458136 580172 458164
rect 505796 458124 505802 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 53098 449868 53104 449880
rect 3384 449840 53104 449868
rect 3384 449828 3390 449840
rect 53098 449828 53104 449840
rect 53156 449828 53162 449880
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 79318 423620 79324 423632
rect 3384 423592 79324 423620
rect 3384 423580 3390 423592
rect 79318 423580 79324 423592
rect 79376 423580 79382 423632
rect 525058 419432 525064 419484
rect 525116 419472 525122 419484
rect 580166 419472 580172 419484
rect 525116 419444 580172 419472
rect 525116 419432 525122 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 536098 405628 536104 405680
rect 536156 405668 536162 405680
rect 580166 405668 580172 405680
rect 536156 405640 580172 405668
rect 536156 405628 536162 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 57238 398800 57244 398812
rect 3384 398772 57244 398800
rect 3384 398760 3390 398772
rect 57238 398760 57244 398772
rect 57296 398760 57302 398812
rect 556798 379448 556804 379500
rect 556856 379488 556862 379500
rect 580166 379488 580172 379500
rect 556856 379460 580172 379488
rect 556856 379448 556862 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 75178 372552 75184 372564
rect 3384 372524 75184 372552
rect 3384 372512 3390 372524
rect 75178 372512 75184 372524
rect 75236 372512 75242 372564
rect 522298 365644 522304 365696
rect 522356 365684 522362 365696
rect 580166 365684 580172 365696
rect 522356 365656 580172 365684
rect 522356 365644 522362 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3142 358572 3148 358624
rect 3200 358612 3206 358624
rect 7558 358612 7564 358624
rect 3200 358584 7564 358612
rect 3200 358572 3206 358584
rect 7558 358572 7564 358584
rect 7616 358572 7622 358624
rect 533338 353200 533344 353252
rect 533396 353240 533402 353252
rect 580166 353240 580172 353252
rect 533396 353212 580172 353240
rect 533396 353200 533402 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 54478 346372 54484 346384
rect 3384 346344 54484 346372
rect 3384 346332 3390 346344
rect 54478 346332 54484 346344
rect 54536 346332 54542 346384
rect 555418 325592 555424 325644
rect 555476 325632 555482 325644
rect 580166 325632 580172 325644
rect 555476 325604 580172 325632
rect 555476 325592 555482 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 77938 320124 77944 320136
rect 3384 320096 77944 320124
rect 3384 320084 3390 320096
rect 77938 320084 77944 320096
rect 77996 320084 78002 320136
rect 520918 313216 520924 313268
rect 520976 313256 520982 313268
rect 580166 313256 580172 313268
rect 520976 313228 580172 313256
rect 520976 313216 520982 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 530578 299412 530584 299464
rect 530636 299452 530642 299464
rect 580166 299452 580172 299464
rect 530636 299424 580172 299452
rect 530636 299412 530642 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 51718 293944 51724 293956
rect 3108 293916 51724 293944
rect 3108 293904 3114 293916
rect 51718 293904 51724 293916
rect 51776 293904 51782 293956
rect 547138 273164 547144 273216
rect 547196 273204 547202 273216
rect 580166 273204 580172 273216
rect 547196 273176 580172 273204
rect 547196 273164 547202 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 76558 267696 76564 267708
rect 3568 267668 76564 267696
rect 3568 267656 3574 267668
rect 76558 267656 76564 267668
rect 76616 267656 76622 267708
rect 519538 259360 519544 259412
rect 519596 259400 519602 259412
rect 580166 259400 580172 259412
rect 519596 259372 580172 259400
rect 519596 259360 519602 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 2774 254328 2780 254380
rect 2832 254368 2838 254380
rect 4890 254368 4896 254380
rect 2832 254340 4896 254368
rect 2832 254328 2838 254340
rect 4890 254328 4896 254340
rect 4948 254328 4954 254380
rect 551278 245556 551284 245608
rect 551336 245596 551342 245608
rect 580166 245596 580172 245608
rect 551336 245568 580172 245596
rect 551336 245556 551342 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 47578 241448 47584 241460
rect 3568 241420 47584 241448
rect 3568 241408 3574 241420
rect 47578 241408 47584 241420
rect 47636 241408 47642 241460
rect 544378 233180 544384 233232
rect 544436 233220 544442 233232
rect 579982 233220 579988 233232
rect 544436 233192 579988 233220
rect 544436 233180 544442 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 518158 219376 518164 219428
rect 518216 219416 518222 219428
rect 580166 219416 580172 219428
rect 518216 219388 580172 219416
rect 518216 219376 518222 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 72418 215268 72424 215280
rect 3384 215240 72424 215268
rect 3384 215228 3390 215240
rect 72418 215228 72424 215240
rect 72476 215228 72482 215280
rect 529198 206932 529204 206984
rect 529256 206972 529262 206984
rect 579798 206972 579804 206984
rect 529256 206944 579804 206972
rect 529256 206932 529262 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 2774 202716 2780 202768
rect 2832 202756 2838 202768
rect 4798 202756 4804 202768
rect 2832 202728 4804 202756
rect 2832 202716 2838 202728
rect 4798 202716 4804 202728
rect 4856 202716 4862 202768
rect 542998 193128 543004 193180
rect 543056 193168 543062 193180
rect 580166 193168 580172 193180
rect 543056 193140 580172 193168
rect 543056 193128 543062 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 32398 189020 32404 189032
rect 3568 188992 32404 189020
rect 3568 188980 3574 188992
rect 32398 188980 32404 188992
rect 32456 188980 32462 189032
rect 515398 179324 515404 179376
rect 515456 179364 515462 179376
rect 580166 179364 580172 179376
rect 515456 179336 580172 179364
rect 515456 179324 515462 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 526438 166948 526444 167000
rect 526496 166988 526502 167000
rect 580166 166988 580172 167000
rect 526496 166960 580172 166988
rect 526496 166948 526502 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 68278 164200 68284 164212
rect 3292 164172 68284 164200
rect 3292 164160 3298 164172
rect 68278 164160 68284 164172
rect 68336 164160 68342 164212
rect 540238 153144 540244 153196
rect 540296 153184 540302 153196
rect 580166 153184 580172 153196
rect 540296 153156 580172 153184
rect 540296 153144 540302 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 17218 150396 17224 150408
rect 3568 150368 17224 150396
rect 3568 150356 3574 150368
rect 17218 150356 17224 150368
rect 17276 150356 17282 150408
rect 512638 139340 512644 139392
rect 512696 139380 512702 139392
rect 580166 139380 580172 139392
rect 512696 139352 580172 139380
rect 512696 139340 512702 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 80054 138388 80060 138440
rect 80112 138428 80118 138440
rect 81020 138428 81026 138440
rect 80112 138400 81026 138428
rect 80112 138388 80118 138400
rect 81020 138388 81026 138400
rect 81078 138388 81084 138440
rect 161566 138388 161572 138440
rect 161624 138428 161630 138440
rect 162808 138428 162814 138440
rect 161624 138400 162814 138428
rect 161624 138388 161630 138400
rect 162808 138388 162814 138400
rect 162866 138388 162872 138440
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 11698 137952 11704 137964
rect 3568 137924 11704 137952
rect 3568 137912 3574 137924
rect 11698 137912 11704 137924
rect 11756 137912 11762 137964
rect 54478 136552 54484 136604
rect 54536 136592 54542 136604
rect 111978 136592 111984 136604
rect 54536 136564 111984 136592
rect 54536 136552 54542 136564
rect 111978 136552 111984 136564
rect 112036 136552 112042 136604
rect 115290 136552 115296 136604
rect 115348 136592 115354 136604
rect 117958 136592 117964 136604
rect 115348 136564 117964 136592
rect 115348 136552 115354 136564
rect 117958 136552 117964 136564
rect 118016 136552 118022 136604
rect 124122 136552 124128 136604
rect 124180 136592 124186 136604
rect 169662 136592 169668 136604
rect 124180 136564 169668 136592
rect 124180 136552 124186 136564
rect 169662 136552 169668 136564
rect 169720 136552 169726 136604
rect 170490 136552 170496 136604
rect 170548 136592 170554 136604
rect 171410 136592 171416 136604
rect 170548 136564 171416 136592
rect 170548 136552 170554 136564
rect 171410 136552 171416 136564
rect 171468 136552 171474 136604
rect 180702 136552 180708 136604
rect 180760 136592 180766 136604
rect 210970 136592 210976 136604
rect 180760 136564 210976 136592
rect 180760 136552 180766 136564
rect 210970 136552 210976 136564
rect 211028 136552 211034 136604
rect 213822 136552 213828 136604
rect 213880 136592 213886 136604
rect 235074 136592 235080 136604
rect 213880 136564 235080 136592
rect 213880 136552 213886 136564
rect 235074 136552 235080 136564
rect 235132 136552 235138 136604
rect 238018 136552 238024 136604
rect 238076 136592 238082 136604
rect 250622 136592 250628 136604
rect 238076 136564 250628 136592
rect 238076 136552 238082 136564
rect 250622 136552 250628 136564
rect 250680 136552 250686 136604
rect 274542 136552 274548 136604
rect 274600 136592 274606 136604
rect 279050 136592 279056 136604
rect 274600 136564 279056 136592
rect 274600 136552 274606 136564
rect 279050 136552 279056 136564
rect 279108 136552 279114 136604
rect 315298 136552 315304 136604
rect 315356 136592 315362 136604
rect 316678 136592 316684 136604
rect 315356 136564 316684 136592
rect 315356 136552 315362 136564
rect 316678 136552 316684 136564
rect 316736 136552 316742 136604
rect 403986 136552 403992 136604
rect 404044 136592 404050 136604
rect 435358 136592 435364 136604
rect 404044 136564 435364 136592
rect 404044 136552 404050 136564
rect 435358 136552 435364 136564
rect 435416 136552 435422 136604
rect 456061 136595 456119 136601
rect 456061 136561 456073 136595
rect 456107 136592 456119 136595
rect 496817 136595 496875 136601
rect 496817 136592 496829 136595
rect 456107 136564 496829 136592
rect 456107 136561 456119 136564
rect 456061 136555 456119 136561
rect 496817 136561 496829 136564
rect 496863 136561 496875 136595
rect 496817 136555 496875 136561
rect 68278 136484 68284 136536
rect 68336 136524 68342 136536
rect 125778 136524 125784 136536
rect 68336 136496 125784 136524
rect 68336 136484 68342 136496
rect 125778 136484 125784 136496
rect 125836 136484 125842 136536
rect 126238 136484 126244 136536
rect 126296 136524 126302 136536
rect 136082 136524 136088 136536
rect 126296 136496 136088 136524
rect 126296 136484 126302 136496
rect 136082 136484 136088 136496
rect 136140 136484 136146 136536
rect 142798 136484 142804 136536
rect 142856 136524 142862 136536
rect 172238 136524 172244 136536
rect 142856 136496 172244 136524
rect 142856 136484 142862 136496
rect 172238 136484 172244 136496
rect 172296 136484 172302 136536
rect 173802 136484 173808 136536
rect 173860 136524 173866 136536
rect 173860 136496 174124 136524
rect 173860 136484 173866 136496
rect 74442 136416 74448 136468
rect 74500 136456 74506 136468
rect 133506 136456 133512 136468
rect 74500 136428 133512 136456
rect 74500 136416 74506 136428
rect 133506 136416 133512 136428
rect 133564 136416 133570 136468
rect 170398 136416 170404 136468
rect 170456 136456 170462 136468
rect 173986 136456 173992 136468
rect 170456 136428 173992 136456
rect 170456 136416 170462 136428
rect 173986 136416 173992 136428
rect 174044 136416 174050 136468
rect 174096 136456 174124 136496
rect 177850 136484 177856 136536
rect 177908 136524 177914 136536
rect 209314 136524 209320 136536
rect 177908 136496 209320 136524
rect 177908 136484 177914 136496
rect 209314 136484 209320 136496
rect 209372 136484 209378 136536
rect 215202 136484 215208 136536
rect 215260 136524 215266 136536
rect 235994 136524 236000 136536
rect 215260 136496 236000 136524
rect 215260 136484 215266 136496
rect 235994 136484 236000 136496
rect 236052 136484 236058 136536
rect 238662 136484 238668 136536
rect 238720 136524 238726 136536
rect 253198 136524 253204 136536
rect 238720 136496 253204 136524
rect 238720 136484 238726 136496
rect 253198 136484 253204 136496
rect 253256 136484 253262 136536
rect 255958 136484 255964 136536
rect 256016 136524 256022 136536
rect 263502 136524 263508 136536
rect 256016 136496 263508 136524
rect 256016 136484 256022 136496
rect 263502 136484 263508 136496
rect 263560 136484 263566 136536
rect 303246 136484 303252 136536
rect 303304 136524 303310 136536
rect 306558 136524 306564 136536
rect 303304 136496 306564 136524
rect 303304 136484 303310 136496
rect 306558 136484 306564 136496
rect 306616 136484 306622 136536
rect 398742 136484 398748 136536
rect 398800 136524 398806 136536
rect 429746 136524 429752 136536
rect 398800 136496 429752 136524
rect 398800 136484 398806 136496
rect 429746 136484 429752 136496
rect 429804 136484 429810 136536
rect 441062 136484 441068 136536
rect 441120 136524 441126 136536
rect 443638 136524 443644 136536
rect 441120 136496 443644 136524
rect 441120 136484 441126 136496
rect 443638 136484 443644 136496
rect 443696 136484 443702 136536
rect 449618 136484 449624 136536
rect 449676 136524 449682 136536
rect 506474 136524 506480 136536
rect 449676 136496 506480 136524
rect 449676 136484 449682 136496
rect 506474 136484 506480 136496
rect 506532 136484 506538 136536
rect 205818 136456 205824 136468
rect 174096 136428 205824 136456
rect 205818 136416 205824 136428
rect 205876 136416 205882 136468
rect 211062 136416 211068 136468
rect 211120 136456 211126 136468
rect 233418 136456 233424 136468
rect 211120 136428 233424 136456
rect 211120 136416 211126 136428
rect 233418 136416 233424 136428
rect 233476 136416 233482 136468
rect 235902 136416 235908 136468
rect 235960 136456 235966 136468
rect 251450 136456 251456 136468
rect 235960 136428 251456 136456
rect 235960 136416 235966 136428
rect 251450 136416 251456 136428
rect 251508 136416 251514 136468
rect 256602 136416 256608 136468
rect 256660 136456 256666 136468
rect 266078 136456 266084 136468
rect 256660 136428 266084 136456
rect 256660 136416 256666 136428
rect 266078 136416 266084 136428
rect 266136 136416 266142 136468
rect 286962 136416 286968 136468
rect 287020 136456 287026 136468
rect 288526 136456 288532 136468
rect 287020 136428 288532 136456
rect 287020 136416 287026 136428
rect 288526 136416 288532 136428
rect 288584 136416 288590 136468
rect 393682 136416 393688 136468
rect 393740 136456 393746 136468
rect 429930 136456 429936 136468
rect 393740 136428 429936 136456
rect 393740 136416 393746 136428
rect 429930 136416 429936 136428
rect 429988 136416 429994 136468
rect 453942 136416 453948 136468
rect 454000 136456 454006 136468
rect 461213 136459 461271 136465
rect 454000 136428 456794 136456
rect 454000 136416 454006 136428
rect 78490 136348 78496 136400
rect 78548 136388 78554 136400
rect 136910 136388 136916 136400
rect 78548 136360 136916 136388
rect 78548 136348 78554 136360
rect 136910 136348 136916 136360
rect 136968 136348 136974 136400
rect 140774 136348 140780 136400
rect 140832 136388 140838 136400
rect 145558 136388 145564 136400
rect 140832 136360 145564 136388
rect 140832 136348 140838 136360
rect 145558 136348 145564 136360
rect 145616 136348 145622 136400
rect 169570 136348 169576 136400
rect 169628 136388 169634 136400
rect 203242 136388 203248 136400
rect 169628 136360 203248 136388
rect 169628 136348 169634 136360
rect 203242 136348 203248 136360
rect 203300 136348 203306 136400
rect 204898 136348 204904 136400
rect 204956 136388 204962 136400
rect 228266 136388 228272 136400
rect 204956 136360 228272 136388
rect 204956 136348 204962 136360
rect 228266 136348 228272 136360
rect 228324 136348 228330 136400
rect 229002 136348 229008 136400
rect 229060 136388 229066 136400
rect 246298 136388 246304 136400
rect 229060 136360 246304 136388
rect 229060 136348 229066 136360
rect 246298 136348 246304 136360
rect 246356 136348 246362 136400
rect 251082 136348 251088 136400
rect 251140 136388 251146 136400
rect 261846 136388 261852 136400
rect 251140 136360 261852 136388
rect 251140 136348 251146 136360
rect 261846 136348 261852 136360
rect 261904 136348 261910 136400
rect 395430 136348 395436 136400
rect 395488 136388 395494 136400
rect 427081 136391 427139 136397
rect 427081 136388 427093 136391
rect 395488 136360 427093 136388
rect 395488 136348 395494 136360
rect 427081 136357 427093 136360
rect 427127 136357 427139 136391
rect 427081 136351 427139 136357
rect 444466 136348 444472 136400
rect 444524 136388 444530 136400
rect 456061 136391 456119 136397
rect 456061 136388 456073 136391
rect 444524 136360 456073 136388
rect 444524 136348 444530 136360
rect 456061 136357 456073 136360
rect 456107 136357 456119 136391
rect 456766 136388 456794 136428
rect 461213 136425 461225 136459
rect 461259 136456 461271 136459
rect 508590 136456 508596 136468
rect 461259 136428 508596 136456
rect 461259 136425 461271 136428
rect 461213 136419 461271 136425
rect 508590 136416 508596 136428
rect 508648 136416 508654 136468
rect 511350 136388 511356 136400
rect 456766 136360 511356 136388
rect 456061 136351 456119 136357
rect 511350 136348 511356 136360
rect 511408 136348 511414 136400
rect 71682 136280 71688 136332
rect 71740 136320 71746 136332
rect 131758 136320 131764 136332
rect 71740 136292 131764 136320
rect 71740 136280 71746 136292
rect 131758 136280 131764 136292
rect 131816 136280 131822 136332
rect 144178 136280 144184 136332
rect 144236 136320 144242 136332
rect 181714 136320 181720 136332
rect 144236 136292 181720 136320
rect 144236 136280 144242 136292
rect 181714 136280 181720 136292
rect 181772 136280 181778 136332
rect 186958 136280 186964 136332
rect 187016 136320 187022 136332
rect 192018 136320 192024 136332
rect 187016 136292 192024 136320
rect 187016 136280 187022 136292
rect 192018 136280 192024 136292
rect 192076 136280 192082 136332
rect 195241 136323 195299 136329
rect 195241 136289 195253 136323
rect 195287 136320 195299 136323
rect 216214 136320 216220 136332
rect 195287 136292 216220 136320
rect 195287 136289 195299 136292
rect 195241 136283 195299 136289
rect 216214 136280 216220 136292
rect 216272 136280 216278 136332
rect 216582 136280 216588 136332
rect 216640 136320 216646 136332
rect 236822 136320 236828 136332
rect 216640 136292 236828 136320
rect 216640 136280 216646 136292
rect 236822 136280 236828 136292
rect 236880 136280 236886 136332
rect 237282 136280 237288 136332
rect 237340 136320 237346 136332
rect 252370 136320 252376 136332
rect 237340 136292 252376 136320
rect 237340 136280 237346 136292
rect 252370 136280 252376 136292
rect 252428 136280 252434 136332
rect 253842 136280 253848 136332
rect 253900 136320 253906 136332
rect 264422 136320 264428 136332
rect 253900 136292 264428 136320
rect 253900 136280 253906 136292
rect 264422 136280 264428 136292
rect 264480 136280 264486 136332
rect 267642 136280 267648 136332
rect 267700 136320 267706 136332
rect 273898 136320 273904 136332
rect 267700 136292 273904 136320
rect 267700 136280 267706 136292
rect 273898 136280 273904 136292
rect 273956 136280 273962 136332
rect 400582 136280 400588 136332
rect 400640 136320 400646 136332
rect 440234 136320 440240 136332
rect 400640 136292 440240 136320
rect 400640 136280 400646 136292
rect 440234 136280 440240 136292
rect 440292 136280 440298 136332
rect 451366 136280 451372 136332
rect 451424 136320 451430 136332
rect 461213 136323 461271 136329
rect 461213 136320 461225 136323
rect 451424 136292 461225 136320
rect 451424 136280 451430 136292
rect 461213 136289 461225 136292
rect 461259 136289 461271 136323
rect 461213 136283 461271 136289
rect 475381 136323 475439 136329
rect 475381 136289 475393 136323
rect 475427 136320 475439 136323
rect 529198 136320 529204 136332
rect 475427 136292 529204 136320
rect 475427 136289 475439 136292
rect 475381 136283 475439 136289
rect 529198 136280 529204 136292
rect 529256 136280 529262 136332
rect 51718 136212 51724 136264
rect 51776 136252 51782 136264
rect 115382 136252 115388 136264
rect 51776 136224 115388 136252
rect 51776 136212 51782 136224
rect 115382 136212 115388 136224
rect 115440 136212 115446 136264
rect 117222 136212 117228 136264
rect 117280 136252 117286 136264
rect 164510 136252 164516 136264
rect 117280 136224 164516 136252
rect 117280 136212 117286 136224
rect 164510 136212 164516 136224
rect 164568 136212 164574 136264
rect 166902 136212 166908 136264
rect 166960 136252 166966 136264
rect 200666 136252 200672 136264
rect 166960 136224 200672 136252
rect 166960 136212 166966 136224
rect 200666 136212 200672 136224
rect 200724 136212 200730 136264
rect 202782 136212 202788 136264
rect 202840 136252 202846 136264
rect 226518 136252 226524 136264
rect 202840 136224 226524 136252
rect 202840 136212 202846 136224
rect 226518 136212 226524 136224
rect 226576 136212 226582 136264
rect 227622 136212 227628 136264
rect 227680 136252 227686 136264
rect 244550 136252 244556 136264
rect 227680 136224 244556 136252
rect 227680 136212 227686 136224
rect 244550 136212 244556 136224
rect 244608 136212 244614 136264
rect 246942 136212 246948 136264
rect 247000 136252 247006 136264
rect 259270 136252 259276 136264
rect 247000 136224 259276 136252
rect 247000 136212 247006 136224
rect 259270 136212 259276 136224
rect 259328 136212 259334 136264
rect 263502 136212 263508 136264
rect 263560 136252 263566 136264
rect 267185 136255 267243 136261
rect 263560 136224 267136 136252
rect 263560 136212 263566 136224
rect 29638 136144 29644 136196
rect 29696 136184 29702 136196
rect 93026 136184 93032 136196
rect 29696 136156 93032 136184
rect 29696 136144 29702 136156
rect 93026 136144 93032 136156
rect 93084 136144 93090 136196
rect 104158 136144 104164 136196
rect 104216 136184 104222 136196
rect 109402 136184 109408 136196
rect 104216 136156 109408 136184
rect 104216 136144 104222 136156
rect 109402 136144 109408 136156
rect 109460 136144 109466 136196
rect 113082 136144 113088 136196
rect 113140 136184 113146 136196
rect 161934 136184 161940 136196
rect 113140 136156 161940 136184
rect 113140 136144 113146 136156
rect 161934 136144 161940 136156
rect 161992 136144 161998 136196
rect 162762 136144 162768 136196
rect 162820 136184 162826 136196
rect 198090 136184 198096 136196
rect 162820 136156 198096 136184
rect 162820 136144 162826 136156
rect 198090 136144 198096 136156
rect 198148 136144 198154 136196
rect 205542 136144 205548 136196
rect 205600 136184 205606 136196
rect 229094 136184 229100 136196
rect 205600 136156 229100 136184
rect 205600 136144 205606 136156
rect 229094 136144 229100 136156
rect 229152 136144 229158 136196
rect 234522 136144 234528 136196
rect 234580 136184 234586 136196
rect 249794 136184 249800 136196
rect 234580 136156 249800 136184
rect 234580 136144 234586 136156
rect 249794 136144 249800 136156
rect 249852 136144 249858 136196
rect 252462 136144 252468 136196
rect 252520 136184 252526 136196
rect 262674 136184 262680 136196
rect 252520 136156 262680 136184
rect 252520 136144 252526 136156
rect 262674 136144 262680 136156
rect 262732 136144 262738 136196
rect 264238 136144 264244 136196
rect 264296 136184 264302 136196
rect 266998 136184 267004 136196
rect 264296 136156 267004 136184
rect 264296 136144 264302 136156
rect 266998 136144 267004 136156
rect 267056 136144 267062 136196
rect 267108 136184 267136 136224
rect 267185 136221 267197 136255
rect 267231 136252 267243 136255
rect 268746 136252 268752 136264
rect 267231 136224 268752 136252
rect 267231 136221 267243 136224
rect 267185 136215 267243 136221
rect 268746 136212 268752 136224
rect 268804 136212 268810 136264
rect 448514 136252 448520 136264
rect 408466 136224 448520 136252
rect 271322 136184 271328 136196
rect 267108 136156 271328 136184
rect 271322 136144 271328 136156
rect 271380 136144 271386 136196
rect 276658 136144 276664 136196
rect 276716 136184 276722 136196
rect 279878 136184 279884 136196
rect 276716 136156 279884 136184
rect 276716 136144 276722 136156
rect 279878 136144 279884 136156
rect 279936 136144 279942 136196
rect 391106 136144 391112 136196
rect 391164 136184 391170 136196
rect 399478 136184 399484 136196
rect 391164 136156 399484 136184
rect 391164 136144 391170 136156
rect 399478 136144 399484 136156
rect 399536 136144 399542 136196
rect 407482 136144 407488 136196
rect 407540 136184 407546 136196
rect 408466 136184 408494 136224
rect 448514 136212 448520 136224
rect 448572 136212 448578 136264
rect 457438 136212 457444 136264
rect 457496 136252 457502 136264
rect 517514 136252 517520 136264
rect 457496 136224 517520 136252
rect 457496 136212 457502 136224
rect 517514 136212 517520 136224
rect 517572 136212 517578 136264
rect 407540 136156 408494 136184
rect 407540 136144 407546 136156
rect 409138 136144 409144 136196
rect 409196 136184 409202 136196
rect 450446 136184 450452 136196
rect 409196 136156 450452 136184
rect 409196 136144 409202 136156
rect 450446 136144 450452 136156
rect 450504 136144 450510 136196
rect 456518 136144 456524 136196
rect 456576 136184 456582 136196
rect 464246 136184 464252 136196
rect 456576 136156 464252 136184
rect 456576 136144 456582 136156
rect 464246 136144 464252 136156
rect 464304 136144 464310 136196
rect 469490 136144 469496 136196
rect 469548 136184 469554 136196
rect 475381 136187 475439 136193
rect 475381 136184 475393 136187
rect 469548 136156 475393 136184
rect 469548 136144 469554 136156
rect 475381 136153 475393 136156
rect 475427 136153 475439 136187
rect 475381 136147 475439 136153
rect 482370 136144 482376 136196
rect 482428 136184 482434 136196
rect 542998 136184 543004 136196
rect 482428 136156 543004 136184
rect 482428 136144 482434 136156
rect 542998 136144 543004 136156
rect 543056 136144 543062 136196
rect 32398 136076 32404 136128
rect 32456 136116 32462 136128
rect 99006 136116 99012 136128
rect 32456 136088 99012 136116
rect 32456 136076 32462 136088
rect 99006 136076 99012 136088
rect 99064 136076 99070 136128
rect 107562 136076 107568 136128
rect 107620 136116 107626 136128
rect 157610 136116 157616 136128
rect 107620 136088 157616 136116
rect 107620 136076 107626 136088
rect 157610 136076 157616 136088
rect 157668 136076 157674 136128
rect 160002 136076 160008 136128
rect 160060 136116 160066 136128
rect 195514 136116 195520 136128
rect 160060 136088 195520 136116
rect 160060 136076 160066 136088
rect 195514 136076 195520 136088
rect 195572 136076 195578 136128
rect 202690 136076 202696 136128
rect 202748 136116 202754 136128
rect 227346 136116 227352 136128
rect 202748 136088 227352 136116
rect 202748 136076 202754 136088
rect 227346 136076 227352 136088
rect 227404 136076 227410 136128
rect 227530 136076 227536 136128
rect 227588 136116 227594 136128
rect 245470 136116 245476 136128
rect 227588 136088 245476 136116
rect 227588 136076 227594 136088
rect 245470 136076 245476 136088
rect 245528 136076 245534 136128
rect 249702 136076 249708 136128
rect 249760 136116 249766 136128
rect 260926 136116 260932 136128
rect 249760 136088 260932 136116
rect 249760 136076 249766 136088
rect 260926 136076 260932 136088
rect 260984 136076 260990 136128
rect 264882 136076 264888 136128
rect 264940 136116 264946 136128
rect 272150 136116 272156 136128
rect 264940 136088 272156 136116
rect 264940 136076 264946 136088
rect 272150 136076 272156 136088
rect 272208 136076 272214 136128
rect 273898 136076 273904 136128
rect 273956 136116 273962 136128
rect 278222 136116 278228 136128
rect 273956 136088 278228 136116
rect 273956 136076 273962 136088
rect 278222 136076 278228 136088
rect 278280 136076 278286 136128
rect 385954 136076 385960 136128
rect 386012 136116 386018 136128
rect 407758 136116 407764 136128
rect 386012 136088 407764 136116
rect 386012 136076 386018 136088
rect 407758 136076 407764 136088
rect 407816 136076 407822 136128
rect 468478 136116 468484 136128
rect 423048 136088 468484 136116
rect 17218 136008 17224 136060
rect 17276 136048 17282 136060
rect 87874 136048 87880 136060
rect 17276 136020 87880 136048
rect 17276 136008 17282 136020
rect 87874 136008 87880 136020
rect 87932 136008 87938 136060
rect 93762 136008 93768 136060
rect 93820 136048 93826 136060
rect 147306 136048 147312 136060
rect 93820 136020 147312 136048
rect 93820 136008 93826 136020
rect 147306 136008 147312 136020
rect 147364 136008 147370 136060
rect 148962 136008 148968 136060
rect 149020 136008 149026 136060
rect 153102 136008 153108 136060
rect 153160 136048 153166 136060
rect 185581 136051 185639 136057
rect 185581 136048 185593 136051
rect 153160 136020 185593 136048
rect 153160 136008 153166 136020
rect 185581 136017 185593 136020
rect 185627 136017 185639 136051
rect 185581 136011 185639 136017
rect 187602 136008 187608 136060
rect 187660 136048 187666 136060
rect 195241 136051 195299 136057
rect 195241 136048 195253 136051
rect 187660 136020 195253 136048
rect 187660 136008 187666 136020
rect 195241 136017 195253 136020
rect 195287 136017 195299 136051
rect 195241 136011 195299 136017
rect 198642 136008 198648 136060
rect 198700 136048 198706 136060
rect 223942 136048 223948 136060
rect 198700 136020 223948 136048
rect 198700 136008 198706 136020
rect 223942 136008 223948 136020
rect 224000 136008 224006 136060
rect 224862 136008 224868 136060
rect 224920 136048 224926 136060
rect 242894 136048 242900 136060
rect 224920 136020 242900 136048
rect 224920 136008 224926 136020
rect 242894 136008 242900 136020
rect 242952 136008 242958 136060
rect 245562 136008 245568 136060
rect 245620 136048 245626 136060
rect 258350 136048 258356 136060
rect 245620 136020 258356 136048
rect 245620 136008 245626 136020
rect 258350 136008 258356 136020
rect 258408 136008 258414 136060
rect 259362 136008 259368 136060
rect 259420 136048 259426 136060
rect 267826 136048 267832 136060
rect 259420 136020 267832 136048
rect 259420 136008 259426 136020
rect 267826 136008 267832 136020
rect 267884 136008 267890 136060
rect 271782 136008 271788 136060
rect 271840 136048 271846 136060
rect 277302 136048 277308 136060
rect 271840 136020 277308 136048
rect 271840 136008 271846 136020
rect 277302 136008 277308 136020
rect 277360 136008 277366 136060
rect 372982 136008 372988 136060
rect 373040 136048 373046 136060
rect 395338 136048 395344 136060
rect 373040 136020 395344 136048
rect 373040 136008 373046 136020
rect 395338 136008 395344 136020
rect 395396 136008 395402 136060
rect 414382 136008 414388 136060
rect 414440 136048 414446 136060
rect 422941 136051 422999 136057
rect 422941 136048 422953 136051
rect 414440 136020 422953 136048
rect 414440 136008 414446 136020
rect 422941 136017 422953 136020
rect 422987 136017 422999 136051
rect 422941 136011 422999 136017
rect 18598 135940 18604 135992
rect 18656 135980 18662 135992
rect 92198 135980 92204 135992
rect 18656 135952 92204 135980
rect 18656 135940 18662 135952
rect 92198 135940 92204 135952
rect 92256 135940 92262 135992
rect 95050 135940 95056 135992
rect 95108 135980 95114 135992
rect 148980 135980 149008 136008
rect 95108 135952 149008 135980
rect 95108 135940 95114 135952
rect 153010 135940 153016 135992
rect 153068 135980 153074 135992
rect 190365 135983 190423 135989
rect 190365 135980 190377 135983
rect 153068 135952 190377 135980
rect 153068 135940 153074 135952
rect 190365 135949 190377 135952
rect 190411 135949 190423 135983
rect 190365 135943 190423 135949
rect 195330 135940 195336 135992
rect 195388 135980 195394 135992
rect 221366 135980 221372 135992
rect 195388 135952 221372 135980
rect 195388 135940 195394 135952
rect 221366 135940 221372 135952
rect 221424 135940 221430 135992
rect 223482 135940 223488 135992
rect 223540 135980 223546 135992
rect 241974 135980 241980 135992
rect 223540 135952 241980 135980
rect 223540 135940 223546 135952
rect 241974 135940 241980 135952
rect 242032 135940 242038 135992
rect 242802 135940 242808 135992
rect 242860 135980 242866 135992
rect 255774 135980 255780 135992
rect 242860 135952 255780 135980
rect 242860 135940 242866 135952
rect 255774 135940 255780 135952
rect 255832 135940 255838 135992
rect 265250 135980 265256 135992
rect 258046 135952 265256 135980
rect 7558 135872 7564 135924
rect 7616 135912 7622 135924
rect 83550 135912 83556 135924
rect 7616 135884 83556 135912
rect 7616 135872 7622 135884
rect 83550 135872 83556 135884
rect 83608 135872 83614 135924
rect 88242 135872 88248 135924
rect 88300 135912 88306 135924
rect 143810 135912 143816 135924
rect 88300 135884 143816 135912
rect 88300 135872 88306 135884
rect 143810 135872 143816 135884
rect 143868 135872 143874 135924
rect 148962 135872 148968 135924
rect 149020 135912 149026 135924
rect 187786 135912 187792 135924
rect 149020 135884 187792 135912
rect 149020 135872 149026 135884
rect 187786 135872 187792 135884
rect 187844 135872 187850 135924
rect 191742 135872 191748 135924
rect 191800 135912 191806 135924
rect 218790 135912 218796 135924
rect 191800 135884 218796 135912
rect 191800 135872 191806 135884
rect 218790 135872 218796 135884
rect 218848 135872 218854 135924
rect 219989 135915 220047 135921
rect 219989 135881 220001 135915
rect 220035 135912 220047 135915
rect 222194 135912 222200 135924
rect 220035 135884 222200 135912
rect 220035 135881 220047 135884
rect 219989 135875 220047 135881
rect 222194 135872 222200 135884
rect 222252 135872 222258 135924
rect 222289 135915 222347 135921
rect 222289 135881 222301 135915
rect 222335 135912 222347 135915
rect 240318 135912 240324 135924
rect 222335 135884 240324 135912
rect 222335 135881 222347 135884
rect 222289 135875 222347 135881
rect 240318 135872 240324 135884
rect 240376 135872 240382 135924
rect 241422 135872 241428 135924
rect 241480 135912 241486 135924
rect 254946 135912 254952 135924
rect 241480 135884 254952 135912
rect 241480 135872 241486 135884
rect 254946 135872 254952 135884
rect 255004 135872 255010 135924
rect 255222 135872 255228 135924
rect 255280 135912 255286 135924
rect 258046 135912 258074 135952
rect 265250 135940 265256 135952
rect 265308 135940 265314 135992
rect 266998 135940 267004 135992
rect 267056 135980 267062 135992
rect 270402 135980 270408 135992
rect 267056 135952 270408 135980
rect 267056 135940 267062 135952
rect 270402 135940 270408 135952
rect 270460 135940 270466 135992
rect 305822 135940 305828 135992
rect 305880 135980 305886 135992
rect 309226 135980 309232 135992
rect 305880 135952 309232 135980
rect 305880 135940 305886 135952
rect 309226 135940 309232 135952
rect 309284 135940 309290 135992
rect 314470 135940 314476 135992
rect 314528 135980 314534 135992
rect 321646 135980 321652 135992
rect 314528 135952 321652 135980
rect 314528 135940 314534 135952
rect 321646 135940 321652 135952
rect 321704 135940 321710 135992
rect 335998 135940 336004 135992
rect 336056 135980 336062 135992
rect 336642 135980 336648 135992
rect 336056 135952 336648 135980
rect 336056 135940 336062 135952
rect 336642 135940 336648 135952
rect 336700 135940 336706 135992
rect 365254 135940 365260 135992
rect 365312 135980 365318 135992
rect 385678 135980 385684 135992
rect 365312 135952 385684 135980
rect 365312 135940 365318 135952
rect 385678 135940 385684 135952
rect 385736 135940 385742 135992
rect 391842 135940 391848 135992
rect 391900 135980 391906 135992
rect 414658 135980 414664 135992
rect 391900 135952 414664 135980
rect 391900 135940 391906 135952
rect 414658 135940 414664 135952
rect 414716 135940 414722 135992
rect 416958 135940 416964 135992
rect 417016 135980 417022 135992
rect 417016 135952 422064 135980
rect 417016 135940 417022 135952
rect 255280 135884 258074 135912
rect 255280 135872 255286 135884
rect 260742 135872 260748 135924
rect 260800 135912 260806 135924
rect 267185 135915 267243 135921
rect 267185 135912 267197 135915
rect 260800 135884 267197 135912
rect 260800 135872 260806 135884
rect 267185 135881 267197 135884
rect 267231 135881 267243 135915
rect 267185 135875 267243 135881
rect 277302 135872 277308 135924
rect 277360 135912 277366 135924
rect 281626 135912 281632 135924
rect 277360 135884 281632 135912
rect 277360 135872 277366 135884
rect 281626 135872 281632 135884
rect 281684 135872 281690 135924
rect 333422 135872 333428 135924
rect 333480 135912 333486 135924
rect 336090 135912 336096 135924
rect 333480 135884 336096 135912
rect 333480 135872 333486 135884
rect 336090 135872 336096 135884
rect 336148 135872 336154 135924
rect 352374 135872 352380 135924
rect 352432 135912 352438 135924
rect 374086 135912 374092 135924
rect 352432 135884 374092 135912
rect 352432 135872 352438 135884
rect 374086 135872 374092 135884
rect 374144 135872 374150 135924
rect 378042 135872 378048 135924
rect 378100 135912 378106 135924
rect 400858 135912 400864 135924
rect 378100 135884 400864 135912
rect 378100 135872 378106 135884
rect 400858 135872 400864 135884
rect 400916 135872 400922 135924
rect 402330 135872 402336 135924
rect 402388 135912 402394 135924
rect 421558 135912 421564 135924
rect 402388 135884 421564 135912
rect 402388 135872 402394 135884
rect 421558 135872 421564 135884
rect 421616 135872 421622 135924
rect 422036 135912 422064 135952
rect 422110 135940 422116 135992
rect 422168 135980 422174 135992
rect 423048 135980 423076 136088
rect 468478 136076 468484 136088
rect 468536 136076 468542 136128
rect 474642 136076 474648 136128
rect 474700 136116 474706 136128
rect 536098 136116 536104 136128
rect 474700 136088 536104 136116
rect 474700 136076 474706 136088
rect 536098 136076 536104 136088
rect 536156 136076 536162 136128
rect 423125 136051 423183 136057
rect 423125 136017 423137 136051
rect 423171 136048 423183 136051
rect 457530 136048 457536 136060
rect 423171 136020 457536 136048
rect 423171 136017 423183 136020
rect 423125 136011 423183 136017
rect 457530 136008 457536 136020
rect 457588 136008 457594 136060
rect 462590 136008 462596 136060
rect 462648 136048 462654 136060
rect 524414 136048 524420 136060
rect 462648 136020 524420 136048
rect 462648 136008 462654 136020
rect 524414 136008 524420 136020
rect 524472 136008 524478 136060
rect 461578 135980 461584 135992
rect 422168 135952 423076 135980
rect 426636 135952 461584 135980
rect 422168 135940 422174 135952
rect 426636 135912 426664 135952
rect 461578 135940 461584 135952
rect 461636 135940 461642 135992
rect 467742 135940 467748 135992
rect 467800 135980 467806 135992
rect 531314 135980 531320 135992
rect 467800 135952 531320 135980
rect 467800 135940 467806 135952
rect 531314 135940 531320 135952
rect 531372 135940 531378 135992
rect 471238 135912 471244 135924
rect 422036 135884 426664 135912
rect 427004 135884 471244 135912
rect 81342 135804 81348 135856
rect 81400 135844 81406 135856
rect 138658 135844 138664 135856
rect 81400 135816 138664 135844
rect 81400 135804 81406 135816
rect 138658 135804 138664 135816
rect 138716 135804 138722 135856
rect 146938 135804 146944 135856
rect 146996 135844 147002 135856
rect 176562 135844 176568 135856
rect 146996 135816 176568 135844
rect 146996 135804 147002 135816
rect 176562 135804 176568 135816
rect 176620 135804 176626 135856
rect 177942 135804 177948 135856
rect 178000 135844 178006 135856
rect 208394 135844 208400 135856
rect 178000 135816 208400 135844
rect 178000 135804 178006 135816
rect 208394 135804 208400 135816
rect 208452 135804 208458 135856
rect 209682 135804 209688 135856
rect 209740 135844 209746 135856
rect 231670 135844 231676 135856
rect 209740 135816 231676 135844
rect 209740 135804 209746 135816
rect 231670 135804 231676 135816
rect 231728 135804 231734 135856
rect 231762 135804 231768 135856
rect 231820 135844 231826 135856
rect 248046 135844 248052 135856
rect 231820 135816 248052 135844
rect 231820 135804 231826 135816
rect 248046 135804 248052 135816
rect 248104 135804 248110 135856
rect 260650 135804 260656 135856
rect 260708 135844 260714 135856
rect 269574 135844 269580 135856
rect 260708 135816 269580 135844
rect 260708 135804 260714 135816
rect 269574 135804 269580 135816
rect 269632 135804 269638 135856
rect 399662 135804 399668 135856
rect 399720 135844 399726 135856
rect 417418 135844 417424 135856
rect 399720 135816 417424 135844
rect 399720 135804 399726 135816
rect 417418 135804 417424 135816
rect 417476 135804 417482 135856
rect 424686 135804 424692 135856
rect 424744 135844 424750 135856
rect 427004 135844 427032 135884
rect 471238 135872 471244 135884
rect 471296 135872 471302 135924
rect 472894 135872 472900 135924
rect 472952 135912 472958 135924
rect 539594 135912 539600 135924
rect 472952 135884 539600 135912
rect 472952 135872 472958 135884
rect 539594 135872 539600 135884
rect 539652 135872 539658 135924
rect 424744 135816 427032 135844
rect 427081 135847 427139 135853
rect 424744 135804 424750 135816
rect 427081 135813 427093 135847
rect 427127 135844 427139 135847
rect 431954 135844 431960 135856
rect 427127 135816 431960 135844
rect 427127 135813 427139 135816
rect 427081 135807 427139 135813
rect 431954 135804 431960 135816
rect 432012 135804 432018 135856
rect 434990 135804 434996 135856
rect 435048 135844 435054 135856
rect 480441 135847 480499 135853
rect 480441 135844 480453 135847
rect 435048 135816 480453 135844
rect 435048 135804 435054 135816
rect 480441 135813 480453 135816
rect 480487 135813 480499 135847
rect 486418 135844 486424 135856
rect 480441 135807 480499 135813
rect 480548 135816 486424 135844
rect 65518 135736 65524 135788
rect 65576 135776 65582 135788
rect 120534 135776 120540 135788
rect 65576 135748 120540 135776
rect 65576 135736 65582 135748
rect 120534 135736 120540 135748
rect 120592 135736 120598 135788
rect 125502 135736 125508 135788
rect 125560 135776 125566 135788
rect 170582 135776 170588 135788
rect 125560 135748 170588 135776
rect 125560 135736 125566 135748
rect 170582 135736 170588 135748
rect 170640 135736 170646 135788
rect 185581 135779 185639 135785
rect 185581 135745 185593 135779
rect 185627 135776 185639 135779
rect 190270 135776 190276 135788
rect 185627 135748 190276 135776
rect 185627 135745 185639 135748
rect 185581 135739 185639 135745
rect 190270 135736 190276 135748
rect 190328 135736 190334 135788
rect 190365 135779 190423 135785
rect 190365 135745 190377 135779
rect 190411 135776 190423 135779
rect 191190 135776 191196 135788
rect 190411 135748 191196 135776
rect 190411 135745 190423 135748
rect 190365 135739 190423 135745
rect 191190 135736 191196 135748
rect 191248 135736 191254 135788
rect 200669 135779 200727 135785
rect 200669 135745 200681 135779
rect 200715 135776 200727 135779
rect 204990 135776 204996 135788
rect 200715 135748 204996 135776
rect 200715 135745 200727 135748
rect 200669 135739 200727 135745
rect 204990 135736 204996 135748
rect 205048 135736 205054 135788
rect 213178 135736 213184 135788
rect 213236 135776 213242 135788
rect 234246 135776 234252 135788
rect 213236 135748 234252 135776
rect 213236 135736 213242 135748
rect 234246 135736 234252 135748
rect 234304 135736 234310 135788
rect 246298 135736 246304 135788
rect 246356 135776 246362 135788
rect 254026 135776 254032 135788
rect 246356 135748 254032 135776
rect 246356 135736 246362 135748
rect 254026 135736 254032 135748
rect 254084 135736 254090 135788
rect 329926 135736 329932 135788
rect 329984 135776 329990 135788
rect 335998 135776 336004 135788
rect 329984 135748 336004 135776
rect 329984 135736 329990 135748
rect 335998 135736 336004 135748
rect 336056 135736 336062 135788
rect 432414 135736 432420 135788
rect 432472 135776 432478 135788
rect 480349 135779 480407 135785
rect 480349 135776 480361 135779
rect 432472 135748 480361 135776
rect 432472 135736 432478 135748
rect 480349 135745 480361 135748
rect 480395 135745 480407 135779
rect 480349 135739 480407 135745
rect 86862 135668 86868 135720
rect 86920 135708 86926 135720
rect 142062 135708 142068 135720
rect 86920 135680 142068 135708
rect 86920 135668 86926 135680
rect 142062 135668 142068 135680
rect 142120 135668 142126 135720
rect 180058 135668 180064 135720
rect 180116 135708 180122 135720
rect 185210 135708 185216 135720
rect 180116 135680 185216 135708
rect 180116 135668 180122 135680
rect 185210 135668 185216 135680
rect 185268 135668 185274 135720
rect 199378 135668 199384 135720
rect 199436 135708 199442 135720
rect 219989 135711 220047 135717
rect 219989 135708 220001 135711
rect 199436 135680 220001 135708
rect 199436 135668 199442 135680
rect 219989 135677 220001 135680
rect 220035 135677 220047 135711
rect 219989 135671 220047 135677
rect 220078 135668 220084 135720
rect 220136 135708 220142 135720
rect 224770 135708 224776 135720
rect 220136 135680 224776 135708
rect 220136 135668 220142 135680
rect 224770 135668 224776 135680
rect 224828 135668 224834 135720
rect 226242 135668 226248 135720
rect 226300 135708 226306 135720
rect 243722 135708 243728 135720
rect 226300 135680 243728 135708
rect 226300 135668 226306 135680
rect 243722 135668 243728 135680
rect 243780 135668 243786 135720
rect 251818 135668 251824 135720
rect 251876 135708 251882 135720
rect 260098 135708 260104 135720
rect 251876 135680 260104 135708
rect 251876 135668 251882 135680
rect 260098 135668 260104 135680
rect 260156 135668 260162 135720
rect 304902 135668 304908 135720
rect 304960 135708 304966 135720
rect 305638 135708 305644 135720
rect 304960 135680 305644 135708
rect 304960 135668 304966 135680
rect 305638 135668 305644 135680
rect 305696 135668 305702 135720
rect 427262 135668 427268 135720
rect 427320 135708 427326 135720
rect 436646 135708 436652 135720
rect 427320 135680 436652 135708
rect 427320 135668 427326 135680
rect 436646 135668 436652 135680
rect 436704 135668 436710 135720
rect 438486 135668 438492 135720
rect 438544 135708 438550 135720
rect 480548 135708 480576 135816
rect 486418 135804 486424 135816
rect 486476 135804 486482 135856
rect 520918 135844 520924 135856
rect 489886 135816 520924 135844
rect 486694 135736 486700 135788
rect 486752 135776 486758 135788
rect 489886 135776 489914 135816
rect 520918 135804 520924 135816
rect 520976 135804 520982 135856
rect 486752 135748 489914 135776
rect 486752 135736 486758 135748
rect 499482 135736 499488 135788
rect 499540 135776 499546 135788
rect 526438 135776 526444 135788
rect 499540 135748 526444 135776
rect 499540 135736 499546 135748
rect 526438 135736 526444 135748
rect 526496 135736 526502 135788
rect 438544 135680 480576 135708
rect 438544 135668 438550 135680
rect 480622 135668 480628 135720
rect 480680 135708 480686 135720
rect 481542 135708 481548 135720
rect 480680 135680 481548 135708
rect 480680 135668 480686 135680
rect 481542 135668 481548 135680
rect 481600 135668 481606 135720
rect 483198 135668 483204 135720
rect 483256 135708 483262 135720
rect 484210 135708 484216 135720
rect 483256 135680 484216 135708
rect 483256 135668 483262 135680
rect 484210 135668 484216 135680
rect 484268 135668 484274 135720
rect 485866 135668 485872 135720
rect 485924 135708 485930 135720
rect 487062 135708 487068 135720
rect 485924 135680 487068 135708
rect 485924 135668 485930 135680
rect 487062 135668 487068 135680
rect 487120 135668 487126 135720
rect 489270 135668 489276 135720
rect 489328 135708 489334 135720
rect 489822 135708 489828 135720
rect 489328 135680 489828 135708
rect 489328 135668 489334 135680
rect 489822 135668 489828 135680
rect 489880 135668 489886 135720
rect 490098 135668 490104 135720
rect 490156 135708 490162 135720
rect 491202 135708 491208 135720
rect 490156 135680 491208 135708
rect 490156 135668 490162 135680
rect 491202 135668 491208 135680
rect 491260 135668 491266 135720
rect 491846 135668 491852 135720
rect 491904 135708 491910 135720
rect 493870 135708 493876 135720
rect 491904 135680 493876 135708
rect 491904 135668 491910 135680
rect 493870 135668 493876 135680
rect 493928 135668 493934 135720
rect 494422 135668 494428 135720
rect 494480 135708 494486 135720
rect 522298 135708 522304 135720
rect 494480 135680 522304 135708
rect 494480 135668 494486 135680
rect 522298 135668 522304 135680
rect 522356 135668 522362 135720
rect 47578 135600 47584 135652
rect 47636 135640 47642 135652
rect 101674 135640 101680 135652
rect 47636 135612 101680 135640
rect 47636 135600 47642 135612
rect 101674 135600 101680 135612
rect 101732 135600 101738 135652
rect 130378 135600 130384 135652
rect 130436 135640 130442 135652
rect 153286 135640 153292 135652
rect 130436 135612 153292 135640
rect 130436 135600 130442 135612
rect 153286 135600 153292 135612
rect 153344 135600 153350 135652
rect 197998 135600 198004 135652
rect 198056 135640 198062 135652
rect 199838 135640 199844 135652
rect 198056 135612 199844 135640
rect 198056 135600 198062 135612
rect 199838 135600 199844 135612
rect 199896 135600 199902 135652
rect 199933 135643 199991 135649
rect 199933 135609 199945 135643
rect 199979 135640 199991 135643
rect 200669 135643 200727 135649
rect 200669 135640 200681 135643
rect 199979 135612 200681 135640
rect 199979 135609 199991 135612
rect 199933 135603 199991 135609
rect 200669 135609 200681 135612
rect 200715 135609 200727 135643
rect 200669 135603 200727 135609
rect 200758 135600 200764 135652
rect 200816 135640 200822 135652
rect 202414 135640 202420 135652
rect 200816 135612 202420 135640
rect 200816 135600 200822 135612
rect 202414 135600 202420 135612
rect 202472 135600 202478 135652
rect 206922 135600 206928 135652
rect 206980 135640 206986 135652
rect 229922 135640 229928 135652
rect 206980 135612 229928 135640
rect 206980 135600 206986 135612
rect 229922 135600 229928 135612
rect 229980 135600 229986 135652
rect 233142 135600 233148 135652
rect 233200 135640 233206 135652
rect 248874 135640 248880 135652
rect 233200 135612 248880 135640
rect 233200 135600 233206 135612
rect 248874 135600 248880 135612
rect 248932 135600 248938 135652
rect 268930 135600 268936 135652
rect 268988 135640 268994 135652
rect 274726 135640 274732 135652
rect 268988 135612 274732 135640
rect 268988 135600 268994 135612
rect 274726 135600 274732 135612
rect 274784 135600 274790 135652
rect 280798 135600 280804 135652
rect 280856 135640 280862 135652
rect 283374 135640 283380 135652
rect 280856 135612 283380 135640
rect 280856 135600 280862 135612
rect 283374 135600 283380 135612
rect 283432 135600 283438 135652
rect 289814 135600 289820 135652
rect 289872 135640 289878 135652
rect 291102 135640 291108 135652
rect 289872 135612 291108 135640
rect 289872 135600 289878 135612
rect 291102 135600 291108 135612
rect 291160 135600 291166 135652
rect 297174 135600 297180 135652
rect 297232 135640 297238 135652
rect 298094 135640 298100 135652
rect 297232 135612 298100 135640
rect 297232 135600 297238 135612
rect 298094 135600 298100 135612
rect 298152 135600 298158 135652
rect 300670 135600 300676 135652
rect 300728 135640 300734 135652
rect 302234 135640 302240 135652
rect 300728 135612 302240 135640
rect 300728 135600 300734 135612
rect 302234 135600 302240 135612
rect 302292 135600 302298 135652
rect 302418 135600 302424 135652
rect 302476 135640 302482 135652
rect 304994 135640 305000 135652
rect 302476 135612 305000 135640
rect 302476 135600 302482 135612
rect 304994 135600 305000 135612
rect 305052 135600 305058 135652
rect 320450 135600 320456 135652
rect 320508 135640 320514 135652
rect 321462 135640 321468 135652
rect 320508 135612 321468 135640
rect 320508 135600 320514 135612
rect 321462 135600 321468 135612
rect 321520 135600 321526 135652
rect 327350 135600 327356 135652
rect 327408 135640 327414 135652
rect 328362 135640 328368 135652
rect 327408 135612 328368 135640
rect 327408 135600 327414 135612
rect 328362 135600 328368 135612
rect 328420 135600 328426 135652
rect 338574 135600 338580 135652
rect 338632 135640 338638 135652
rect 339402 135640 339408 135652
rect 338632 135612 339408 135640
rect 338632 135600 338638 135612
rect 339402 135600 339408 135612
rect 339460 135600 339466 135652
rect 354950 135600 354956 135652
rect 355008 135640 355014 135652
rect 356698 135640 356704 135652
rect 355008 135612 356704 135640
rect 355008 135600 355014 135612
rect 356698 135600 356704 135612
rect 356756 135600 356762 135652
rect 362678 135600 362684 135652
rect 362736 135640 362742 135652
rect 363598 135640 363604 135652
rect 362736 135612 363604 135640
rect 362736 135600 362742 135612
rect 363598 135600 363604 135612
rect 363656 135600 363662 135652
rect 429838 135600 429844 135652
rect 429896 135640 429902 135652
rect 429896 135612 453068 135640
rect 429896 135600 429902 135612
rect 72418 135532 72424 135584
rect 72476 135572 72482 135584
rect 123202 135572 123208 135584
rect 72476 135544 123208 135572
rect 72476 135532 72482 135544
rect 123202 135532 123208 135544
rect 123260 135532 123266 135584
rect 137278 135532 137284 135584
rect 137336 135572 137342 135584
rect 140406 135572 140412 135584
rect 137336 135544 140412 135572
rect 137336 135532 137342 135544
rect 140406 135532 140412 135544
rect 140464 135532 140470 135584
rect 163682 135572 163688 135584
rect 142126 135544 163688 135572
rect 75178 135464 75184 135516
rect 75236 135504 75242 135516
rect 82722 135504 82728 135516
rect 75236 135476 82728 135504
rect 75236 135464 75242 135476
rect 82722 135464 82728 135476
rect 82780 135464 82786 135516
rect 83458 135464 83464 135516
rect 83516 135504 83522 135516
rect 130010 135504 130016 135516
rect 83516 135476 130016 135504
rect 83516 135464 83522 135476
rect 130010 135464 130016 135476
rect 130068 135464 130074 135516
rect 133138 135464 133144 135516
rect 133196 135504 133202 135516
rect 142126 135504 142154 135544
rect 163682 135532 163688 135544
rect 163740 135532 163746 135584
rect 188338 135532 188344 135584
rect 188396 135572 188402 135584
rect 189442 135572 189448 135584
rect 188396 135544 189448 135572
rect 188396 135532 188402 135544
rect 189442 135532 189448 135544
rect 189500 135532 189506 135584
rect 213546 135572 213552 135584
rect 190426 135544 213552 135572
rect 133196 135476 142154 135504
rect 133196 135464 133202 135476
rect 184842 135464 184848 135516
rect 184900 135504 184906 135516
rect 190426 135504 190454 135544
rect 213546 135532 213552 135544
rect 213604 135532 213610 135584
rect 217962 135532 217968 135584
rect 218020 135572 218026 135584
rect 237742 135572 237748 135584
rect 218020 135544 237748 135572
rect 218020 135532 218026 135544
rect 237742 135532 237748 135544
rect 237800 135532 237806 135584
rect 249058 135532 249064 135584
rect 249116 135572 249122 135584
rect 256694 135572 256700 135584
rect 249116 135544 256700 135572
rect 249116 135532 249122 135544
rect 256694 135532 256700 135544
rect 256752 135532 256758 135584
rect 269758 135532 269764 135584
rect 269816 135572 269822 135584
rect 272978 135572 272984 135584
rect 269816 135544 272984 135572
rect 269816 135532 269822 135544
rect 272978 135532 272984 135544
rect 273036 135532 273042 135584
rect 282178 135532 282184 135584
rect 282236 135572 282242 135584
rect 284202 135572 284208 135584
rect 282236 135544 284208 135572
rect 282236 135532 282242 135544
rect 284202 135532 284208 135544
rect 284260 135532 284266 135584
rect 284938 135532 284944 135584
rect 284996 135572 285002 135584
rect 285950 135572 285956 135584
rect 284996 135544 285956 135572
rect 284996 135532 285002 135544
rect 285950 135532 285956 135544
rect 286008 135532 286014 135584
rect 288342 135532 288348 135584
rect 288400 135572 288406 135584
rect 289354 135572 289360 135584
rect 288400 135544 289360 135572
rect 288400 135532 288406 135544
rect 289354 135532 289360 135544
rect 289412 135532 289418 135584
rect 289722 135532 289728 135584
rect 289780 135572 289786 135584
rect 290274 135572 290280 135584
rect 289780 135544 290280 135572
rect 289780 135532 289786 135544
rect 290274 135532 290280 135544
rect 290332 135532 290338 135584
rect 292574 135532 292580 135584
rect 292632 135572 292638 135584
rect 293678 135572 293684 135584
rect 292632 135544 293684 135572
rect 292632 135532 292638 135544
rect 293678 135532 293684 135544
rect 293736 135532 293742 135584
rect 298002 135532 298008 135584
rect 298060 135572 298066 135584
rect 298738 135572 298744 135584
rect 298060 135544 298744 135572
rect 298060 135532 298066 135544
rect 298738 135532 298744 135544
rect 298796 135532 298802 135584
rect 298922 135532 298928 135584
rect 298980 135572 298986 135584
rect 299566 135572 299572 135584
rect 298980 135544 299572 135572
rect 298980 135532 298986 135544
rect 299566 135532 299572 135544
rect 299624 135532 299630 135584
rect 299842 135532 299848 135584
rect 299900 135572 299906 135584
rect 300762 135572 300768 135584
rect 299900 135544 300768 135572
rect 299900 135532 299906 135544
rect 300762 135532 300768 135544
rect 300820 135532 300826 135584
rect 301498 135532 301504 135584
rect 301556 135572 301562 135584
rect 303614 135572 303620 135584
rect 301556 135544 303620 135572
rect 301556 135532 301562 135544
rect 303614 135532 303620 135544
rect 303672 135532 303678 135584
rect 304074 135532 304080 135584
rect 304132 135572 304138 135584
rect 304902 135572 304908 135584
rect 304132 135544 304908 135572
rect 304132 135532 304138 135544
rect 304902 135532 304908 135544
rect 304960 135532 304966 135584
rect 306650 135532 306656 135584
rect 306708 135572 306714 135584
rect 307662 135572 307668 135584
rect 306708 135544 307668 135572
rect 306708 135532 306714 135544
rect 307662 135532 307668 135544
rect 307720 135532 307726 135584
rect 309318 135532 309324 135584
rect 309376 135572 309382 135584
rect 310330 135572 310336 135584
rect 309376 135544 310336 135572
rect 309376 135532 309382 135544
rect 310330 135532 310336 135544
rect 310388 135532 310394 135584
rect 310974 135532 310980 135584
rect 311032 135572 311038 135584
rect 311710 135572 311716 135584
rect 311032 135544 311716 135572
rect 311032 135532 311038 135544
rect 311710 135532 311716 135544
rect 311768 135532 311774 135584
rect 312722 135532 312728 135584
rect 312780 135572 312786 135584
rect 313182 135572 313188 135584
rect 312780 135544 313188 135572
rect 312780 135532 312786 135544
rect 313182 135532 313188 135544
rect 313240 135532 313246 135584
rect 313550 135532 313556 135584
rect 313608 135572 313614 135584
rect 314562 135572 314568 135584
rect 313608 135544 314568 135572
rect 313608 135532 313614 135544
rect 314562 135532 314568 135544
rect 314620 135532 314626 135584
rect 316126 135532 316132 135584
rect 316184 135572 316190 135584
rect 317322 135572 317328 135584
rect 316184 135544 317328 135572
rect 316184 135532 316190 135544
rect 317322 135532 317328 135544
rect 317380 135532 317386 135584
rect 317874 135532 317880 135584
rect 317932 135572 317938 135584
rect 318702 135572 318708 135584
rect 317932 135544 318708 135572
rect 317932 135532 317938 135544
rect 318702 135532 318708 135544
rect 318760 135532 318766 135584
rect 319622 135532 319628 135584
rect 319680 135572 319686 135584
rect 320818 135572 320824 135584
rect 319680 135544 320824 135572
rect 319680 135532 319686 135544
rect 320818 135532 320824 135544
rect 320876 135532 320882 135584
rect 322198 135532 322204 135584
rect 322256 135572 322262 135584
rect 322842 135572 322848 135584
rect 322256 135544 322848 135572
rect 322256 135532 322262 135544
rect 322842 135532 322848 135544
rect 322900 135532 322906 135584
rect 323026 135532 323032 135584
rect 323084 135572 323090 135584
rect 324222 135572 324228 135584
rect 323084 135544 324228 135572
rect 323084 135532 323090 135544
rect 324222 135532 324228 135544
rect 324280 135532 324286 135584
rect 324774 135532 324780 135584
rect 324832 135572 324838 135584
rect 325602 135572 325608 135584
rect 324832 135544 325608 135572
rect 324832 135532 324838 135544
rect 325602 135532 325608 135544
rect 325660 135532 325666 135584
rect 326522 135532 326528 135584
rect 326580 135572 326586 135584
rect 327718 135572 327724 135584
rect 326580 135544 327724 135572
rect 326580 135532 326586 135544
rect 327718 135532 327724 135544
rect 327776 135532 327782 135584
rect 329098 135532 329104 135584
rect 329156 135572 329162 135584
rect 329742 135572 329748 135584
rect 329156 135544 329748 135572
rect 329156 135532 329162 135544
rect 329742 135532 329748 135544
rect 329800 135532 329806 135584
rect 331674 135532 331680 135584
rect 331732 135572 331738 135584
rect 332410 135572 332416 135584
rect 331732 135544 332416 135572
rect 331732 135532 331738 135544
rect 332410 135532 332416 135544
rect 332468 135532 332474 135584
rect 334250 135532 334256 135584
rect 334308 135572 334314 135584
rect 335170 135572 335176 135584
rect 334308 135544 335176 135572
rect 334308 135532 334314 135544
rect 335170 135532 335176 135544
rect 335228 135532 335234 135584
rect 336826 135532 336832 135584
rect 336884 135572 336890 135584
rect 338758 135572 338764 135584
rect 336884 135544 338764 135572
rect 336884 135532 336890 135544
rect 338758 135532 338764 135544
rect 338816 135532 338822 135584
rect 340322 135532 340328 135584
rect 340380 135572 340386 135584
rect 340782 135572 340788 135584
rect 340380 135544 340788 135572
rect 340380 135532 340386 135544
rect 340782 135532 340788 135544
rect 340840 135532 340846 135584
rect 341150 135532 341156 135584
rect 341208 135572 341214 135584
rect 342162 135572 342168 135584
rect 341208 135544 342168 135572
rect 341208 135532 341214 135544
rect 342162 135532 342168 135544
rect 342220 135532 342226 135584
rect 342898 135532 342904 135584
rect 342956 135572 342962 135584
rect 343542 135572 343548 135584
rect 342956 135544 343548 135572
rect 342956 135532 342962 135544
rect 343542 135532 343548 135544
rect 343600 135532 343606 135584
rect 343726 135532 343732 135584
rect 343784 135572 343790 135584
rect 344922 135572 344928 135584
rect 343784 135544 344928 135572
rect 343784 135532 343790 135544
rect 344922 135532 344928 135544
rect 344980 135532 344986 135584
rect 345474 135532 345480 135584
rect 345532 135572 345538 135584
rect 346302 135572 346308 135584
rect 345532 135544 346308 135572
rect 345532 135532 345538 135544
rect 346302 135532 346308 135544
rect 346360 135532 346366 135584
rect 347130 135532 347136 135584
rect 347188 135572 347194 135584
rect 347682 135572 347688 135584
rect 347188 135544 347688 135572
rect 347188 135532 347194 135544
rect 347682 135532 347688 135544
rect 347740 135532 347746 135584
rect 348050 135532 348056 135584
rect 348108 135572 348114 135584
rect 349062 135572 349068 135584
rect 348108 135544 349068 135572
rect 348108 135532 348114 135544
rect 349062 135532 349068 135544
rect 349120 135532 349126 135584
rect 349798 135532 349804 135584
rect 349856 135572 349862 135584
rect 350442 135572 350448 135584
rect 349856 135544 350448 135572
rect 349856 135532 349862 135544
rect 350442 135532 350448 135544
rect 350500 135532 350506 135584
rect 350626 135532 350632 135584
rect 350684 135572 350690 135584
rect 351730 135572 351736 135584
rect 350684 135544 351736 135572
rect 350684 135532 350690 135544
rect 351730 135532 351736 135544
rect 351788 135532 351794 135584
rect 354030 135532 354036 135584
rect 354088 135572 354094 135584
rect 354582 135572 354588 135584
rect 354088 135544 354588 135572
rect 354088 135532 354094 135544
rect 354582 135532 354588 135544
rect 354640 135532 354646 135584
rect 356606 135532 356612 135584
rect 356664 135572 356670 135584
rect 357342 135572 357348 135584
rect 356664 135544 357348 135572
rect 356664 135532 356670 135544
rect 357342 135532 357348 135544
rect 357400 135532 357406 135584
rect 357526 135532 357532 135584
rect 357584 135572 357590 135584
rect 358630 135572 358636 135584
rect 357584 135544 358636 135572
rect 357584 135532 357590 135544
rect 358630 135532 358636 135544
rect 358688 135532 358694 135584
rect 359182 135532 359188 135584
rect 359240 135572 359246 135584
rect 360102 135572 360108 135584
rect 359240 135544 360108 135572
rect 359240 135532 359246 135544
rect 360102 135532 360108 135544
rect 360160 135532 360166 135584
rect 360930 135532 360936 135584
rect 360988 135572 360994 135584
rect 361482 135572 361488 135584
rect 360988 135544 361488 135572
rect 360988 135532 360994 135544
rect 361482 135532 361488 135544
rect 361540 135532 361546 135584
rect 361850 135532 361856 135584
rect 361908 135572 361914 135584
rect 362862 135572 362868 135584
rect 361908 135544 362868 135572
rect 361908 135532 361914 135544
rect 362862 135532 362868 135544
rect 362920 135532 362926 135584
rect 363506 135532 363512 135584
rect 363564 135572 363570 135584
rect 364242 135572 364248 135584
rect 363564 135544 364248 135572
rect 363564 135532 363570 135544
rect 364242 135532 364248 135544
rect 364300 135532 364306 135584
rect 364426 135532 364432 135584
rect 364484 135572 364490 135584
rect 365622 135572 365628 135584
rect 364484 135544 365628 135572
rect 364484 135532 364490 135544
rect 365622 135532 365628 135544
rect 365680 135532 365686 135584
rect 366082 135532 366088 135584
rect 366140 135572 366146 135584
rect 367002 135572 367008 135584
rect 366140 135544 367008 135572
rect 366140 135532 366146 135544
rect 367002 135532 367008 135544
rect 367060 135532 367066 135584
rect 367830 135532 367836 135584
rect 367888 135572 367894 135584
rect 368382 135572 368388 135584
rect 367888 135544 368388 135572
rect 367888 135532 367894 135544
rect 368382 135532 368388 135544
rect 368440 135532 368446 135584
rect 368658 135532 368664 135584
rect 368716 135572 368722 135584
rect 369762 135572 369768 135584
rect 368716 135544 369768 135572
rect 368716 135532 368722 135544
rect 369762 135532 369768 135544
rect 369820 135532 369826 135584
rect 370406 135532 370412 135584
rect 370464 135572 370470 135584
rect 371142 135572 371148 135584
rect 370464 135544 371148 135572
rect 370464 135532 370470 135544
rect 371142 135532 371148 135544
rect 371200 135532 371206 135584
rect 371326 135532 371332 135584
rect 371384 135572 371390 135584
rect 372430 135572 372436 135584
rect 371384 135544 372436 135572
rect 371384 135532 371390 135544
rect 372430 135532 372436 135544
rect 372488 135532 372494 135584
rect 374730 135532 374736 135584
rect 374788 135572 374794 135584
rect 375282 135572 375288 135584
rect 374788 135544 375288 135572
rect 374788 135532 374794 135544
rect 375282 135532 375288 135544
rect 375340 135532 375346 135584
rect 375558 135532 375564 135584
rect 375616 135572 375622 135584
rect 376570 135572 376576 135584
rect 375616 135544 376576 135572
rect 375616 135532 375622 135544
rect 376570 135532 376576 135544
rect 376628 135532 376634 135584
rect 381630 135532 381636 135584
rect 381688 135572 381694 135584
rect 382182 135572 382188 135584
rect 381688 135544 382188 135572
rect 381688 135532 381694 135544
rect 382182 135532 382188 135544
rect 382240 135532 382246 135584
rect 382458 135532 382464 135584
rect 382516 135572 382522 135584
rect 383562 135572 383568 135584
rect 382516 135544 383568 135572
rect 382516 135532 382522 135544
rect 383562 135532 383568 135544
rect 383620 135532 383626 135584
rect 384206 135532 384212 135584
rect 384264 135572 384270 135584
rect 384942 135572 384948 135584
rect 384264 135544 384948 135572
rect 384264 135532 384270 135544
rect 384942 135532 384948 135544
rect 385000 135532 385006 135584
rect 386782 135532 386788 135584
rect 386840 135572 386846 135584
rect 387610 135572 387616 135584
rect 386840 135544 387616 135572
rect 386840 135532 386846 135544
rect 387610 135532 387616 135544
rect 387668 135532 387674 135584
rect 388530 135532 388536 135584
rect 388588 135572 388594 135584
rect 389082 135572 389088 135584
rect 388588 135544 389088 135572
rect 388588 135532 388594 135544
rect 389082 135532 389088 135544
rect 389140 135532 389146 135584
rect 389358 135532 389364 135584
rect 389416 135572 389422 135584
rect 390462 135572 390468 135584
rect 389416 135544 390468 135572
rect 389416 135532 389422 135544
rect 390462 135532 390468 135544
rect 390520 135532 390526 135584
rect 396258 135532 396264 135584
rect 396316 135572 396322 135584
rect 397362 135572 397368 135584
rect 396316 135544 397368 135572
rect 396316 135532 396322 135544
rect 397362 135532 397368 135544
rect 397420 135532 397426 135584
rect 398006 135532 398012 135584
rect 398064 135572 398070 135584
rect 398742 135572 398748 135584
rect 398064 135544 398748 135572
rect 398064 135532 398070 135544
rect 398742 135532 398748 135544
rect 398800 135532 398806 135584
rect 403158 135532 403164 135584
rect 403216 135572 403222 135584
rect 404262 135572 404268 135584
rect 403216 135544 404268 135572
rect 403216 135532 403222 135544
rect 404262 135532 404268 135544
rect 404320 135532 404326 135584
rect 404906 135532 404912 135584
rect 404964 135572 404970 135584
rect 406378 135572 406384 135584
rect 404964 135544 406384 135572
rect 404964 135532 404970 135544
rect 406378 135532 406384 135544
rect 406436 135532 406442 135584
rect 406562 135532 406568 135584
rect 406620 135572 406626 135584
rect 407022 135572 407028 135584
rect 406620 135544 407028 135572
rect 406620 135532 406626 135544
rect 407022 135532 407028 135544
rect 407080 135532 407086 135584
rect 418614 135532 418620 135584
rect 418672 135572 418678 135584
rect 419442 135572 419448 135584
rect 418672 135544 419448 135572
rect 418672 135532 418678 135544
rect 419442 135532 419448 135544
rect 419500 135532 419506 135584
rect 420362 135532 420368 135584
rect 420420 135572 420426 135584
rect 420822 135572 420828 135584
rect 420420 135544 420828 135572
rect 420420 135532 420426 135544
rect 420822 135532 420828 135544
rect 420880 135532 420886 135584
rect 421190 135532 421196 135584
rect 421248 135572 421254 135584
rect 422202 135572 422208 135584
rect 421248 135544 422208 135572
rect 421248 135532 421254 135544
rect 422202 135532 422208 135544
rect 422260 135532 422266 135584
rect 422938 135532 422944 135584
rect 422996 135572 423002 135584
rect 423582 135572 423588 135584
rect 422996 135544 423588 135572
rect 422996 135532 423002 135544
rect 423582 135532 423588 135544
rect 423640 135532 423646 135584
rect 423858 135532 423864 135584
rect 423916 135572 423922 135584
rect 424962 135572 424968 135584
rect 423916 135544 424968 135572
rect 423916 135532 423922 135544
rect 424962 135532 424968 135544
rect 425020 135532 425026 135584
rect 428090 135532 428096 135584
rect 428148 135572 428154 135584
rect 429102 135572 429108 135584
rect 428148 135544 429108 135572
rect 428148 135532 428154 135544
rect 429102 135532 429108 135544
rect 429160 135532 429166 135584
rect 430666 135532 430672 135584
rect 430724 135572 430730 135584
rect 431770 135572 431776 135584
rect 430724 135544 431776 135572
rect 430724 135532 430730 135544
rect 431770 135532 431776 135544
rect 431828 135532 431834 135584
rect 434162 135532 434168 135584
rect 434220 135572 434226 135584
rect 434622 135572 434628 135584
rect 434220 135544 434628 135572
rect 434220 135532 434226 135544
rect 434622 135532 434628 135544
rect 434680 135532 434686 135584
rect 436738 135532 436744 135584
rect 436796 135572 436802 135584
rect 437382 135572 437388 135584
rect 436796 135544 437388 135572
rect 436796 135532 436802 135544
rect 437382 135532 437388 135544
rect 437440 135532 437446 135584
rect 437566 135532 437572 135584
rect 437624 135572 437630 135584
rect 438762 135572 438768 135584
rect 437624 135544 438768 135572
rect 437624 135532 437630 135544
rect 438762 135532 438768 135544
rect 438820 135532 438826 135584
rect 439314 135532 439320 135584
rect 439372 135572 439378 135584
rect 440142 135572 440148 135584
rect 439372 135544 440148 135572
rect 439372 135532 439378 135544
rect 440142 135532 440148 135544
rect 440200 135532 440206 135584
rect 441890 135532 441896 135584
rect 441948 135572 441954 135584
rect 442902 135572 442908 135584
rect 441948 135544 442908 135572
rect 441948 135532 441954 135544
rect 442902 135532 442908 135544
rect 442960 135532 442966 135584
rect 446214 135532 446220 135584
rect 446272 135572 446278 135584
rect 446950 135572 446956 135584
rect 446272 135544 446956 135572
rect 446272 135532 446278 135544
rect 446950 135532 446956 135544
rect 447008 135532 447014 135584
rect 447962 135532 447968 135584
rect 448020 135572 448026 135584
rect 448422 135572 448428 135584
rect 448020 135544 448428 135572
rect 448020 135532 448026 135544
rect 448422 135532 448428 135544
rect 448480 135532 448486 135584
rect 448790 135532 448796 135584
rect 448848 135572 448854 135584
rect 449802 135572 449808 135584
rect 448848 135544 449808 135572
rect 448848 135532 448854 135544
rect 449802 135532 449808 135544
rect 449860 135532 449866 135584
rect 449912 135544 452976 135572
rect 184900 135476 190454 135504
rect 184900 135464 184906 135476
rect 191098 135464 191104 135516
rect 191156 135504 191162 135516
rect 199933 135507 199991 135513
rect 199933 135504 199945 135507
rect 191156 135476 199945 135504
rect 191156 135464 191162 135476
rect 199933 135473 199945 135476
rect 199979 135473 199991 135507
rect 199933 135467 199991 135473
rect 220722 135464 220728 135516
rect 220780 135504 220786 135516
rect 222289 135507 222347 135513
rect 222289 135504 222301 135507
rect 220780 135476 222301 135504
rect 220780 135464 220786 135476
rect 222289 135473 222301 135476
rect 222335 135473 222347 135507
rect 222289 135467 222347 135473
rect 224218 135464 224224 135516
rect 224276 135504 224282 135516
rect 232498 135504 232504 135516
rect 224276 135476 232504 135504
rect 224276 135464 224282 135476
rect 232498 135464 232504 135476
rect 232556 135464 232562 135516
rect 233878 135464 233884 135516
rect 233936 135504 233942 135516
rect 247218 135504 247224 135516
rect 233936 135476 247224 135504
rect 233936 135464 233942 135476
rect 247218 135464 247224 135476
rect 247276 135464 247282 135516
rect 251910 135464 251916 135516
rect 251968 135504 251974 135516
rect 257522 135504 257528 135516
rect 251968 135476 257528 135504
rect 251968 135464 251974 135476
rect 257522 135464 257528 135476
rect 257580 135464 257586 135516
rect 269022 135464 269028 135516
rect 269080 135504 269086 135516
rect 275554 135504 275560 135516
rect 269080 135476 275560 135504
rect 269080 135464 269086 135476
rect 275554 135464 275560 135476
rect 275612 135464 275618 135516
rect 278682 135464 278688 135516
rect 278740 135504 278746 135516
rect 282454 135504 282460 135516
rect 278740 135476 282460 135504
rect 278740 135464 278746 135476
rect 282454 135464 282460 135476
rect 282512 135464 282518 135516
rect 308398 135464 308404 135516
rect 308456 135504 308462 135516
rect 313366 135504 313372 135516
rect 308456 135476 313372 135504
rect 308456 135464 308462 135476
rect 313366 135464 313372 135476
rect 313424 135464 313430 135516
rect 317046 135464 317052 135516
rect 317104 135504 317110 135516
rect 324498 135504 324504 135516
rect 317104 135476 324504 135504
rect 317104 135464 317110 135476
rect 324498 135464 324504 135476
rect 324556 135464 324562 135516
rect 337654 135464 337660 135516
rect 337712 135504 337718 135516
rect 340138 135504 340144 135516
rect 337712 135476 340144 135504
rect 337712 135464 337718 135476
rect 340138 135464 340144 135476
rect 340196 135464 340202 135516
rect 377306 135464 377312 135516
rect 377364 135504 377370 135516
rect 378042 135504 378048 135516
rect 377364 135476 378048 135504
rect 377364 135464 377370 135476
rect 378042 135464 378048 135476
rect 378100 135464 378106 135516
rect 380802 135464 380808 135516
rect 380860 135504 380866 135516
rect 381538 135504 381544 135516
rect 380860 135476 381544 135504
rect 380860 135464 380866 135476
rect 381538 135464 381544 135476
rect 381596 135464 381602 135516
rect 425514 135464 425520 135516
rect 425572 135504 425578 135516
rect 426342 135504 426348 135516
rect 425572 135476 426348 135504
rect 425572 135464 425578 135476
rect 426342 135464 426348 135476
rect 426400 135464 426406 135516
rect 443546 135464 443552 135516
rect 443604 135504 443610 135516
rect 449912 135504 449940 135544
rect 443604 135476 449940 135504
rect 443604 135464 443610 135476
rect 450538 135464 450544 135516
rect 450596 135504 450602 135516
rect 451182 135504 451188 135516
rect 450596 135476 451188 135504
rect 450596 135464 450602 135476
rect 451182 135464 451188 135476
rect 451240 135464 451246 135516
rect 76926 135396 76932 135448
rect 76984 135436 76990 135448
rect 95602 135436 95608 135448
rect 76984 135408 95608 135436
rect 76984 135396 76990 135408
rect 95602 135396 95608 135408
rect 95660 135396 95666 135448
rect 219342 135396 219348 135448
rect 219400 135436 219406 135448
rect 238570 135436 238576 135448
rect 219400 135408 238576 135436
rect 219400 135396 219406 135408
rect 238570 135396 238576 135408
rect 238628 135396 238634 135448
rect 270402 135396 270408 135448
rect 270460 135436 270466 135448
rect 276474 135436 276480 135448
rect 270460 135408 276480 135436
rect 270460 135396 270466 135408
rect 276474 135396 276480 135408
rect 276532 135396 276538 135448
rect 452948 135436 452976 135544
rect 453040 135504 453068 135612
rect 453114 135600 453120 135652
rect 453172 135640 453178 135652
rect 453942 135640 453948 135652
rect 453172 135612 453948 135640
rect 453172 135600 453178 135612
rect 453942 135600 453948 135612
rect 454000 135600 454006 135652
rect 454862 135600 454868 135652
rect 454920 135640 454926 135652
rect 455322 135640 455328 135652
rect 454920 135612 455328 135640
rect 454920 135600 454926 135612
rect 455322 135600 455328 135612
rect 455380 135600 455386 135652
rect 455690 135600 455696 135652
rect 455748 135640 455754 135652
rect 456702 135640 456708 135652
rect 455748 135612 456708 135640
rect 455748 135600 455754 135612
rect 456702 135600 456708 135612
rect 456760 135600 456766 135652
rect 466914 135600 466920 135652
rect 466972 135640 466978 135652
rect 467742 135640 467748 135652
rect 466972 135612 467748 135640
rect 466972 135600 466978 135612
rect 467742 135600 467748 135612
rect 467800 135600 467806 135652
rect 468570 135600 468576 135652
rect 468628 135640 468634 135652
rect 469122 135640 469128 135652
rect 468628 135612 469128 135640
rect 468628 135600 468634 135612
rect 469122 135600 469128 135612
rect 469180 135600 469186 135652
rect 512638 135640 512644 135652
rect 469324 135612 512644 135640
rect 457438 135504 457444 135516
rect 453040 135476 457444 135504
rect 457438 135464 457444 135476
rect 457496 135464 457502 135516
rect 465994 135464 466000 135516
rect 466052 135504 466058 135516
rect 469324 135504 469352 135612
rect 512638 135600 512644 135612
rect 512696 135600 512702 135652
rect 471146 135532 471152 135584
rect 471204 135572 471210 135584
rect 471882 135572 471888 135584
rect 471204 135544 471888 135572
rect 471204 135532 471210 135544
rect 471882 135532 471888 135544
rect 471940 135532 471946 135584
rect 472066 135532 472072 135584
rect 472124 135572 472130 135584
rect 473262 135572 473268 135584
rect 472124 135544 473268 135572
rect 472124 135532 472130 135544
rect 473262 135532 473268 135544
rect 473320 135532 473326 135584
rect 475470 135532 475476 135584
rect 475528 135572 475534 135584
rect 476022 135572 476028 135584
rect 475528 135544 476028 135572
rect 475528 135532 475534 135544
rect 476022 135532 476028 135544
rect 476080 135532 476086 135584
rect 478046 135532 478052 135584
rect 478104 135572 478110 135584
rect 478782 135572 478788 135584
rect 478104 135544 478788 135572
rect 478104 135532 478110 135544
rect 478782 135532 478788 135544
rect 478840 135532 478846 135584
rect 519538 135572 519544 135584
rect 478892 135544 519544 135572
rect 466052 135476 469352 135504
rect 466052 135464 466058 135476
rect 473814 135464 473820 135516
rect 473872 135504 473878 135516
rect 473872 135476 476344 135504
rect 473872 135464 473878 135476
rect 475378 135436 475384 135448
rect 452948 135408 475384 135436
rect 475378 135396 475384 135408
rect 475436 135396 475442 135448
rect 476316 135436 476344 135476
rect 476390 135464 476396 135516
rect 476448 135504 476454 135516
rect 478892 135504 478920 135544
rect 519538 135532 519544 135544
rect 519596 135532 519602 135584
rect 515398 135504 515404 135516
rect 476448 135476 478920 135504
rect 480226 135476 515404 135504
rect 476448 135464 476454 135476
rect 480226 135436 480254 135476
rect 515398 135464 515404 135476
rect 515456 135464 515462 135516
rect 476316 135408 480254 135436
rect 480441 135439 480499 135445
rect 480441 135405 480453 135439
rect 480487 135436 480499 135439
rect 485038 135436 485044 135448
rect 480487 135408 485044 135436
rect 480487 135405 480499 135408
rect 480441 135399 480499 135405
rect 485038 135396 485044 135408
rect 485096 135396 485102 135448
rect 496170 135396 496176 135448
rect 496228 135436 496234 135448
rect 496722 135436 496728 135448
rect 496228 135408 496728 135436
rect 496228 135396 496234 135408
rect 496722 135396 496728 135408
rect 496780 135396 496786 135448
rect 496817 135439 496875 135445
rect 496817 135405 496829 135439
rect 496863 135436 496875 135439
rect 499574 135436 499580 135448
rect 496863 135408 499580 135436
rect 496863 135405 496875 135408
rect 496817 135399 496875 135405
rect 499574 135396 499580 135408
rect 499632 135396 499638 135448
rect 501322 135396 501328 135448
rect 501380 135436 501386 135448
rect 502150 135436 502156 135448
rect 501380 135408 502156 135436
rect 501380 135396 501386 135408
rect 502150 135396 502156 135408
rect 502208 135396 502214 135448
rect 503070 135396 503076 135448
rect 503128 135436 503134 135448
rect 503622 135436 503628 135448
rect 503128 135408 503628 135436
rect 503128 135396 503134 135408
rect 503622 135396 503628 135408
rect 503680 135396 503686 135448
rect 503898 135396 503904 135448
rect 503956 135436 503962 135448
rect 505002 135436 505008 135448
rect 503956 135408 505008 135436
rect 503956 135396 503962 135408
rect 505002 135396 505008 135408
rect 505060 135396 505066 135448
rect 79318 135328 79324 135380
rect 79376 135368 79382 135380
rect 88702 135368 88708 135380
rect 79376 135340 88708 135368
rect 79376 135328 79382 135340
rect 88702 135328 88708 135340
rect 88760 135328 88766 135380
rect 228358 135328 228364 135380
rect 228416 135368 228422 135380
rect 241146 135368 241152 135380
rect 228416 135340 241152 135368
rect 228416 135328 228422 135340
rect 241146 135328 241152 135340
rect 241204 135328 241210 135380
rect 379882 135328 379888 135380
rect 379940 135368 379946 135380
rect 380802 135368 380808 135380
rect 379940 135340 380808 135368
rect 379940 135328 379946 135340
rect 380802 135328 380808 135340
rect 380860 135328 380866 135380
rect 480349 135371 480407 135377
rect 480349 135337 480361 135371
rect 480395 135368 480407 135371
rect 482278 135368 482284 135380
rect 480395 135340 482284 135368
rect 480395 135337 480407 135340
rect 480349 135331 480407 135337
rect 482278 135328 482284 135340
rect 482336 135328 482342 135380
rect 498746 135328 498752 135380
rect 498804 135368 498810 135380
rect 499482 135368 499488 135380
rect 498804 135340 499488 135368
rect 498804 135328 498810 135340
rect 499482 135328 499488 135340
rect 499540 135328 499546 135380
rect 231118 135260 231124 135312
rect 231176 135300 231182 135312
rect 239398 135300 239404 135312
rect 231176 135272 239404 135300
rect 231176 135260 231182 135272
rect 239398 135260 239404 135272
rect 239456 135260 239462 135312
rect 410058 135260 410064 135312
rect 410116 135300 410122 135312
rect 411162 135300 411168 135312
rect 410116 135272 411168 135300
rect 410116 135260 410122 135272
rect 411162 135260 411168 135272
rect 411220 135260 411226 135312
rect 411806 135260 411812 135312
rect 411864 135300 411870 135312
rect 412450 135300 412456 135312
rect 411864 135272 412456 135300
rect 411864 135260 411870 135272
rect 412450 135260 412456 135272
rect 412508 135260 412514 135312
rect 413462 135260 413468 135312
rect 413520 135300 413526 135312
rect 413922 135300 413928 135312
rect 413520 135272 413928 135300
rect 413520 135260 413526 135272
rect 413922 135260 413928 135272
rect 413980 135260 413986 135312
rect 416038 135260 416044 135312
rect 416096 135300 416102 135312
rect 416682 135300 416688 135312
rect 416096 135272 416688 135300
rect 416096 135260 416102 135272
rect 416682 135260 416688 135272
rect 416740 135260 416746 135312
rect 458266 135260 458272 135312
rect 458324 135300 458330 135312
rect 459370 135300 459376 135312
rect 458324 135272 459376 135300
rect 458324 135260 458330 135272
rect 459370 135260 459376 135272
rect 459428 135260 459434 135312
rect 460014 135260 460020 135312
rect 460072 135300 460078 135312
rect 460842 135300 460848 135312
rect 460072 135272 460848 135300
rect 460072 135260 460078 135272
rect 460842 135260 460848 135272
rect 460900 135260 460906 135312
rect 461670 135260 461676 135312
rect 461728 135300 461734 135312
rect 462222 135300 462228 135312
rect 461728 135272 462228 135300
rect 461728 135260 461734 135272
rect 462222 135260 462228 135272
rect 462280 135260 462286 135312
rect 464338 135260 464344 135312
rect 464396 135300 464402 135312
rect 464982 135300 464988 135312
rect 464396 135272 464988 135300
rect 464396 135260 464402 135272
rect 464982 135260 464988 135272
rect 465040 135260 465046 135312
rect 465166 135260 465172 135312
rect 465224 135300 465230 135312
rect 466362 135300 466368 135312
rect 465224 135272 466368 135300
rect 465224 135260 465230 135272
rect 466362 135260 466368 135272
rect 466420 135260 466426 135312
rect 481450 135260 481456 135312
rect 481508 135300 481514 135312
rect 488626 135300 488632 135312
rect 481508 135272 488632 135300
rect 481508 135260 481514 135272
rect 488626 135260 488632 135272
rect 488684 135260 488690 135312
rect 43438 135124 43444 135176
rect 43496 135164 43502 135176
rect 96430 135164 96436 135176
rect 43496 135136 96436 135164
rect 43496 135124 43502 135136
rect 96430 135124 96436 135136
rect 96488 135124 96494 135176
rect 22002 135056 22008 135108
rect 22060 135096 22066 135108
rect 76926 135096 76932 135108
rect 22060 135068 76932 135096
rect 22060 135056 22066 135068
rect 76926 135056 76932 135068
rect 76984 135056 76990 135108
rect 77202 135056 77208 135108
rect 77260 135096 77266 135108
rect 135162 135096 135168 135108
rect 77260 135068 135168 135096
rect 77260 135056 77266 135068
rect 135162 135056 135168 135068
rect 135220 135056 135226 135108
rect 53742 134988 53748 135040
rect 53800 135028 53806 135040
rect 115290 135028 115296 135040
rect 53800 135000 115296 135028
rect 53800 134988 53806 135000
rect 115290 134988 115296 135000
rect 115348 134988 115354 135040
rect 487522 134988 487528 135040
rect 487580 135028 487586 135040
rect 547138 135028 547144 135040
rect 487580 135000 547144 135028
rect 487580 134988 487586 135000
rect 547138 134988 547144 135000
rect 547196 134988 547202 135040
rect 62022 134920 62028 134972
rect 62080 134960 62086 134972
rect 124858 134960 124864 134972
rect 62080 134932 124864 134960
rect 62080 134920 62086 134932
rect 124858 134920 124864 134932
rect 124916 134920 124922 134972
rect 459094 134920 459100 134972
rect 459152 134960 459158 134972
rect 520274 134960 520280 134972
rect 459152 134932 520280 134960
rect 459152 134920 459158 134932
rect 520274 134920 520280 134932
rect 520332 134920 520338 134972
rect 41322 134852 41328 134904
rect 41380 134892 41386 134904
rect 104158 134892 104164 134904
rect 41380 134864 104164 134892
rect 41380 134852 41386 134864
rect 104158 134852 104164 134864
rect 104216 134852 104222 134904
rect 488626 134852 488632 134904
rect 488684 134892 488690 134904
rect 550634 134892 550640 134904
rect 488684 134864 550640 134892
rect 488684 134852 488690 134864
rect 550634 134852 550640 134864
rect 550692 134852 550698 134904
rect 39390 134784 39396 134836
rect 39448 134824 39454 134836
rect 102502 134824 102508 134836
rect 39448 134796 102508 134824
rect 39448 134784 39454 134796
rect 102502 134784 102508 134796
rect 102560 134784 102566 134836
rect 477218 134784 477224 134836
rect 477276 134824 477282 134836
rect 544378 134824 544384 134836
rect 477276 134796 544384 134824
rect 477276 134784 477282 134796
rect 544378 134784 544384 134796
rect 544436 134784 544442 134836
rect 35158 134716 35164 134768
rect 35216 134756 35222 134768
rect 99926 134756 99932 134768
rect 35216 134728 99932 134756
rect 35216 134716 35222 134728
rect 99926 134716 99932 134728
rect 99984 134716 99990 134768
rect 478966 134716 478972 134768
rect 479024 134756 479030 134768
rect 547874 134756 547880 134768
rect 479024 134728 547880 134756
rect 479024 134716 479030 134728
rect 547874 134716 547880 134728
rect 547932 134716 547938 134768
rect 37182 134648 37188 134700
rect 37240 134688 37246 134700
rect 106826 134688 106832 134700
rect 37240 134660 106832 134688
rect 37240 134648 37246 134660
rect 106826 134648 106832 134660
rect 106884 134648 106890 134700
rect 484118 134648 484124 134700
rect 484176 134688 484182 134700
rect 554774 134688 554780 134700
rect 484176 134660 554780 134688
rect 484176 134648 484182 134660
rect 554774 134648 554780 134660
rect 554832 134648 554838 134700
rect 15838 134580 15844 134632
rect 15896 134620 15902 134632
rect 89530 134620 89536 134632
rect 15896 134592 89536 134620
rect 15896 134580 15902 134592
rect 89530 134580 89536 134592
rect 89588 134580 89594 134632
rect 135162 134580 135168 134632
rect 135220 134620 135226 134632
rect 177390 134620 177396 134632
rect 135220 134592 177396 134620
rect 135220 134580 135226 134592
rect 177390 134580 177396 134592
rect 177448 134580 177454 134632
rect 493870 134580 493876 134632
rect 493928 134620 493934 134632
rect 564526 134620 564532 134632
rect 493928 134592 564532 134620
rect 493928 134580 493934 134592
rect 564526 134580 564532 134592
rect 564584 134580 564590 134632
rect 11698 134512 11704 134564
rect 11756 134552 11762 134564
rect 86126 134552 86132 134564
rect 11756 134524 86132 134552
rect 11756 134512 11762 134524
rect 86126 134512 86132 134524
rect 86184 134512 86190 134564
rect 91002 134512 91008 134564
rect 91060 134552 91066 134564
rect 140774 134552 140780 134564
rect 91060 134524 140780 134552
rect 91060 134512 91066 134524
rect 140774 134512 140780 134524
rect 140832 134512 140838 134564
rect 142062 134512 142068 134564
rect 142120 134552 142126 134564
rect 182542 134552 182548 134564
rect 142120 134524 182548 134552
rect 142120 134512 142126 134524
rect 182542 134512 182548 134524
rect 182600 134512 182606 134564
rect 496998 134512 497004 134564
rect 497056 134552 497062 134564
rect 572806 134552 572812 134564
rect 497056 134524 572812 134552
rect 497056 134512 497062 134524
rect 572806 134512 572812 134524
rect 572864 134512 572870 134564
rect 57238 133152 57244 133204
rect 57296 133192 57302 133204
rect 105078 133192 105084 133204
rect 57296 133164 105084 133192
rect 57296 133152 57302 133164
rect 105078 133152 105084 133164
rect 105136 133152 105142 133204
rect 484946 133152 484952 133204
rect 485004 133192 485010 133204
rect 556246 133192 556252 133204
rect 485004 133164 556252 133192
rect 485004 133152 485010 133164
rect 556246 133152 556252 133164
rect 556304 133152 556310 133204
rect 511258 126896 511264 126948
rect 511316 126936 511322 126948
rect 580166 126936 580172 126948
rect 511316 126908 580172 126936
rect 511316 126896 511322 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 538858 113092 538864 113144
rect 538916 113132 538922 113144
rect 579798 113132 579804 113144
rect 538916 113104 579804 113132
rect 538916 113092 538922 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 58618 111772 58624 111784
rect 3200 111744 58624 111772
rect 3200 111732 3206 111744
rect 58618 111732 58624 111744
rect 58676 111732 58682 111784
rect 560938 100648 560944 100700
rect 560996 100688 561002 100700
rect 580166 100688 580172 100700
rect 560996 100660 580172 100688
rect 560996 100648 561002 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 22738 97968 22744 97980
rect 3568 97940 22744 97968
rect 3568 97928 3574 97940
rect 22738 97928 22744 97940
rect 22796 97928 22802 97980
rect 508498 86912 508504 86964
rect 508556 86952 508562 86964
rect 580166 86952 580172 86964
rect 508556 86924 580172 86952
rect 508556 86912 508562 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 25498 85524 25504 85536
rect 3568 85496 25504 85524
rect 3568 85484 3574 85496
rect 25498 85484 25504 85496
rect 25556 85484 25562 85536
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 69658 71720 69664 71732
rect 3568 71692 69664 71720
rect 3568 71680 3574 71692
rect 69658 71680 69664 71692
rect 69716 71680 69722 71732
rect 70302 71000 70308 71052
rect 70360 71040 70366 71052
rect 130930 71040 130936 71052
rect 70360 71012 130936 71040
rect 70360 71000 70366 71012
rect 130930 71000 130936 71012
rect 130988 71000 130994 71052
rect 558178 60664 558184 60716
rect 558236 60704 558242 60716
rect 580166 60704 580172 60716
rect 558236 60676 580172 60704
rect 558236 60664 558242 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 473262 48968 473268 49020
rect 473320 49008 473326 49020
rect 538214 49008 538220 49020
rect 473320 48980 538220 49008
rect 473320 48968 473326 48980
rect 538214 48968 538220 48980
rect 538272 48968 538278 49020
rect 446950 47540 446956 47592
rect 447008 47580 447014 47592
rect 502334 47580 502340 47592
rect 447008 47552 502340 47580
rect 447008 47540 447014 47552
rect 502334 47540 502340 47552
rect 502392 47540 502398 47592
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 39298 45540 39304 45552
rect 3476 45512 39304 45540
rect 3476 45500 3482 45512
rect 39298 45500 39304 45512
rect 39356 45500 39362 45552
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 50338 33096 50344 33108
rect 3200 33068 50344 33096
rect 3200 33056 3206 33068
rect 50338 33056 50344 33068
rect 50396 33056 50402 33108
rect 50430 32376 50436 32428
rect 50488 32416 50494 32428
rect 107654 32416 107660 32428
rect 50488 32388 107660 32416
rect 50488 32376 50494 32388
rect 107654 32376 107660 32388
rect 107712 32376 107718 32428
rect 35250 26868 35256 26920
rect 35308 26908 35314 26920
rect 104250 26908 104256 26920
rect 35308 26880 104256 26908
rect 35308 26868 35314 26880
rect 104250 26868 104256 26880
rect 104308 26868 104314 26920
rect 104802 25508 104808 25560
rect 104860 25548 104866 25560
rect 155862 25548 155868 25560
rect 104860 25520 155868 25548
rect 104860 25508 104866 25520
rect 155862 25508 155868 25520
rect 155920 25508 155926 25560
rect 97902 24080 97908 24132
rect 97960 24120 97966 24132
rect 150710 24120 150716 24132
rect 97960 24092 150716 24120
rect 97960 24080 97966 24092
rect 150710 24080 150716 24092
rect 150768 24080 150774 24132
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 14458 20652 14464 20664
rect 3476 20624 14464 20652
rect 3476 20612 3482 20624
rect 14458 20612 14464 20624
rect 14516 20612 14522 20664
rect 368382 15852 368388 15904
rect 368440 15892 368446 15904
rect 395246 15892 395252 15904
rect 368440 15864 395252 15892
rect 368440 15852 368446 15864
rect 395246 15852 395252 15864
rect 395304 15852 395310 15904
rect 436002 15852 436008 15904
rect 436060 15892 436066 15904
rect 488810 15892 488816 15904
rect 436060 15864 488816 15892
rect 436060 15852 436066 15864
rect 488810 15852 488816 15864
rect 488868 15852 488874 15904
rect 489822 15852 489828 15904
rect 489880 15892 489886 15904
rect 562042 15892 562048 15904
rect 489880 15864 562048 15892
rect 489880 15852 489886 15864
rect 562042 15852 562048 15864
rect 562100 15852 562106 15904
rect 381538 14424 381544 14476
rect 381596 14464 381602 14476
rect 412634 14464 412640 14476
rect 381596 14436 412640 14464
rect 381596 14424 381602 14436
rect 412634 14424 412640 14436
rect 412692 14424 412698 14476
rect 471882 14424 471888 14476
rect 471940 14464 471946 14476
rect 537202 14464 537208 14476
rect 471940 14436 537208 14464
rect 471940 14424 471946 14436
rect 537202 14424 537208 14436
rect 537260 14424 537266 14476
rect 376570 11704 376576 11756
rect 376628 11744 376634 11756
rect 406010 11744 406016 11756
rect 376628 11716 406016 11744
rect 376628 11704 376634 11716
rect 406010 11704 406016 11716
rect 406068 11704 406074 11756
rect 406378 11704 406384 11756
rect 406436 11744 406442 11756
rect 445754 11744 445760 11756
rect 406436 11716 445760 11744
rect 406436 11704 406442 11716
rect 445754 11704 445760 11716
rect 445812 11704 445818 11756
rect 449802 11704 449808 11756
rect 449860 11744 449866 11756
rect 506566 11744 506572 11756
rect 449860 11716 506572 11744
rect 449860 11704 449866 11716
rect 506566 11704 506572 11716
rect 506624 11704 506630 11756
rect 512638 11704 512644 11756
rect 512696 11744 512702 11756
rect 530118 11744 530124 11756
rect 512696 11716 530124 11744
rect 512696 11704 512702 11716
rect 530118 11704 530124 11716
rect 530176 11704 530182 11756
rect 526438 10276 526444 10328
rect 526496 10316 526502 10328
rect 575842 10316 575848 10328
rect 526496 10288 575848 10316
rect 526496 10276 526502 10288
rect 575842 10276 575848 10288
rect 575900 10276 575906 10328
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 75178 8956 75184 8968
rect 4120 8928 75184 8956
rect 4120 8916 4126 8928
rect 75178 8916 75184 8928
rect 75236 8916 75242 8968
rect 83274 8916 83280 8968
rect 83332 8956 83338 8968
rect 137278 8956 137284 8968
rect 83332 8928 137284 8956
rect 83332 8916 83338 8928
rect 137278 8916 137284 8928
rect 137336 8916 137342 8968
rect 137646 8916 137652 8968
rect 137704 8956 137710 8968
rect 179966 8956 179972 8968
rect 137704 8928 179972 8956
rect 137704 8916 137710 8928
rect 179966 8916 179972 8928
rect 180024 8916 180030 8968
rect 363598 8916 363604 8968
rect 363656 8956 363662 8968
rect 388254 8956 388260 8968
rect 363656 8928 388260 8956
rect 363656 8916 363662 8928
rect 388254 8916 388260 8928
rect 388312 8916 388318 8968
rect 469122 8916 469128 8968
rect 469180 8956 469186 8968
rect 533706 8956 533712 8968
rect 469180 8928 533712 8956
rect 469180 8916 469186 8928
rect 533706 8916 533712 8928
rect 533764 8916 533770 8968
rect 132954 7692 132960 7744
rect 133012 7732 133018 7744
rect 146938 7732 146944 7744
rect 133012 7704 146944 7732
rect 133012 7692 133018 7704
rect 146938 7692 146944 7704
rect 146996 7692 147002 7744
rect 115198 7624 115204 7676
rect 115256 7664 115262 7676
rect 133138 7664 133144 7676
rect 115256 7636 133144 7664
rect 115256 7624 115262 7636
rect 133138 7624 133144 7636
rect 133196 7624 133202 7676
rect 147122 7624 147128 7676
rect 147180 7664 147186 7676
rect 186866 7664 186872 7676
rect 147180 7636 186872 7664
rect 147180 7624 147186 7636
rect 186866 7624 186872 7636
rect 186924 7624 186930 7676
rect 397270 7624 397276 7676
rect 397328 7664 397334 7676
rect 435542 7664 435548 7676
rect 397328 7636 435548 7664
rect 397328 7624 397334 7636
rect 435542 7624 435548 7636
rect 435600 7624 435606 7676
rect 520918 7624 520924 7676
rect 520976 7664 520982 7676
rect 558546 7664 558552 7676
rect 520976 7636 558552 7664
rect 520976 7624 520982 7636
rect 558546 7624 558552 7636
rect 558604 7624 558610 7676
rect 12342 7556 12348 7608
rect 12400 7596 12406 7608
rect 79318 7596 79324 7608
rect 12400 7568 79324 7596
rect 12400 7556 12406 7568
rect 79318 7556 79324 7568
rect 79376 7556 79382 7608
rect 111610 7556 111616 7608
rect 111668 7596 111674 7608
rect 161014 7596 161020 7608
rect 111668 7568 161020 7596
rect 111668 7556 111674 7568
rect 161014 7556 161020 7568
rect 161072 7556 161078 7608
rect 358630 7556 358636 7608
rect 358688 7596 358694 7608
rect 381170 7596 381176 7608
rect 358688 7568 381176 7596
rect 358688 7556 358694 7568
rect 381170 7556 381176 7568
rect 381228 7556 381234 7608
rect 419350 7556 419356 7608
rect 419408 7596 419414 7608
rect 466270 7596 466276 7608
rect 419408 7568 466276 7596
rect 419408 7556 419414 7568
rect 466270 7556 466276 7568
rect 466328 7556 466334 7608
rect 522298 7556 522304 7608
rect 522356 7596 522362 7608
rect 569126 7596 569132 7608
rect 522356 7568 569132 7596
rect 522356 7556 522362 7568
rect 569126 7556 569132 7568
rect 569184 7556 569190 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 33778 6848 33784 6860
rect 3476 6820 33784 6848
rect 3476 6808 3482 6820
rect 33778 6808 33784 6820
rect 33836 6808 33842 6860
rect 431770 6604 431776 6656
rect 431828 6644 431834 6656
rect 481726 6644 481732 6656
rect 431828 6616 481732 6644
rect 431828 6604 431834 6616
rect 481726 6604 481732 6616
rect 481784 6604 481790 6656
rect 433242 6536 433248 6588
rect 433300 6576 433306 6588
rect 485222 6576 485228 6588
rect 433300 6548 485228 6576
rect 433300 6536 433306 6548
rect 485222 6536 485228 6548
rect 485280 6536 485286 6588
rect 144730 6468 144736 6520
rect 144788 6508 144794 6520
rect 180058 6508 180064 6520
rect 144788 6480 180064 6508
rect 144788 6468 144794 6480
rect 180058 6468 180064 6480
rect 180116 6468 180122 6520
rect 464338 6468 464344 6520
rect 464396 6508 464402 6520
rect 517146 6508 517152 6520
rect 464396 6480 517152 6508
rect 464396 6468 464402 6480
rect 517146 6468 517152 6480
rect 517204 6468 517210 6520
rect 138842 6400 138848 6452
rect 138900 6440 138906 6452
rect 180886 6440 180892 6452
rect 138900 6412 180892 6440
rect 138900 6400 138906 6412
rect 180886 6400 180892 6412
rect 180944 6400 180950 6452
rect 443638 6400 443644 6452
rect 443696 6440 443702 6452
rect 495894 6440 495900 6452
rect 443696 6412 495900 6440
rect 443696 6400 443702 6412
rect 495894 6400 495900 6412
rect 495952 6400 495958 6452
rect 519538 6400 519544 6452
rect 519596 6440 519602 6452
rect 544286 6440 544292 6452
rect 519596 6412 544292 6440
rect 519596 6400 519602 6412
rect 544286 6400 544292 6412
rect 544344 6400 544350 6452
rect 122374 6332 122380 6384
rect 122432 6372 122438 6384
rect 168834 6372 168840 6384
rect 122432 6344 168840 6372
rect 122432 6332 122438 6344
rect 168834 6332 168840 6344
rect 168892 6332 168898 6384
rect 462222 6332 462228 6384
rect 462280 6372 462286 6384
rect 524230 6372 524236 6384
rect 462280 6344 524236 6372
rect 462280 6332 462286 6344
rect 524230 6332 524236 6344
rect 524288 6332 524294 6384
rect 118786 6264 118792 6316
rect 118844 6304 118850 6316
rect 166258 6304 166264 6316
rect 118844 6276 166264 6304
rect 118844 6264 118850 6276
rect 166258 6264 166264 6276
rect 166316 6264 166322 6316
rect 464982 6264 464988 6316
rect 465040 6304 465046 6316
rect 527818 6304 527824 6316
rect 465040 6276 527824 6304
rect 465040 6264 465046 6276
rect 527818 6264 527824 6276
rect 527876 6264 527882 6316
rect 108114 6196 108120 6248
rect 108172 6236 108178 6248
rect 158438 6236 158444 6248
rect 108172 6208 158444 6236
rect 108172 6196 108178 6208
rect 158438 6196 158444 6208
rect 158496 6196 158502 6248
rect 467742 6196 467748 6248
rect 467800 6236 467806 6248
rect 531314 6236 531320 6248
rect 467800 6208 531320 6236
rect 467800 6196 467806 6208
rect 531314 6196 531320 6208
rect 531372 6196 531378 6248
rect 69106 6128 69112 6180
rect 69164 6168 69170 6180
rect 83458 6168 83464 6180
rect 69164 6140 83464 6168
rect 69164 6128 69170 6140
rect 83458 6128 83464 6140
rect 83516 6128 83522 6180
rect 86862 6128 86868 6180
rect 86920 6168 86926 6180
rect 142982 6168 142988 6180
rect 86920 6140 142988 6168
rect 86920 6128 86926 6140
rect 142982 6128 142988 6140
rect 143040 6128 143046 6180
rect 183462 6168 183468 6180
rect 151786 6140 183468 6168
rect 142430 6060 142436 6112
rect 142488 6100 142494 6112
rect 151786 6100 151814 6140
rect 183462 6128 183468 6140
rect 183520 6128 183526 6180
rect 436738 6128 436744 6180
rect 436796 6168 436802 6180
rect 476942 6168 476948 6180
rect 436796 6140 476948 6168
rect 436796 6128 436802 6140
rect 476942 6128 476948 6140
rect 477000 6128 477006 6180
rect 480070 6128 480076 6180
rect 480128 6168 480134 6180
rect 549070 6168 549076 6180
rect 480128 6140 549076 6168
rect 480128 6128 480134 6140
rect 549070 6128 549076 6140
rect 549128 6128 549134 6180
rect 142488 6072 151814 6100
rect 142488 6060 142494 6072
rect 59630 5448 59636 5500
rect 59688 5488 59694 5500
rect 72418 5488 72424 5500
rect 59688 5460 72424 5488
rect 59688 5448 59694 5460
rect 72418 5448 72424 5460
rect 72476 5448 72482 5500
rect 72602 5448 72608 5500
rect 72660 5488 72666 5500
rect 132678 5488 132684 5500
rect 72660 5460 132684 5488
rect 72660 5448 72666 5460
rect 132678 5448 132684 5460
rect 132736 5448 132742 5500
rect 161290 5448 161296 5500
rect 161348 5488 161354 5500
rect 197262 5488 197268 5500
rect 161348 5460 197268 5488
rect 161348 5448 161354 5460
rect 197262 5448 197268 5460
rect 197320 5448 197326 5500
rect 438762 5448 438768 5500
rect 438820 5488 438826 5500
rect 491018 5488 491024 5500
rect 438820 5460 491024 5488
rect 438820 5448 438826 5460
rect 491018 5448 491024 5460
rect 491076 5448 491082 5500
rect 65610 5380 65616 5432
rect 65668 5420 65674 5432
rect 127434 5420 127440 5432
rect 65668 5392 127440 5420
rect 65668 5380 65674 5392
rect 127434 5380 127440 5392
rect 127492 5380 127498 5432
rect 135254 5380 135260 5432
rect 135312 5420 135318 5432
rect 178310 5420 178316 5432
rect 135312 5392 178316 5420
rect 135312 5380 135318 5392
rect 178310 5380 178316 5392
rect 178368 5380 178374 5432
rect 414658 5380 414664 5432
rect 414716 5420 414722 5432
rect 428458 5420 428464 5432
rect 414716 5392 428464 5420
rect 414716 5380 414722 5392
rect 428458 5380 428464 5392
rect 428516 5380 428522 5432
rect 440050 5380 440056 5432
rect 440108 5420 440114 5432
rect 494698 5420 494704 5432
rect 440108 5392 494704 5420
rect 440108 5380 440114 5392
rect 494698 5380 494704 5392
rect 494756 5380 494762 5432
rect 56042 5312 56048 5364
rect 56100 5352 56106 5364
rect 65518 5352 65524 5364
rect 56100 5324 65524 5352
rect 56100 5312 56106 5324
rect 65518 5312 65524 5324
rect 65576 5312 65582 5364
rect 66714 5312 66720 5364
rect 66772 5352 66778 5364
rect 128354 5352 128360 5364
rect 66772 5324 128360 5352
rect 66772 5312 66778 5324
rect 128354 5312 128360 5324
rect 128412 5312 128418 5364
rect 129366 5312 129372 5364
rect 129424 5352 129430 5364
rect 170398 5352 170404 5364
rect 129424 5324 170404 5352
rect 129424 5312 129430 5324
rect 170398 5312 170404 5324
rect 170456 5312 170462 5364
rect 407758 5312 407764 5364
rect 407816 5352 407822 5364
rect 420178 5352 420184 5364
rect 407816 5324 420184 5352
rect 407816 5312 407822 5324
rect 420178 5312 420184 5324
rect 420236 5312 420242 5364
rect 421558 5312 421564 5364
rect 421616 5352 421622 5364
rect 442626 5352 442632 5364
rect 421616 5324 442632 5352
rect 421616 5312 421622 5324
rect 442626 5312 442632 5324
rect 442684 5312 442690 5364
rect 445662 5312 445668 5364
rect 445720 5352 445726 5364
rect 501782 5352 501788 5364
rect 445720 5324 501788 5352
rect 445720 5312 445726 5324
rect 501782 5312 501788 5324
rect 501840 5312 501846 5364
rect 58434 5244 58440 5296
rect 58492 5284 58498 5296
rect 122282 5284 122288 5296
rect 58492 5256 122288 5284
rect 58492 5244 58498 5256
rect 122282 5244 122288 5256
rect 122340 5244 122346 5296
rect 136450 5244 136456 5296
rect 136508 5284 136514 5296
rect 179138 5284 179144 5296
rect 136508 5256 179144 5284
rect 136508 5244 136514 5256
rect 179138 5244 179144 5256
rect 179196 5244 179202 5296
rect 399478 5244 399484 5296
rect 399536 5284 399542 5296
rect 427262 5284 427268 5296
rect 399536 5256 427268 5284
rect 399536 5244 399542 5256
rect 427262 5244 427268 5256
rect 427320 5244 427326 5296
rect 442810 5244 442816 5296
rect 442868 5284 442874 5296
rect 498194 5284 498200 5296
rect 442868 5256 498200 5284
rect 442868 5244 442874 5256
rect 498194 5244 498200 5256
rect 498252 5244 498258 5296
rect 44266 5176 44272 5228
rect 44324 5216 44330 5228
rect 54478 5216 54484 5228
rect 44324 5188 54484 5216
rect 44324 5176 44330 5188
rect 54478 5176 54484 5188
rect 54536 5176 54542 5228
rect 54938 5176 54944 5228
rect 54996 5216 55002 5228
rect 119706 5216 119712 5228
rect 54996 5188 119712 5216
rect 54996 5176 55002 5188
rect 119706 5176 119712 5188
rect 119764 5176 119770 5228
rect 131758 5176 131764 5228
rect 131816 5216 131822 5228
rect 175734 5216 175740 5228
rect 131816 5188 175740 5216
rect 131816 5176 131822 5188
rect 175734 5176 175740 5188
rect 175792 5176 175798 5228
rect 383470 5176 383476 5228
rect 383528 5216 383534 5228
rect 416682 5216 416688 5228
rect 383528 5188 416688 5216
rect 383528 5176 383534 5188
rect 416682 5176 416688 5188
rect 416740 5176 416746 5228
rect 417418 5176 417424 5228
rect 417476 5216 417482 5228
rect 439130 5216 439136 5228
rect 417476 5188 439136 5216
rect 417476 5176 417482 5188
rect 439130 5176 439136 5188
rect 439188 5176 439194 5228
rect 448422 5176 448428 5228
rect 448480 5216 448486 5228
rect 505370 5216 505376 5228
rect 448480 5188 505376 5216
rect 448480 5176 448486 5188
rect 505370 5176 505376 5188
rect 505428 5176 505434 5228
rect 51350 5108 51356 5160
rect 51408 5148 51414 5160
rect 117130 5148 117136 5160
rect 51408 5120 117136 5148
rect 51408 5108 51414 5120
rect 117130 5108 117136 5120
rect 117188 5108 117194 5160
rect 130562 5108 130568 5160
rect 130620 5148 130626 5160
rect 174814 5148 174820 5160
rect 130620 5120 174820 5148
rect 130620 5108 130626 5120
rect 174814 5108 174820 5120
rect 174872 5108 174878 5160
rect 389082 5108 389088 5160
rect 389140 5148 389146 5160
rect 423766 5148 423772 5160
rect 389140 5120 423772 5148
rect 389140 5108 389146 5120
rect 423766 5108 423772 5120
rect 423824 5108 423830 5160
rect 429838 5108 429844 5160
rect 429896 5148 429902 5160
rect 437934 5148 437940 5160
rect 429896 5120 437940 5148
rect 429896 5108 429902 5120
rect 437934 5108 437940 5120
rect 437992 5108 437998 5160
rect 451182 5108 451188 5160
rect 451240 5148 451246 5160
rect 508866 5148 508872 5160
rect 451240 5120 508872 5148
rect 451240 5108 451246 5120
rect 508866 5108 508872 5120
rect 508924 5108 508930 5160
rect 30098 5040 30104 5092
rect 30156 5080 30162 5092
rect 47578 5080 47584 5092
rect 30156 5052 47584 5080
rect 30156 5040 30162 5052
rect 47578 5040 47584 5052
rect 47636 5040 47642 5092
rect 47854 5040 47860 5092
rect 47912 5080 47918 5092
rect 114554 5080 114560 5092
rect 47912 5052 114560 5080
rect 47912 5040 47918 5052
rect 114554 5040 114560 5052
rect 114612 5040 114618 5092
rect 125870 5040 125876 5092
rect 125928 5080 125934 5092
rect 170490 5080 170496 5092
rect 125928 5052 170496 5080
rect 125928 5040 125934 5052
rect 170490 5040 170496 5052
rect 170548 5040 170554 5092
rect 171962 5040 171968 5092
rect 172020 5080 172026 5092
rect 191098 5080 191104 5092
rect 172020 5052 191104 5080
rect 172020 5040 172026 5052
rect 191098 5040 191104 5052
rect 191156 5040 191162 5092
rect 397362 5040 397368 5092
rect 397420 5080 397426 5092
rect 426989 5083 427047 5089
rect 426989 5080 427001 5083
rect 397420 5052 427001 5080
rect 397420 5040 397426 5052
rect 426989 5049 427001 5052
rect 427035 5049 427047 5083
rect 432046 5080 432052 5092
rect 426989 5043 427047 5049
rect 427096 5052 432052 5080
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 85298 5012 85304 5024
rect 7708 4984 85304 5012
rect 7708 4972 7714 4984
rect 85298 4972 85304 4984
rect 85356 4972 85362 5024
rect 128170 4972 128176 5024
rect 128228 5012 128234 5024
rect 173066 5012 173072 5024
rect 128228 4984 173072 5012
rect 128228 4972 128234 4984
rect 173066 4972 173072 4984
rect 173124 4972 173130 5024
rect 394602 4972 394608 5024
rect 394660 5012 394666 5024
rect 427096 5012 427124 5052
rect 432046 5040 432052 5052
rect 432104 5040 432110 5092
rect 453942 5040 453948 5092
rect 454000 5080 454006 5092
rect 512454 5080 512460 5092
rect 454000 5052 512460 5080
rect 454000 5040 454006 5052
rect 512454 5040 512460 5052
rect 512512 5040 512518 5092
rect 394660 4984 427124 5012
rect 394660 4972 394666 4984
rect 435358 4972 435364 5024
rect 435416 5012 435422 5024
rect 445018 5012 445024 5024
rect 435416 4984 445024 5012
rect 435416 4972 435422 4984
rect 445018 4972 445024 4984
rect 445076 4972 445082 5024
rect 456702 4972 456708 5024
rect 456760 5012 456766 5024
rect 456760 4984 515352 5012
rect 456760 4972 456766 4984
rect 1670 4904 1676 4956
rect 1728 4944 1734 4956
rect 80054 4944 80060 4956
rect 1728 4916 80060 4944
rect 1728 4904 1734 4916
rect 80054 4904 80060 4916
rect 80112 4904 80118 4956
rect 93946 4904 93952 4956
rect 94004 4944 94010 4956
rect 148134 4944 148140 4956
rect 94004 4916 148140 4944
rect 94004 4904 94010 4916
rect 148134 4904 148140 4916
rect 148192 4904 148198 4956
rect 157794 4904 157800 4956
rect 157852 4944 157858 4956
rect 194686 4944 194692 4956
rect 157852 4916 194692 4944
rect 157852 4904 157858 4916
rect 194686 4904 194692 4916
rect 194744 4904 194750 4956
rect 356698 4904 356704 4956
rect 356756 4944 356762 4956
rect 377674 4944 377680 4956
rect 356756 4916 377680 4944
rect 356756 4904 356762 4916
rect 377674 4904 377680 4916
rect 377732 4904 377738 4956
rect 401502 4904 401508 4956
rect 401560 4944 401566 4956
rect 441522 4944 441528 4956
rect 401560 4916 441528 4944
rect 401560 4904 401566 4916
rect 441522 4904 441528 4916
rect 441580 4904 441586 4956
rect 459370 4904 459376 4956
rect 459428 4944 459434 4956
rect 514021 4947 514079 4953
rect 514021 4944 514033 4947
rect 459428 4916 514033 4944
rect 459428 4904 459434 4916
rect 514021 4913 514033 4916
rect 514067 4913 514079 4947
rect 515324 4944 515352 4984
rect 515398 4972 515404 5024
rect 515456 5012 515462 5024
rect 540790 5012 540796 5024
rect 515456 4984 540796 5012
rect 515456 4972 515462 4984
rect 540790 4972 540796 4984
rect 540848 4972 540854 5024
rect 515950 4944 515956 4956
rect 515324 4916 515956 4944
rect 514021 4907 514079 4913
rect 515950 4904 515956 4916
rect 516008 4904 516014 4956
rect 2866 4836 2872 4888
rect 2924 4876 2930 4888
rect 81802 4876 81808 4888
rect 2924 4848 81808 4876
rect 2924 4836 2930 4848
rect 81802 4836 81808 4848
rect 81860 4836 81866 4888
rect 91554 4836 91560 4888
rect 91612 4876 91618 4888
rect 146386 4876 146392 4888
rect 91612 4848 146392 4876
rect 91612 4836 91618 4848
rect 146386 4836 146392 4848
rect 146444 4836 146450 4888
rect 150618 4836 150624 4888
rect 150676 4876 150682 4888
rect 188338 4876 188344 4888
rect 150676 4848 188344 4876
rect 150676 4836 150682 4848
rect 188338 4836 188344 4848
rect 188396 4836 188402 4888
rect 360010 4836 360016 4888
rect 360068 4876 360074 4888
rect 384758 4876 384764 4888
rect 360068 4848 384764 4876
rect 360068 4836 360074 4848
rect 384758 4836 384764 4848
rect 384816 4836 384822 4888
rect 407022 4836 407028 4888
rect 407080 4876 407086 4888
rect 448606 4876 448612 4888
rect 407080 4848 448612 4876
rect 407080 4836 407086 4848
rect 448606 4836 448612 4848
rect 448664 4836 448670 4888
rect 463602 4836 463608 4888
rect 463660 4876 463666 4888
rect 526622 4876 526628 4888
rect 463660 4848 526628 4876
rect 463660 4836 463666 4848
rect 526622 4836 526628 4848
rect 526680 4836 526686 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 80146 4808 80152 4820
rect 624 4780 80152 4808
rect 624 4768 630 4780
rect 80146 4768 80152 4780
rect 80204 4768 80210 4820
rect 84470 4768 84476 4820
rect 84528 4808 84534 4820
rect 141234 4808 141240 4820
rect 84528 4780 141240 4808
rect 84528 4768 84534 4780
rect 141234 4768 141240 4780
rect 141292 4768 141298 4820
rect 143534 4768 143540 4820
rect 143592 4808 143598 4820
rect 184290 4808 184296 4820
rect 143592 4780 184296 4808
rect 143592 4768 143598 4780
rect 184290 4768 184296 4780
rect 184348 4768 184354 4820
rect 371142 4768 371148 4820
rect 371200 4808 371206 4820
rect 398926 4808 398932 4820
rect 371200 4780 398932 4808
rect 371200 4768 371206 4780
rect 398926 4768 398932 4780
rect 398984 4768 398990 4820
rect 400858 4768 400864 4820
rect 400916 4808 400922 4820
rect 409598 4808 409604 4820
rect 400916 4780 409604 4808
rect 400916 4768 400922 4780
rect 409598 4768 409604 4780
rect 409656 4768 409662 4820
rect 412450 4768 412456 4820
rect 412508 4808 412514 4820
rect 455690 4808 455696 4820
rect 412508 4780 455696 4808
rect 412508 4768 412514 4780
rect 455690 4768 455696 4780
rect 455748 4768 455754 4820
rect 460750 4768 460756 4820
rect 460808 4808 460814 4820
rect 523034 4808 523040 4820
rect 460808 4780 523040 4808
rect 460808 4768 460814 4780
rect 523034 4768 523040 4780
rect 523092 4768 523098 4820
rect 536098 4768 536104 4820
rect 536156 4808 536162 4820
rect 541986 4808 541992 4820
rect 536156 4780 541992 4808
rect 536156 4768 536162 4780
rect 541986 4768 541992 4780
rect 542044 4768 542050 4820
rect 542998 4768 543004 4820
rect 543056 4808 543062 4820
rect 552658 4808 552664 4820
rect 543056 4780 552664 4808
rect 543056 4768 543062 4780
rect 552658 4768 552664 4780
rect 552716 4768 552722 4820
rect 63218 4700 63224 4752
rect 63276 4740 63282 4752
rect 68278 4740 68284 4752
rect 63276 4712 68284 4740
rect 63276 4700 63282 4712
rect 68278 4700 68284 4712
rect 68336 4700 68342 4752
rect 79686 4700 79692 4752
rect 79744 4740 79750 4752
rect 137830 4740 137836 4752
rect 79744 4712 137836 4740
rect 79744 4700 79750 4712
rect 137830 4700 137836 4712
rect 137888 4700 137894 4752
rect 154206 4700 154212 4752
rect 154264 4740 154270 4752
rect 186958 4740 186964 4752
rect 154264 4712 186964 4740
rect 154264 4700 154270 4712
rect 186958 4700 186964 4712
rect 187016 4700 187022 4752
rect 426989 4743 427047 4749
rect 426989 4709 427001 4743
rect 427035 4740 427047 4743
rect 434438 4740 434444 4752
rect 427035 4712 434444 4740
rect 427035 4709 427047 4712
rect 426989 4703 427047 4709
rect 434438 4700 434444 4712
rect 434496 4700 434502 4752
rect 475378 4700 475384 4752
rect 475436 4740 475442 4752
rect 499390 4740 499396 4752
rect 475436 4712 499396 4740
rect 475436 4700 475442 4712
rect 499390 4700 499396 4712
rect 499448 4700 499454 4752
rect 508590 4700 508596 4752
rect 508648 4740 508654 4752
rect 510062 4740 510068 4752
rect 508648 4712 510068 4740
rect 508648 4700 508654 4712
rect 510062 4700 510068 4712
rect 510120 4700 510126 4752
rect 514021 4743 514079 4749
rect 514021 4709 514033 4743
rect 514067 4740 514079 4743
rect 519538 4740 519544 4752
rect 514067 4712 519544 4740
rect 514067 4709 514079 4712
rect 514021 4703 514079 4709
rect 519538 4700 519544 4712
rect 519596 4700 519602 4752
rect 77386 4632 77392 4684
rect 77444 4672 77450 4684
rect 126238 4672 126244 4684
rect 77444 4644 126244 4672
rect 77444 4632 77450 4644
rect 126238 4632 126244 4644
rect 126296 4632 126302 4684
rect 126974 4632 126980 4684
rect 127032 4672 127038 4684
rect 142798 4672 142804 4684
rect 127032 4644 142804 4672
rect 127032 4632 127038 4644
rect 142798 4632 142804 4644
rect 142856 4632 142862 4684
rect 164878 4632 164884 4684
rect 164936 4672 164942 4684
rect 197998 4672 198004 4684
rect 164936 4644 198004 4672
rect 164936 4632 164942 4644
rect 197998 4632 198004 4644
rect 198056 4632 198062 4684
rect 457438 4632 457444 4684
rect 457496 4672 457502 4684
rect 480530 4672 480536 4684
rect 457496 4644 480536 4672
rect 457496 4632 457502 4644
rect 480530 4632 480536 4644
rect 480588 4632 480594 4684
rect 486418 4632 486424 4684
rect 486476 4672 486482 4684
rect 492306 4672 492312 4684
rect 486476 4644 492312 4672
rect 486476 4632 486482 4644
rect 492306 4632 492312 4644
rect 492364 4632 492370 4684
rect 101030 4564 101036 4616
rect 101088 4604 101094 4616
rect 130378 4604 130384 4616
rect 101088 4576 130384 4604
rect 101088 4564 101094 4576
rect 130378 4564 130384 4576
rect 130436 4564 130442 4616
rect 168374 4564 168380 4616
rect 168432 4604 168438 4616
rect 200758 4604 200764 4616
rect 168432 4576 200764 4604
rect 168432 4564 168438 4576
rect 200758 4564 200764 4576
rect 200816 4564 200822 4616
rect 140038 4496 140044 4548
rect 140096 4536 140102 4548
rect 144178 4536 144184 4548
rect 140096 4508 144184 4536
rect 140096 4496 140102 4508
rect 144178 4496 144184 4508
rect 144236 4496 144242 4548
rect 450538 4360 450544 4412
rect 450596 4400 450602 4412
rect 452102 4400 452108 4412
rect 450596 4372 452108 4400
rect 450596 4360 450602 4372
rect 452102 4360 452108 4372
rect 452160 4360 452166 4412
rect 26510 4156 26516 4208
rect 26568 4196 26574 4208
rect 32398 4196 32404 4208
rect 26568 4168 32404 4196
rect 26568 4156 26574 4168
rect 32398 4156 32404 4168
rect 32456 4156 32462 4208
rect 48958 4156 48964 4208
rect 49016 4196 49022 4208
rect 51718 4196 51724 4208
rect 49016 4168 51724 4196
rect 49016 4156 49022 4168
rect 51718 4156 51724 4168
rect 51776 4156 51782 4208
rect 85485 4199 85543 4205
rect 85485 4165 85497 4199
rect 85531 4196 85543 4199
rect 87046 4196 87052 4208
rect 85531 4168 87052 4196
rect 85531 4165 85543 4168
rect 85485 4159 85543 4165
rect 87046 4156 87052 4168
rect 87104 4156 87110 4208
rect 90269 4199 90327 4205
rect 90269 4165 90281 4199
rect 90315 4196 90327 4199
rect 94038 4196 94044 4208
rect 90315 4168 94044 4196
rect 90315 4165 90327 4168
rect 90269 4159 90327 4165
rect 94038 4156 94044 4168
rect 94096 4156 94102 4208
rect 106829 4199 106887 4205
rect 106829 4165 106841 4199
rect 106875 4196 106887 4199
rect 106875 4168 110368 4196
rect 106875 4165 106887 4168
rect 106829 4159 106887 4165
rect 41874 4088 41880 4140
rect 41932 4128 41938 4140
rect 110230 4128 110236 4140
rect 41932 4100 110236 4128
rect 41932 4088 41938 4100
rect 110230 4088 110236 4100
rect 110288 4088 110294 4140
rect 110340 4128 110368 4168
rect 385678 4156 385684 4208
rect 385736 4196 385742 4208
rect 391842 4196 391848 4208
rect 385736 4168 391848 4196
rect 385736 4156 385742 4168
rect 391842 4156 391848 4168
rect 391900 4156 391906 4208
rect 395338 4156 395344 4208
rect 395396 4196 395402 4208
rect 402514 4196 402520 4208
rect 395396 4168 402520 4196
rect 395396 4156 395402 4168
rect 402514 4156 402520 4168
rect 402572 4156 402578 4208
rect 429930 4156 429936 4208
rect 429988 4196 429994 4208
rect 430850 4196 430856 4208
rect 429988 4168 430856 4196
rect 429988 4156 429994 4168
rect 430850 4156 430856 4168
rect 430908 4156 430914 4208
rect 431954 4156 431960 4208
rect 432012 4196 432018 4208
rect 433242 4196 433248 4208
rect 432012 4168 433248 4196
rect 432012 4156 432018 4168
rect 433242 4156 433248 4168
rect 433300 4156 433306 4208
rect 457530 4156 457536 4208
rect 457588 4196 457594 4208
rect 459186 4196 459192 4208
rect 457588 4168 459192 4196
rect 457588 4156 457594 4168
rect 459186 4156 459192 4168
rect 459244 4156 459250 4208
rect 461578 4156 461584 4208
rect 461636 4196 461642 4208
rect 462774 4196 462780 4208
rect 461636 4168 462780 4196
rect 461636 4156 461642 4168
rect 462774 4156 462780 4168
rect 462832 4156 462838 4208
rect 468478 4156 468484 4208
rect 468536 4196 468542 4208
rect 469858 4196 469864 4208
rect 468536 4168 469864 4196
rect 468536 4156 468542 4168
rect 469858 4156 469864 4168
rect 469916 4156 469922 4208
rect 471238 4156 471244 4208
rect 471296 4196 471302 4208
rect 473446 4196 473452 4208
rect 471296 4168 473452 4196
rect 471296 4156 471302 4168
rect 473446 4156 473452 4168
rect 473504 4156 473510 4208
rect 482278 4156 482284 4208
rect 482336 4196 482342 4208
rect 484026 4196 484032 4208
rect 482336 4168 484032 4196
rect 482336 4156 482342 4168
rect 484026 4156 484032 4168
rect 484084 4156 484090 4208
rect 485038 4156 485044 4208
rect 485096 4196 485102 4208
rect 487614 4196 487620 4208
rect 485096 4168 487620 4196
rect 485096 4156 485102 4168
rect 487614 4156 487620 4168
rect 487672 4156 487678 4208
rect 506474 4156 506480 4208
rect 506532 4196 506538 4208
rect 507670 4196 507676 4208
rect 506532 4168 507676 4196
rect 506532 4156 506538 4168
rect 507670 4156 507676 4168
rect 507728 4156 507734 4208
rect 511350 4156 511356 4208
rect 511408 4196 511414 4208
rect 513558 4196 513564 4208
rect 511408 4168 513564 4196
rect 511408 4156 511414 4168
rect 513558 4156 513564 4168
rect 513616 4156 513622 4208
rect 529198 4156 529204 4208
rect 529256 4196 529262 4208
rect 534902 4196 534908 4208
rect 529256 4168 534908 4196
rect 529256 4156 529262 4168
rect 534902 4156 534908 4168
rect 534960 4156 534966 4208
rect 112806 4128 112812 4140
rect 110340 4100 112812 4128
rect 112806 4088 112812 4100
rect 112864 4088 112870 4140
rect 159358 4128 159364 4140
rect 113146 4100 159364 4128
rect 31294 4020 31300 4072
rect 31352 4060 31358 4072
rect 39390 4060 39396 4072
rect 31352 4032 39396 4060
rect 31352 4020 31358 4032
rect 39390 4020 39396 4032
rect 39448 4020 39454 4072
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 43128 4032 108436 4060
rect 43128 4020 43134 4032
rect 23014 3952 23020 4004
rect 23072 3992 23078 4004
rect 43438 3992 43444 4004
rect 23072 3964 43444 3992
rect 23072 3952 23078 3964
rect 43438 3952 43444 3964
rect 43496 3952 43502 4004
rect 46658 3952 46664 4004
rect 46716 3992 46722 4004
rect 108301 3995 108359 4001
rect 108301 3992 108313 3995
rect 46716 3964 108313 3992
rect 46716 3952 46722 3964
rect 108301 3961 108313 3964
rect 108347 3961 108359 3995
rect 108408 3992 108436 4032
rect 109310 4020 109316 4072
rect 109368 4060 109374 4072
rect 113146 4060 113174 4100
rect 159358 4088 159364 4100
rect 159416 4088 159422 4140
rect 175458 4088 175464 4140
rect 175516 4128 175522 4140
rect 207566 4128 207572 4140
rect 175516 4100 207572 4128
rect 175516 4088 175522 4100
rect 207566 4088 207572 4100
rect 207624 4088 207630 4140
rect 285398 4088 285404 4140
rect 285456 4128 285462 4140
rect 287698 4128 287704 4140
rect 285456 4100 287704 4128
rect 285456 4088 285462 4100
rect 287698 4088 287704 4100
rect 287756 4088 287762 4140
rect 296622 4088 296628 4140
rect 296680 4128 296686 4140
rect 297266 4128 297272 4140
rect 296680 4100 297272 4128
rect 296680 4088 296686 4100
rect 297266 4088 297272 4100
rect 297324 4088 297330 4140
rect 304902 4088 304908 4140
rect 304960 4128 304966 4140
rect 307938 4128 307944 4140
rect 304960 4100 307944 4128
rect 304960 4088 304966 4100
rect 307938 4088 307944 4100
rect 307996 4088 308002 4140
rect 335262 4088 335268 4140
rect 335320 4128 335326 4140
rect 350442 4128 350448 4140
rect 335320 4100 350448 4128
rect 335320 4088 335326 4100
rect 350442 4088 350448 4100
rect 350500 4088 350506 4140
rect 353202 4088 353208 4140
rect 353260 4128 353266 4140
rect 375282 4128 375288 4140
rect 353260 4100 375288 4128
rect 353260 4088 353266 4100
rect 375282 4088 375288 4100
rect 375340 4088 375346 4140
rect 382182 4088 382188 4140
rect 382240 4128 382246 4140
rect 384669 4131 384727 4137
rect 384669 4128 384681 4131
rect 382240 4100 384681 4128
rect 382240 4088 382246 4100
rect 384669 4097 384681 4100
rect 384715 4097 384727 4131
rect 384669 4091 384727 4097
rect 384761 4131 384819 4137
rect 384761 4097 384773 4131
rect 384807 4128 384819 4131
rect 410794 4128 410800 4140
rect 384807 4100 410800 4128
rect 384807 4097 384819 4100
rect 384761 4091 384819 4097
rect 410794 4088 410800 4100
rect 410852 4088 410858 4140
rect 419442 4088 419448 4140
rect 419500 4128 419506 4140
rect 465166 4128 465172 4140
rect 419500 4100 465172 4128
rect 419500 4088 419506 4100
rect 465166 4088 465172 4100
rect 465224 4088 465230 4140
rect 487062 4088 487068 4140
rect 487120 4128 487126 4140
rect 557350 4128 557356 4140
rect 487120 4100 557356 4128
rect 487120 4088 487126 4100
rect 557350 4088 557356 4100
rect 557408 4088 557414 4140
rect 109368 4032 113174 4060
rect 123389 4063 123447 4069
rect 109368 4020 109374 4032
rect 123389 4029 123401 4063
rect 123435 4060 123447 4063
rect 166994 4060 167000 4072
rect 123435 4032 167000 4060
rect 123435 4029 123447 4032
rect 123389 4023 123447 4029
rect 166994 4020 167000 4032
rect 167052 4020 167058 4072
rect 179046 4020 179052 4072
rect 179104 4060 179110 4072
rect 179104 4032 209774 4060
rect 179104 4020 179110 4032
rect 111058 3992 111064 4004
rect 108408 3964 111064 3992
rect 108301 3955 108359 3961
rect 111058 3952 111064 3964
rect 111116 3952 111122 4004
rect 114002 3952 114008 4004
rect 114060 3992 114066 4004
rect 161566 3992 161572 4004
rect 114060 3964 161572 3992
rect 114060 3952 114066 3964
rect 161566 3952 161572 3964
rect 161624 3952 161630 4004
rect 174262 3952 174268 4004
rect 174320 3992 174326 4004
rect 206738 3992 206744 4004
rect 174320 3964 206744 3992
rect 174320 3952 174326 3964
rect 206738 3952 206744 3964
rect 206796 3952 206802 4004
rect 35986 3884 35992 3936
rect 36044 3924 36050 3936
rect 95513 3927 95571 3933
rect 95513 3924 95525 3927
rect 36044 3896 95525 3924
rect 36044 3884 36050 3896
rect 95513 3893 95525 3896
rect 95559 3893 95571 3927
rect 95513 3887 95571 3893
rect 95605 3927 95663 3933
rect 95605 3893 95617 3927
rect 95651 3924 95663 3927
rect 100754 3924 100760 3936
rect 95651 3896 100760 3924
rect 95651 3893 95663 3896
rect 95605 3887 95663 3893
rect 100754 3884 100760 3896
rect 100812 3884 100818 3936
rect 102226 3884 102232 3936
rect 102284 3924 102290 3936
rect 146941 3927 146999 3933
rect 146941 3924 146953 3927
rect 102284 3896 146953 3924
rect 102284 3884 102290 3896
rect 146941 3893 146953 3896
rect 146987 3893 146999 3927
rect 146941 3887 146999 3893
rect 147033 3927 147091 3933
rect 147033 3893 147045 3927
rect 147079 3924 147091 3927
rect 149882 3924 149888 3936
rect 147079 3896 149888 3924
rect 147079 3893 147091 3896
rect 147033 3887 147091 3893
rect 149882 3884 149888 3896
rect 149940 3884 149946 3936
rect 160094 3924 160100 3936
rect 151786 3896 160100 3924
rect 5258 3816 5264 3868
rect 5316 3856 5322 3868
rect 7558 3856 7564 3868
rect 5316 3828 7564 3856
rect 5316 3816 5322 3828
rect 7558 3816 7564 3828
rect 7616 3816 7622 3868
rect 39574 3816 39580 3868
rect 39632 3856 39638 3868
rect 108482 3856 108488 3868
rect 39632 3828 108488 3856
rect 39632 3816 39638 3828
rect 108482 3816 108488 3828
rect 108540 3816 108546 3868
rect 110506 3816 110512 3868
rect 110564 3856 110570 3868
rect 151786 3856 151814 3896
rect 160094 3884 160100 3896
rect 160152 3884 160158 3936
rect 170766 3884 170772 3936
rect 170824 3924 170830 3936
rect 204070 3924 204076 3936
rect 170824 3896 204076 3924
rect 170824 3884 170830 3896
rect 204070 3884 204076 3896
rect 204128 3884 204134 3936
rect 110564 3828 151814 3856
rect 110564 3816 110570 3828
rect 167178 3816 167184 3868
rect 167236 3856 167242 3868
rect 193309 3859 193367 3865
rect 193309 3856 193321 3859
rect 167236 3828 193321 3856
rect 167236 3816 167242 3828
rect 193309 3825 193321 3828
rect 193355 3825 193367 3859
rect 209746 3856 209774 4032
rect 311802 4020 311808 4072
rect 311860 4060 311866 4072
rect 318518 4060 318524 4072
rect 311860 4032 318524 4060
rect 311860 4020 311866 4032
rect 318518 4020 318524 4032
rect 318576 4020 318582 4072
rect 322842 4020 322848 4072
rect 322900 4060 322906 4072
rect 332686 4060 332692 4072
rect 322900 4032 332692 4060
rect 322900 4020 322906 4032
rect 332686 4020 332692 4032
rect 332744 4020 332750 4072
rect 342162 4020 342168 4072
rect 342220 4060 342226 4072
rect 358630 4060 358636 4072
rect 342220 4032 358636 4060
rect 342220 4020 342226 4032
rect 358630 4020 358636 4032
rect 358688 4020 358694 4072
rect 360102 4020 360108 4072
rect 360160 4060 360166 4072
rect 383470 4060 383476 4072
rect 360160 4032 383476 4060
rect 360160 4020 360166 4032
rect 383470 4020 383476 4032
rect 383528 4020 383534 4072
rect 415486 4060 415492 4072
rect 384776 4032 415492 4060
rect 324130 3952 324136 4004
rect 324188 3992 324194 4004
rect 335078 3992 335084 4004
rect 324188 3964 335084 3992
rect 324188 3952 324194 3964
rect 335078 3952 335084 3964
rect 335136 3952 335142 4004
rect 336642 3952 336648 4004
rect 336700 3992 336706 4004
rect 351638 3992 351644 4004
rect 336700 3964 351644 3992
rect 336700 3952 336706 3964
rect 351638 3952 351644 3964
rect 351696 3952 351702 4004
rect 357342 3952 357348 4004
rect 357400 3992 357406 4004
rect 379974 3992 379980 4004
rect 357400 3964 379980 3992
rect 357400 3952 357406 3964
rect 379974 3952 379980 3964
rect 380032 3952 380038 4004
rect 383562 3952 383568 4004
rect 383620 3992 383626 4004
rect 384776 3992 384804 4032
rect 415486 4020 415492 4032
rect 415544 4020 415550 4072
rect 420822 4020 420828 4072
rect 420880 4060 420886 4072
rect 467466 4060 467472 4072
rect 420880 4032 467472 4060
rect 420880 4020 420886 4032
rect 467466 4020 467472 4032
rect 467524 4020 467530 4072
rect 491202 4020 491208 4072
rect 491260 4060 491266 4072
rect 563238 4060 563244 4072
rect 491260 4032 563244 4060
rect 491260 4020 491266 4032
rect 563238 4020 563244 4032
rect 563296 4020 563302 4072
rect 383620 3964 384804 3992
rect 384853 3995 384911 4001
rect 383620 3952 383626 3964
rect 384853 3961 384865 3995
rect 384899 3992 384911 3995
rect 414290 3992 414296 4004
rect 384899 3964 414296 3992
rect 384899 3961 384911 3964
rect 384853 3955 384911 3961
rect 414290 3952 414296 3964
rect 414348 3952 414354 4004
rect 418062 3952 418068 4004
rect 418120 3992 418126 4004
rect 463970 3992 463976 4004
rect 418120 3964 463976 3992
rect 418120 3952 418126 3964
rect 463970 3952 463976 3964
rect 464028 3952 464034 4004
rect 488350 3952 488356 4004
rect 488408 3992 488414 4004
rect 560846 3992 560852 4004
rect 488408 3964 560852 3992
rect 488408 3952 488414 3964
rect 560846 3952 560852 3964
rect 560904 3952 560910 4004
rect 305638 3884 305644 3936
rect 305696 3924 305702 3936
rect 309042 3924 309048 3936
rect 305696 3896 309048 3924
rect 305696 3884 305702 3896
rect 309042 3884 309048 3896
rect 309100 3884 309106 3936
rect 328362 3884 328368 3936
rect 328420 3924 328426 3936
rect 339862 3924 339868 3936
rect 328420 3896 339868 3924
rect 328420 3884 328426 3896
rect 339862 3884 339868 3896
rect 339920 3884 339926 3936
rect 340782 3884 340788 3936
rect 340840 3924 340846 3936
rect 357526 3924 357532 3936
rect 340840 3896 357532 3924
rect 340840 3884 340846 3896
rect 357526 3884 357532 3896
rect 357584 3884 357590 3936
rect 362862 3884 362868 3936
rect 362920 3924 362926 3936
rect 362920 3896 384896 3924
rect 362920 3884 362926 3896
rect 210142 3856 210148 3868
rect 209746 3828 210148 3856
rect 193309 3819 193367 3825
rect 210142 3816 210148 3828
rect 210200 3816 210206 3868
rect 224218 3856 224224 3868
rect 210252 3828 224224 3856
rect 18230 3748 18236 3800
rect 18288 3788 18294 3800
rect 29638 3788 29644 3800
rect 18288 3760 29644 3788
rect 18288 3748 18294 3760
rect 29638 3748 29644 3760
rect 29696 3748 29702 3800
rect 32398 3748 32404 3800
rect 32456 3788 32462 3800
rect 95513 3791 95571 3797
rect 32456 3760 95464 3788
rect 32456 3748 32462 3760
rect 28902 3680 28908 3732
rect 28960 3720 28966 3732
rect 95329 3723 95387 3729
rect 95329 3720 95341 3723
rect 28960 3692 95341 3720
rect 28960 3680 28966 3692
rect 95329 3689 95341 3692
rect 95375 3689 95387 3723
rect 95436 3720 95464 3760
rect 95513 3757 95525 3791
rect 95559 3788 95571 3791
rect 105630 3788 105636 3800
rect 95559 3760 105636 3788
rect 95559 3757 95571 3760
rect 95513 3751 95571 3757
rect 105630 3748 105636 3760
rect 105688 3748 105694 3800
rect 105722 3748 105728 3800
rect 105780 3788 105786 3800
rect 156782 3788 156788 3800
rect 105780 3760 156788 3788
rect 105780 3748 105786 3760
rect 156782 3748 156788 3760
rect 156840 3748 156846 3800
rect 160094 3748 160100 3800
rect 160152 3788 160158 3800
rect 196342 3788 196348 3800
rect 160152 3760 196348 3788
rect 160152 3748 160158 3760
rect 196342 3748 196348 3760
rect 196400 3748 196406 3800
rect 198918 3788 198924 3800
rect 196452 3760 198924 3788
rect 103238 3720 103244 3732
rect 95436 3692 103244 3720
rect 95329 3683 95387 3689
rect 103238 3680 103244 3692
rect 103296 3680 103302 3732
rect 103330 3680 103336 3732
rect 103388 3720 103394 3732
rect 155034 3720 155040 3732
rect 103388 3692 155040 3720
rect 103388 3680 103394 3692
rect 155034 3680 155040 3692
rect 155092 3680 155098 3732
rect 163682 3680 163688 3732
rect 163740 3720 163746 3732
rect 196452 3720 196480 3760
rect 198918 3748 198924 3760
rect 198976 3748 198982 3800
rect 209774 3748 209780 3800
rect 209832 3788 209838 3800
rect 210252 3788 210280 3828
rect 224218 3816 224224 3828
rect 224276 3816 224282 3868
rect 313182 3816 313188 3868
rect 313240 3856 313246 3868
rect 319714 3856 319720 3868
rect 313240 3828 319720 3856
rect 313240 3816 313246 3828
rect 319714 3816 319720 3828
rect 319772 3816 319778 3868
rect 321462 3816 321468 3868
rect 321520 3856 321526 3868
rect 330386 3856 330392 3868
rect 321520 3828 330392 3856
rect 321520 3816 321526 3828
rect 330386 3816 330392 3828
rect 330444 3816 330450 3868
rect 331122 3816 331128 3868
rect 331180 3856 331186 3868
rect 344554 3856 344560 3868
rect 331180 3828 344560 3856
rect 331180 3816 331186 3828
rect 344554 3816 344560 3828
rect 344612 3816 344618 3868
rect 346302 3816 346308 3868
rect 346360 3856 346366 3868
rect 364610 3856 364616 3868
rect 346360 3828 364616 3856
rect 346360 3816 346366 3828
rect 364610 3816 364616 3828
rect 364668 3816 364674 3868
rect 367002 3816 367008 3868
rect 367060 3856 367066 3868
rect 384669 3859 384727 3865
rect 384669 3856 384681 3859
rect 367060 3828 384681 3856
rect 367060 3816 367066 3828
rect 384669 3825 384681 3828
rect 384715 3825 384727 3859
rect 384868 3856 384896 3896
rect 384942 3884 384948 3936
rect 385000 3924 385006 3936
rect 417878 3924 417884 3936
rect 385000 3896 417884 3924
rect 385000 3884 385006 3896
rect 417878 3884 417884 3896
rect 417936 3884 417942 3936
rect 424870 3884 424876 3936
rect 424928 3924 424934 3936
rect 472250 3924 472256 3936
rect 424928 3896 472256 3924
rect 424928 3884 424934 3896
rect 472250 3884 472256 3896
rect 472308 3884 472314 3936
rect 492582 3884 492588 3936
rect 492640 3924 492646 3936
rect 566826 3924 566832 3936
rect 492640 3896 566832 3924
rect 492640 3884 492646 3896
rect 566826 3884 566832 3896
rect 566884 3884 566890 3936
rect 387150 3856 387156 3868
rect 384868 3828 387156 3856
rect 384669 3819 384727 3825
rect 387150 3816 387156 3828
rect 387208 3816 387214 3868
rect 387521 3859 387579 3865
rect 387521 3825 387533 3859
rect 387567 3856 387579 3859
rect 390373 3859 390431 3865
rect 390373 3856 390385 3859
rect 387567 3828 390385 3856
rect 387567 3825 387579 3828
rect 387521 3819 387579 3825
rect 390373 3825 390385 3828
rect 390419 3825 390431 3859
rect 390373 3819 390431 3825
rect 390462 3816 390468 3868
rect 390520 3856 390526 3868
rect 424962 3856 424968 3868
rect 390520 3828 424968 3856
rect 390520 3816 390526 3828
rect 424962 3816 424968 3828
rect 425020 3816 425026 3868
rect 426342 3816 426348 3868
rect 426400 3856 426406 3868
rect 474550 3856 474556 3868
rect 426400 3828 474556 3856
rect 426400 3816 426406 3828
rect 474550 3816 474556 3828
rect 474608 3816 474614 3868
rect 493962 3816 493968 3868
rect 494020 3856 494026 3868
rect 568022 3856 568028 3868
rect 494020 3828 568028 3856
rect 494020 3816 494026 3828
rect 568022 3816 568028 3828
rect 568080 3816 568086 3868
rect 209832 3760 210280 3788
rect 214561 3791 214619 3797
rect 209832 3748 209838 3760
rect 214561 3757 214573 3791
rect 214607 3788 214619 3791
rect 230842 3788 230848 3800
rect 214607 3760 230848 3788
rect 214607 3757 214619 3760
rect 214561 3751 214619 3757
rect 230842 3748 230848 3760
rect 230900 3748 230906 3800
rect 327718 3748 327724 3800
rect 327776 3788 327782 3800
rect 338666 3788 338672 3800
rect 327776 3760 338672 3788
rect 327776 3748 327782 3760
rect 338666 3748 338672 3760
rect 338724 3748 338730 3800
rect 339402 3748 339408 3800
rect 339460 3788 339466 3800
rect 355226 3788 355232 3800
rect 339460 3760 355232 3788
rect 339460 3748 339466 3760
rect 355226 3748 355232 3760
rect 355284 3748 355290 3800
rect 355962 3748 355968 3800
rect 356020 3788 356026 3800
rect 378870 3788 378876 3800
rect 356020 3760 378876 3788
rect 356020 3748 356026 3760
rect 378870 3748 378876 3760
rect 378928 3748 378934 3800
rect 379422 3748 379428 3800
rect 379480 3788 379486 3800
rect 384761 3791 384819 3797
rect 384761 3788 384773 3791
rect 379480 3760 384773 3788
rect 379480 3748 379486 3760
rect 384761 3757 384773 3760
rect 384807 3757 384819 3791
rect 384761 3751 384819 3757
rect 384850 3748 384856 3800
rect 384908 3788 384914 3800
rect 418982 3788 418988 3800
rect 384908 3760 418988 3788
rect 384908 3748 384914 3760
rect 418982 3748 418988 3760
rect 419040 3748 419046 3800
rect 423582 3748 423588 3800
rect 423640 3788 423646 3800
rect 471054 3788 471060 3800
rect 423640 3760 471060 3788
rect 423640 3748 423646 3760
rect 471054 3748 471060 3760
rect 471112 3748 471118 3800
rect 491110 3748 491116 3800
rect 491168 3788 491174 3800
rect 564434 3788 564440 3800
rect 491168 3760 564440 3788
rect 491168 3748 491174 3760
rect 564434 3748 564440 3760
rect 564492 3748 564498 3800
rect 163740 3692 196480 3720
rect 163740 3680 163746 3692
rect 196802 3680 196808 3732
rect 196860 3720 196866 3732
rect 196860 3692 200114 3720
rect 196860 3680 196866 3692
rect 24210 3612 24216 3664
rect 24268 3652 24274 3664
rect 97350 3652 97356 3664
rect 24268 3624 97356 3652
rect 24268 3612 24274 3624
rect 97350 3612 97356 3624
rect 97408 3612 97414 3664
rect 97442 3612 97448 3664
rect 97500 3652 97506 3664
rect 97902 3652 97908 3664
rect 97500 3624 97908 3652
rect 97500 3612 97506 3624
rect 97902 3612 97908 3624
rect 97960 3612 97966 3664
rect 98638 3612 98644 3664
rect 98696 3652 98702 3664
rect 151538 3652 151544 3664
rect 98696 3624 151544 3652
rect 98696 3612 98702 3624
rect 151538 3612 151544 3624
rect 151596 3612 151602 3664
rect 156598 3612 156604 3664
rect 156656 3652 156662 3664
rect 193766 3652 193772 3664
rect 156656 3624 193772 3652
rect 156656 3612 156662 3624
rect 193766 3612 193772 3624
rect 193824 3612 193830 3664
rect 195606 3612 195612 3664
rect 195664 3652 195670 3664
rect 199378 3652 199384 3664
rect 195664 3624 199384 3652
rect 195664 3612 195670 3624
rect 199378 3612 199384 3624
rect 199436 3612 199442 3664
rect 200086 3652 200114 3692
rect 200298 3680 200304 3732
rect 200356 3720 200362 3732
rect 225690 3720 225696 3732
rect 200356 3692 225696 3720
rect 200356 3680 200362 3692
rect 225690 3680 225696 3692
rect 225748 3680 225754 3732
rect 314562 3680 314568 3732
rect 314620 3720 314626 3732
rect 320910 3720 320916 3732
rect 314620 3692 320916 3720
rect 314620 3680 314626 3692
rect 320910 3680 320916 3692
rect 320968 3680 320974 3732
rect 321002 3680 321008 3732
rect 321060 3720 321066 3732
rect 329190 3720 329196 3732
rect 321060 3692 329196 3720
rect 321060 3680 321066 3692
rect 329190 3680 329196 3692
rect 329248 3680 329254 3732
rect 329742 3680 329748 3732
rect 329800 3720 329806 3732
rect 329800 3692 342024 3720
rect 329800 3680 329806 3692
rect 223022 3652 223028 3664
rect 200086 3624 223028 3652
rect 223022 3612 223028 3624
rect 223080 3612 223086 3664
rect 318610 3612 318616 3664
rect 318668 3652 318674 3664
rect 324593 3655 324651 3661
rect 324593 3652 324605 3655
rect 318668 3624 324605 3652
rect 318668 3612 318674 3624
rect 324593 3621 324605 3624
rect 324639 3621 324651 3655
rect 324593 3615 324651 3621
rect 325510 3612 325516 3664
rect 325568 3652 325574 3664
rect 337470 3652 337476 3664
rect 325568 3624 337476 3652
rect 325568 3612 325574 3624
rect 337470 3612 337476 3624
rect 337528 3612 337534 3664
rect 339310 3612 339316 3664
rect 339368 3652 339374 3664
rect 341996 3652 342024 3692
rect 342070 3680 342076 3732
rect 342128 3720 342134 3732
rect 359918 3720 359924 3732
rect 342128 3692 359924 3720
rect 342128 3680 342134 3692
rect 359918 3680 359924 3692
rect 359976 3680 359982 3732
rect 361482 3680 361488 3732
rect 361540 3720 361546 3732
rect 385954 3720 385960 3732
rect 361540 3692 385960 3720
rect 361540 3680 361546 3692
rect 385954 3680 385960 3692
rect 386012 3680 386018 3732
rect 387702 3680 387708 3732
rect 387760 3720 387766 3732
rect 394881 3723 394939 3729
rect 387760 3692 394832 3720
rect 387760 3680 387766 3692
rect 342162 3652 342168 3664
rect 339368 3624 341196 3652
rect 341996 3624 342168 3652
rect 339368 3612 339374 3624
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 98178 3584 98184 3596
rect 25372 3556 98184 3584
rect 25372 3544 25378 3556
rect 98178 3544 98184 3556
rect 98236 3544 98242 3596
rect 99834 3544 99840 3596
rect 99892 3584 99898 3596
rect 146849 3587 146907 3593
rect 146849 3584 146861 3587
rect 99892 3556 146861 3584
rect 99892 3544 99898 3556
rect 146849 3553 146861 3556
rect 146895 3553 146907 3587
rect 146849 3547 146907 3553
rect 146941 3587 146999 3593
rect 146941 3553 146953 3587
rect 146987 3584 146999 3587
rect 154114 3584 154120 3596
rect 146987 3556 154120 3584
rect 146987 3553 146999 3556
rect 146941 3547 146999 3553
rect 154114 3544 154120 3556
rect 154172 3544 154178 3596
rect 155402 3544 155408 3596
rect 155460 3584 155466 3596
rect 193309 3587 193367 3593
rect 155460 3556 185624 3584
rect 155460 3544 155466 3556
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 18598 3516 18604 3528
rect 17092 3488 18604 3516
rect 17092 3476 17098 3488
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 19484 3488 85620 3516
rect 19484 3476 19490 3488
rect 9950 3408 9956 3460
rect 10008 3448 10014 3460
rect 85485 3451 85543 3457
rect 85485 3448 85497 3451
rect 10008 3420 85497 3448
rect 10008 3408 10014 3420
rect 85485 3417 85497 3420
rect 85531 3417 85543 3451
rect 85592 3448 85620 3488
rect 85666 3476 85672 3528
rect 85724 3516 85730 3528
rect 86678 3516 86684 3528
rect 85724 3488 86684 3516
rect 85724 3476 85730 3488
rect 86678 3476 86684 3488
rect 86736 3476 86742 3528
rect 90269 3519 90327 3525
rect 90269 3516 90281 3519
rect 86788 3488 90281 3516
rect 86788 3448 86816 3488
rect 90269 3485 90281 3488
rect 90315 3485 90327 3519
rect 90269 3479 90327 3485
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 96246 3476 96252 3528
rect 96304 3516 96310 3528
rect 147033 3519 147091 3525
rect 147033 3516 147045 3519
rect 96304 3488 147045 3516
rect 96304 3476 96310 3488
rect 147033 3485 147045 3488
rect 147079 3485 147091 3519
rect 147033 3479 147091 3485
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 153102 3516 153108 3528
rect 151872 3488 153108 3516
rect 151872 3476 151878 3488
rect 153102 3476 153108 3488
rect 153160 3476 153166 3528
rect 158898 3476 158904 3528
rect 158956 3516 158962 3528
rect 160002 3516 160008 3528
rect 158956 3488 160008 3516
rect 158956 3476 158962 3488
rect 160002 3476 160008 3488
rect 160060 3476 160066 3528
rect 166074 3476 166080 3528
rect 166132 3516 166138 3528
rect 166902 3516 166908 3528
rect 166132 3488 166908 3516
rect 166132 3476 166138 3488
rect 166902 3476 166908 3488
rect 166960 3476 166966 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173802 3516 173808 3528
rect 173216 3488 173808 3516
rect 173216 3476 173222 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177942 3516 177948 3528
rect 176712 3488 177948 3516
rect 176712 3476 176718 3488
rect 177942 3476 177948 3488
rect 178000 3476 178006 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180702 3516 180708 3528
rect 180300 3488 180708 3516
rect 180300 3476 180306 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 85592 3420 86816 3448
rect 85485 3411 85543 3417
rect 89162 3408 89168 3460
rect 89220 3448 89226 3460
rect 134061 3451 134119 3457
rect 134061 3448 134073 3451
rect 89220 3420 134073 3448
rect 89220 3408 89226 3420
rect 134061 3417 134073 3420
rect 134107 3417 134119 3451
rect 134061 3411 134119 3417
rect 134150 3408 134156 3460
rect 134208 3448 134214 3460
rect 135162 3448 135168 3460
rect 134208 3420 135168 3448
rect 134208 3408 134214 3420
rect 135162 3408 135168 3420
rect 135220 3408 135226 3460
rect 141234 3408 141240 3460
rect 141292 3448 141298 3460
rect 142062 3448 142068 3460
rect 141292 3420 142068 3448
rect 141292 3408 141298 3420
rect 142062 3408 142068 3420
rect 142120 3408 142126 3460
rect 145926 3408 145932 3460
rect 145984 3448 145990 3460
rect 145984 3420 181392 3448
rect 145984 3408 145990 3420
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 17218 3380 17224 3392
rect 11204 3352 17224 3380
rect 11204 3340 11210 3352
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 35250 3380 35256 3392
rect 33652 3352 35256 3380
rect 33652 3340 33658 3352
rect 35250 3340 35256 3352
rect 35308 3340 35314 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 45462 3340 45468 3392
rect 45520 3380 45526 3392
rect 106829 3383 106887 3389
rect 106829 3380 106841 3383
rect 45520 3352 106841 3380
rect 45520 3340 45526 3352
rect 106829 3349 106841 3352
rect 106875 3349 106887 3383
rect 106829 3343 106887 3349
rect 106918 3340 106924 3392
rect 106976 3380 106982 3392
rect 107562 3380 107568 3392
rect 106976 3352 107568 3380
rect 106976 3340 106982 3352
rect 107562 3340 107568 3352
rect 107620 3340 107626 3392
rect 108301 3383 108359 3389
rect 108301 3349 108313 3383
rect 108347 3380 108359 3383
rect 113726 3380 113732 3392
rect 108347 3352 113732 3380
rect 108347 3349 108359 3352
rect 108301 3343 108359 3349
rect 113726 3340 113732 3352
rect 113784 3340 113790 3392
rect 116394 3340 116400 3392
rect 116452 3380 116458 3392
rect 117222 3380 117228 3392
rect 116452 3352 117228 3380
rect 116452 3340 116458 3352
rect 117222 3340 117228 3352
rect 117280 3340 117286 3392
rect 121086 3340 121092 3392
rect 121144 3380 121150 3392
rect 167914 3380 167920 3392
rect 121144 3352 167920 3380
rect 121144 3340 121150 3352
rect 167914 3340 167920 3352
rect 167972 3340 167978 3392
rect 52546 3272 52552 3324
rect 52604 3312 52610 3324
rect 53742 3312 53748 3324
rect 52604 3284 53748 3312
rect 52604 3272 52610 3284
rect 53742 3272 53748 3284
rect 53800 3272 53806 3324
rect 53837 3315 53895 3321
rect 53837 3281 53849 3315
rect 53883 3312 53895 3315
rect 116302 3312 116308 3324
rect 53883 3284 116308 3312
rect 53883 3281 53895 3284
rect 53837 3275 53895 3281
rect 116302 3272 116308 3284
rect 116360 3272 116366 3324
rect 117590 3272 117596 3324
rect 117648 3312 117654 3324
rect 165338 3312 165344 3324
rect 117648 3284 165344 3312
rect 117648 3272 117654 3284
rect 165338 3272 165344 3284
rect 165396 3272 165402 3324
rect 8754 3204 8760 3256
rect 8812 3244 8818 3256
rect 11698 3244 11704 3256
rect 8812 3216 11704 3244
rect 8812 3204 8818 3216
rect 11698 3204 11704 3216
rect 11756 3204 11762 3256
rect 38378 3204 38384 3256
rect 38436 3244 38442 3256
rect 50430 3244 50436 3256
rect 38436 3216 50436 3244
rect 38436 3204 38442 3216
rect 50430 3204 50436 3216
rect 50488 3204 50494 3256
rect 118878 3244 118884 3256
rect 53760 3216 118884 3244
rect 53760 3188 53788 3216
rect 118878 3204 118884 3216
rect 118936 3204 118942 3256
rect 119890 3204 119896 3256
rect 119948 3244 119954 3256
rect 123389 3247 123447 3253
rect 123389 3244 123401 3247
rect 119948 3216 123401 3244
rect 119948 3204 119954 3216
rect 123389 3213 123401 3216
rect 123435 3213 123447 3247
rect 123389 3207 123447 3213
rect 123478 3204 123484 3256
rect 123536 3244 123542 3256
rect 124122 3244 124128 3256
rect 123536 3216 124128 3244
rect 123536 3204 123542 3216
rect 124122 3204 124128 3216
rect 124180 3204 124186 3256
rect 124674 3204 124680 3256
rect 124732 3244 124738 3256
rect 125502 3244 125508 3256
rect 124732 3216 125508 3244
rect 124732 3204 124738 3216
rect 125502 3204 125508 3216
rect 125560 3204 125566 3256
rect 134061 3247 134119 3253
rect 134061 3213 134073 3247
rect 134107 3244 134119 3247
rect 144638 3244 144644 3256
rect 134107 3216 144644 3244
rect 134107 3213 134119 3216
rect 134061 3207 134119 3213
rect 144638 3204 144644 3216
rect 144696 3204 144702 3256
rect 146849 3247 146907 3253
rect 146849 3213 146861 3247
rect 146895 3244 146907 3247
rect 152458 3244 152464 3256
rect 146895 3216 152464 3244
rect 146895 3213 146907 3216
rect 146849 3207 146907 3213
rect 152458 3204 152464 3216
rect 152516 3204 152522 3256
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 15838 3176 15844 3188
rect 13596 3148 15844 3176
rect 13596 3136 13602 3148
rect 15838 3136 15844 3148
rect 15896 3136 15902 3188
rect 53742 3136 53748 3188
rect 53800 3136 53806 3188
rect 57238 3136 57244 3188
rect 57296 3176 57302 3188
rect 121638 3176 121644 3188
rect 57296 3148 121644 3176
rect 57296 3136 57302 3148
rect 121638 3136 121644 3148
rect 121696 3136 121702 3188
rect 149514 3136 149520 3188
rect 149572 3176 149578 3188
rect 181364 3176 181392 3420
rect 183738 3408 183744 3460
rect 183796 3448 183802 3460
rect 184842 3448 184848 3460
rect 183796 3420 184848 3448
rect 183796 3408 183802 3420
rect 184842 3408 184848 3420
rect 184900 3408 184906 3460
rect 185596 3448 185624 3556
rect 193309 3553 193321 3587
rect 193355 3584 193367 3587
rect 201586 3584 201592 3596
rect 193355 3556 201592 3584
rect 193355 3553 193367 3556
rect 193309 3547 193367 3553
rect 201586 3544 201592 3556
rect 201644 3544 201650 3596
rect 207382 3544 207388 3596
rect 207440 3584 207446 3596
rect 214561 3587 214619 3593
rect 214561 3584 214573 3587
rect 207440 3556 214573 3584
rect 207440 3544 207446 3556
rect 214561 3553 214573 3556
rect 214607 3553 214619 3587
rect 214561 3547 214619 3553
rect 221550 3544 221556 3596
rect 221608 3584 221614 3596
rect 228358 3584 228364 3596
rect 221608 3556 228364 3584
rect 221608 3544 221614 3556
rect 228358 3544 228364 3556
rect 228416 3544 228422 3596
rect 247586 3544 247592 3596
rect 247644 3584 247650 3596
rect 251818 3584 251824 3596
rect 247644 3556 251824 3584
rect 247644 3544 247650 3556
rect 251818 3544 251824 3556
rect 251876 3544 251882 3596
rect 267734 3544 267740 3596
rect 267792 3584 267798 3596
rect 268930 3584 268936 3596
rect 267792 3556 268936 3584
rect 267792 3544 267798 3556
rect 268930 3544 268936 3556
rect 268988 3544 268994 3596
rect 318702 3544 318708 3596
rect 318760 3584 318766 3596
rect 326798 3584 326804 3596
rect 318760 3556 326804 3584
rect 318760 3544 318766 3556
rect 326798 3544 326804 3556
rect 326856 3544 326862 3596
rect 328270 3544 328276 3596
rect 328328 3584 328334 3596
rect 340966 3584 340972 3596
rect 328328 3556 340972 3584
rect 328328 3544 328334 3556
rect 340966 3544 340972 3556
rect 341024 3544 341030 3596
rect 341168 3584 341196 3624
rect 342162 3612 342168 3624
rect 342220 3612 342226 3664
rect 356330 3652 356336 3664
rect 342272 3624 356336 3652
rect 342272 3584 342300 3624
rect 356330 3612 356336 3624
rect 356388 3612 356394 3664
rect 358722 3612 358728 3664
rect 358780 3652 358786 3664
rect 382366 3652 382372 3664
rect 358780 3624 382372 3652
rect 358780 3612 358786 3624
rect 382366 3612 382372 3624
rect 382424 3612 382430 3664
rect 384669 3655 384727 3661
rect 384669 3621 384681 3655
rect 384715 3652 384727 3655
rect 387521 3655 387579 3661
rect 387521 3652 387533 3655
rect 384715 3624 387533 3652
rect 384715 3621 384727 3624
rect 384669 3615 384727 3621
rect 387521 3621 387533 3624
rect 387567 3621 387579 3655
rect 387521 3615 387579 3621
rect 387610 3612 387616 3664
rect 387668 3652 387674 3664
rect 394697 3655 394755 3661
rect 394697 3652 394709 3655
rect 387668 3624 394709 3652
rect 387668 3612 387674 3624
rect 394697 3621 394709 3624
rect 394743 3621 394755 3655
rect 394804 3652 394832 3692
rect 394881 3689 394893 3723
rect 394927 3720 394939 3723
rect 421374 3720 421380 3732
rect 394927 3692 421380 3720
rect 394927 3689 394939 3692
rect 394881 3683 394939 3689
rect 421374 3680 421380 3692
rect 421432 3680 421438 3732
rect 429102 3680 429108 3732
rect 429160 3720 429166 3732
rect 478138 3720 478144 3732
rect 429160 3692 478144 3720
rect 429160 3680 429166 3692
rect 478138 3680 478144 3692
rect 478196 3680 478202 3732
rect 495342 3680 495348 3732
rect 495400 3720 495406 3732
rect 570322 3720 570328 3732
rect 495400 3692 570328 3720
rect 495400 3680 495406 3692
rect 570322 3680 570328 3692
rect 570380 3680 570386 3732
rect 422570 3652 422576 3664
rect 394804 3624 422576 3652
rect 394697 3615 394755 3621
rect 422570 3612 422576 3624
rect 422628 3612 422634 3664
rect 426250 3612 426256 3664
rect 426308 3652 426314 3664
rect 475746 3652 475752 3664
rect 426308 3624 475752 3652
rect 426308 3612 426314 3624
rect 475746 3612 475752 3624
rect 475804 3612 475810 3664
rect 499482 3612 499488 3664
rect 499540 3652 499546 3664
rect 575106 3652 575112 3664
rect 499540 3624 575112 3652
rect 499540 3612 499546 3624
rect 575106 3612 575112 3624
rect 575164 3612 575170 3664
rect 341168 3556 342300 3584
rect 344830 3544 344836 3596
rect 344888 3584 344894 3596
rect 363506 3584 363512 3596
rect 344888 3556 363512 3584
rect 344888 3544 344894 3556
rect 363506 3544 363512 3556
rect 363564 3544 363570 3596
rect 364242 3544 364248 3596
rect 364300 3584 364306 3596
rect 389450 3584 389456 3596
rect 364300 3556 389456 3584
rect 364300 3544 364306 3556
rect 389450 3544 389456 3556
rect 389508 3544 389514 3596
rect 390373 3587 390431 3593
rect 390373 3553 390385 3587
rect 390419 3584 390431 3587
rect 393038 3584 393044 3596
rect 390419 3556 393044 3584
rect 390419 3553 390431 3556
rect 390373 3547 390431 3553
rect 393038 3544 393044 3556
rect 393096 3544 393102 3596
rect 393222 3544 393228 3596
rect 393280 3584 393286 3596
rect 429654 3584 429660 3596
rect 393280 3556 429660 3584
rect 393280 3544 393286 3556
rect 429654 3544 429660 3556
rect 429712 3544 429718 3596
rect 431862 3544 431868 3596
rect 431920 3584 431926 3596
rect 482830 3584 482836 3596
rect 431920 3556 482836 3584
rect 431920 3544 431926 3556
rect 482830 3544 482836 3556
rect 482888 3544 482894 3596
rect 496722 3544 496728 3596
rect 496780 3584 496786 3596
rect 571518 3584 571524 3596
rect 496780 3556 571524 3584
rect 496780 3544 496786 3556
rect 571518 3544 571524 3556
rect 571576 3544 571582 3596
rect 188522 3476 188528 3528
rect 188580 3516 188586 3528
rect 188580 3488 200114 3516
rect 188580 3476 188586 3488
rect 192938 3448 192944 3460
rect 185596 3420 192944 3448
rect 192938 3408 192944 3420
rect 192996 3408 193002 3460
rect 194410 3408 194416 3460
rect 194468 3448 194474 3460
rect 195238 3448 195244 3460
rect 194468 3420 195244 3448
rect 194468 3408 194474 3420
rect 195238 3408 195244 3420
rect 195296 3408 195302 3460
rect 197906 3408 197912 3460
rect 197964 3448 197970 3460
rect 198642 3448 198648 3460
rect 197964 3420 198648 3448
rect 197964 3408 197970 3420
rect 198642 3408 198648 3420
rect 198700 3408 198706 3460
rect 200086 3448 200114 3488
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 202782 3516 202788 3528
rect 201552 3488 202788 3516
rect 201552 3476 201558 3488
rect 202782 3476 202788 3488
rect 202840 3476 202846 3528
rect 203886 3476 203892 3528
rect 203944 3516 203950 3528
rect 204898 3516 204904 3528
rect 203944 3488 204904 3516
rect 203944 3476 203950 3488
rect 204898 3476 204904 3488
rect 204956 3476 204962 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 205542 3516 205548 3528
rect 205140 3488 205548 3516
rect 205140 3476 205146 3488
rect 205542 3476 205548 3488
rect 205600 3476 205606 3528
rect 206186 3476 206192 3528
rect 206244 3516 206250 3528
rect 206922 3516 206928 3528
rect 206244 3488 206928 3516
rect 206244 3476 206250 3488
rect 206922 3476 206928 3488
rect 206980 3476 206986 3528
rect 208578 3476 208584 3528
rect 208636 3516 208642 3528
rect 209682 3516 209688 3528
rect 208636 3488 209688 3516
rect 208636 3476 208642 3488
rect 209682 3476 209688 3488
rect 209740 3476 209746 3528
rect 212166 3476 212172 3528
rect 212224 3516 212230 3528
rect 213178 3516 213184 3528
rect 212224 3488 213184 3516
rect 212224 3476 212230 3488
rect 213178 3476 213184 3488
rect 213236 3476 213242 3528
rect 213362 3476 213368 3528
rect 213420 3516 213426 3528
rect 213822 3516 213828 3528
rect 213420 3488 213828 3516
rect 213420 3476 213426 3488
rect 213822 3476 213828 3488
rect 213880 3476 213886 3528
rect 214466 3476 214472 3528
rect 214524 3516 214530 3528
rect 215202 3516 215208 3528
rect 214524 3488 215208 3516
rect 214524 3476 214530 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 216582 3516 216588 3528
rect 215720 3488 216588 3516
rect 215720 3476 215726 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 216858 3476 216864 3528
rect 216916 3516 216922 3528
rect 217962 3516 217968 3528
rect 216916 3488 217968 3516
rect 216916 3476 216922 3488
rect 217962 3476 217968 3488
rect 218020 3476 218026 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 219342 3516 219348 3528
rect 218112 3488 219348 3516
rect 218112 3476 218118 3488
rect 219342 3476 219348 3488
rect 219400 3476 219406 3528
rect 222746 3476 222752 3528
rect 222804 3516 222810 3528
rect 223482 3516 223488 3528
rect 222804 3488 223488 3516
rect 222804 3476 222810 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 225138 3476 225144 3528
rect 225196 3516 225202 3528
rect 226242 3516 226248 3528
rect 225196 3488 226248 3516
rect 225196 3476 225202 3488
rect 226242 3476 226248 3488
rect 226300 3476 226306 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 227622 3516 227628 3528
rect 226392 3488 227628 3516
rect 226392 3476 226398 3488
rect 227622 3476 227628 3488
rect 227680 3476 227686 3528
rect 231026 3476 231032 3528
rect 231084 3516 231090 3528
rect 231762 3516 231768 3528
rect 231084 3488 231768 3516
rect 231084 3476 231090 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 238110 3476 238116 3528
rect 238168 3516 238174 3528
rect 238662 3516 238668 3528
rect 238168 3488 238668 3516
rect 238168 3476 238174 3488
rect 238662 3476 238668 3488
rect 238720 3476 238726 3528
rect 240502 3476 240508 3528
rect 240560 3516 240566 3528
rect 241422 3516 241428 3528
rect 240560 3488 241428 3516
rect 240560 3476 240566 3488
rect 241422 3476 241428 3488
rect 241480 3476 241486 3528
rect 248782 3476 248788 3528
rect 248840 3516 248846 3528
rect 249702 3516 249708 3528
rect 248840 3488 249708 3516
rect 248840 3476 248846 3488
rect 249702 3476 249708 3488
rect 249760 3476 249766 3528
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 251082 3516 251088 3528
rect 250036 3488 251088 3516
rect 250036 3476 250042 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 251174 3476 251180 3528
rect 251232 3516 251238 3528
rect 252462 3516 252468 3528
rect 251232 3488 252468 3516
rect 251232 3476 251238 3488
rect 252462 3476 252468 3488
rect 252520 3476 252526 3528
rect 254670 3476 254676 3528
rect 254728 3516 254734 3528
rect 255222 3516 255228 3528
rect 254728 3488 255228 3516
rect 254728 3476 254734 3488
rect 255222 3476 255228 3488
rect 255280 3476 255286 3528
rect 255866 3476 255872 3528
rect 255924 3516 255930 3528
rect 256602 3516 256608 3528
rect 255924 3488 256608 3516
rect 255924 3476 255930 3488
rect 256602 3476 256608 3488
rect 256660 3476 256666 3528
rect 258258 3476 258264 3528
rect 258316 3516 258322 3528
rect 259362 3516 259368 3528
rect 258316 3488 259368 3516
rect 258316 3476 258322 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 259454 3476 259460 3528
rect 259512 3516 259518 3528
rect 260742 3516 260748 3528
rect 259512 3488 260748 3516
rect 259512 3476 259518 3488
rect 260742 3476 260748 3488
rect 260800 3476 260806 3528
rect 262950 3476 262956 3528
rect 263008 3516 263014 3528
rect 263502 3516 263508 3528
rect 263008 3488 263508 3516
rect 263008 3476 263014 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 264882 3516 264888 3528
rect 264204 3488 264888 3516
rect 264204 3476 264210 3488
rect 264882 3476 264888 3488
rect 264940 3476 264946 3528
rect 266538 3476 266544 3528
rect 266596 3516 266602 3528
rect 267642 3516 267648 3528
rect 266596 3488 267648 3516
rect 266596 3476 266602 3488
rect 267642 3476 267648 3488
rect 267700 3476 267706 3528
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 274542 3516 274548 3528
rect 273680 3488 274548 3516
rect 273680 3476 273686 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 279510 3476 279516 3528
rect 279568 3516 279574 3528
rect 280798 3516 280804 3528
rect 279568 3488 280804 3516
rect 279568 3476 279574 3488
rect 280798 3476 280804 3488
rect 280856 3476 280862 3528
rect 288986 3476 288992 3528
rect 289044 3516 289050 3528
rect 289722 3516 289728 3528
rect 289044 3488 289728 3516
rect 289044 3476 289050 3488
rect 289722 3476 289728 3488
rect 289780 3476 289786 3528
rect 291378 3476 291384 3528
rect 291436 3516 291442 3528
rect 291930 3516 291936 3528
rect 291436 3488 291936 3516
rect 291436 3476 291442 3488
rect 291930 3476 291936 3488
rect 291988 3476 291994 3528
rect 292574 3476 292580 3528
rect 292632 3516 292638 3528
rect 293678 3516 293684 3528
rect 292632 3488 293684 3516
rect 292632 3476 292638 3488
rect 293678 3476 293684 3488
rect 293736 3476 293742 3528
rect 295334 3476 295340 3528
rect 295392 3516 295398 3528
rect 296070 3516 296076 3528
rect 295392 3488 296076 3516
rect 295392 3476 295398 3488
rect 296070 3476 296076 3488
rect 296128 3476 296134 3528
rect 298738 3476 298744 3528
rect 298796 3516 298802 3528
rect 299658 3516 299664 3528
rect 298796 3488 299664 3516
rect 298796 3476 298802 3488
rect 299658 3476 299664 3488
rect 299716 3476 299722 3528
rect 300762 3476 300768 3528
rect 300820 3516 300826 3528
rect 301958 3516 301964 3528
rect 300820 3488 301964 3516
rect 300820 3476 300826 3488
rect 301958 3476 301964 3488
rect 302016 3476 302022 3528
rect 310330 3476 310336 3528
rect 310388 3516 310394 3528
rect 315022 3516 315028 3528
rect 310388 3488 315028 3516
rect 310388 3476 310394 3488
rect 315022 3476 315028 3488
rect 315080 3476 315086 3528
rect 321370 3476 321376 3528
rect 321428 3516 321434 3528
rect 324593 3519 324651 3525
rect 321428 3488 324544 3516
rect 321428 3476 321434 3488
rect 217042 3448 217048 3460
rect 200086 3420 217048 3448
rect 217042 3408 217048 3420
rect 217100 3408 217106 3460
rect 231118 3448 231124 3460
rect 219406 3420 231124 3448
rect 181438 3340 181444 3392
rect 181496 3380 181502 3392
rect 211890 3380 211896 3392
rect 181496 3352 211896 3380
rect 181496 3340 181502 3352
rect 211890 3340 211896 3352
rect 211948 3340 211954 3392
rect 219250 3340 219256 3392
rect 219308 3380 219314 3392
rect 219406 3380 219434 3420
rect 231118 3408 231124 3420
rect 231176 3408 231182 3460
rect 244090 3408 244096 3460
rect 244148 3448 244154 3460
rect 251910 3448 251916 3460
rect 244148 3420 251916 3448
rect 244148 3408 244154 3420
rect 251910 3408 251916 3420
rect 251968 3408 251974 3460
rect 257062 3408 257068 3460
rect 257120 3448 257126 3460
rect 264238 3448 264244 3460
rect 257120 3420 264244 3448
rect 257120 3408 257126 3420
rect 264238 3408 264244 3420
rect 264296 3408 264302 3460
rect 272426 3408 272432 3460
rect 272484 3448 272490 3460
rect 273898 3448 273904 3460
rect 272484 3420 273904 3448
rect 272484 3408 272490 3420
rect 273898 3408 273904 3420
rect 273956 3408 273962 3460
rect 276014 3408 276020 3460
rect 276072 3448 276078 3460
rect 280154 3448 280160 3460
rect 276072 3420 280160 3448
rect 276072 3408 276078 3420
rect 280154 3408 280160 3420
rect 280212 3408 280218 3460
rect 280706 3408 280712 3460
rect 280764 3448 280770 3460
rect 282178 3448 282184 3460
rect 280764 3420 282184 3448
rect 280764 3408 280770 3420
rect 282178 3408 282184 3420
rect 282236 3408 282242 3460
rect 307570 3408 307576 3460
rect 307628 3448 307634 3460
rect 312630 3448 312636 3460
rect 307628 3420 312636 3448
rect 307628 3408 307634 3420
rect 312630 3408 312636 3420
rect 312688 3408 312694 3460
rect 317322 3408 317328 3460
rect 317380 3448 317386 3460
rect 324406 3448 324412 3460
rect 317380 3420 324412 3448
rect 317380 3408 317386 3420
rect 324406 3408 324412 3420
rect 324464 3408 324470 3460
rect 324516 3448 324544 3488
rect 324593 3485 324605 3519
rect 324639 3516 324651 3519
rect 327994 3516 328000 3528
rect 324639 3488 328000 3516
rect 324639 3485 324651 3488
rect 324593 3479 324651 3485
rect 327994 3476 328000 3488
rect 328052 3476 328058 3528
rect 332410 3476 332416 3528
rect 332468 3516 332474 3528
rect 345750 3516 345756 3528
rect 332468 3488 345756 3516
rect 332468 3476 332474 3488
rect 345750 3476 345756 3488
rect 345808 3476 345814 3528
rect 346210 3476 346216 3528
rect 346268 3516 346274 3528
rect 365806 3516 365812 3528
rect 346268 3488 365812 3516
rect 346268 3476 346274 3488
rect 365806 3476 365812 3488
rect 365864 3476 365870 3528
rect 369670 3476 369676 3528
rect 369728 3516 369734 3528
rect 397730 3516 397736 3528
rect 369728 3488 397736 3516
rect 369728 3476 369734 3488
rect 397730 3476 397736 3488
rect 397788 3476 397794 3528
rect 398742 3476 398748 3528
rect 398800 3516 398806 3528
rect 436738 3516 436744 3528
rect 398800 3488 436744 3516
rect 398800 3476 398806 3488
rect 436738 3476 436744 3488
rect 436796 3476 436802 3528
rect 437382 3476 437388 3528
rect 437440 3516 437446 3528
rect 489914 3516 489920 3528
rect 437440 3488 489920 3516
rect 437440 3476 437446 3488
rect 489914 3476 489920 3488
rect 489972 3476 489978 3528
rect 498010 3476 498016 3528
rect 498068 3516 498074 3528
rect 573910 3516 573916 3528
rect 498068 3488 573916 3516
rect 498068 3476 498074 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 331582 3448 331588 3460
rect 324516 3420 331588 3448
rect 331582 3408 331588 3420
rect 331640 3408 331646 3460
rect 335170 3408 335176 3460
rect 335228 3448 335234 3460
rect 349246 3448 349252 3460
rect 335228 3420 349252 3448
rect 335228 3408 335234 3420
rect 349246 3408 349252 3420
rect 349304 3408 349310 3460
rect 351822 3408 351828 3460
rect 351880 3448 351886 3460
rect 372890 3448 372896 3460
rect 351880 3420 372896 3448
rect 351880 3408 351886 3420
rect 372890 3408 372896 3420
rect 372948 3408 372954 3460
rect 373902 3408 373908 3460
rect 373960 3448 373966 3460
rect 403618 3448 403624 3460
rect 373960 3420 403624 3448
rect 373960 3408 373966 3420
rect 403618 3408 403624 3420
rect 403676 3408 403682 3460
rect 404262 3408 404268 3460
rect 404320 3448 404326 3460
rect 443822 3448 443828 3460
rect 404320 3420 443828 3448
rect 404320 3408 404326 3420
rect 443822 3408 443828 3420
rect 443880 3408 443886 3460
rect 447042 3408 447048 3460
rect 447100 3448 447106 3460
rect 504174 3448 504180 3460
rect 447100 3420 504180 3448
rect 447100 3408 447106 3420
rect 504174 3408 504180 3420
rect 504232 3408 504238 3460
rect 505002 3408 505008 3460
rect 505060 3448 505066 3460
rect 583386 3448 583392 3460
rect 505060 3420 583392 3448
rect 505060 3408 505066 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 219308 3352 219434 3380
rect 219308 3340 219314 3352
rect 332502 3340 332508 3392
rect 332560 3380 332566 3392
rect 346946 3380 346952 3392
rect 332560 3352 346952 3380
rect 332560 3340 332566 3352
rect 346946 3340 346952 3352
rect 347004 3340 347010 3392
rect 349062 3340 349068 3392
rect 349120 3380 349126 3392
rect 352929 3383 352987 3389
rect 352929 3380 352941 3383
rect 349120 3352 352941 3380
rect 349120 3340 349126 3352
rect 352929 3349 352941 3352
rect 352975 3349 352987 3383
rect 352929 3343 352987 3349
rect 354582 3340 354588 3392
rect 354640 3380 354646 3392
rect 376478 3380 376484 3392
rect 354640 3352 376484 3380
rect 354640 3340 354646 3352
rect 376478 3340 376484 3352
rect 376536 3340 376542 3392
rect 376662 3340 376668 3392
rect 376720 3380 376726 3392
rect 407206 3380 407212 3392
rect 376720 3352 407212 3380
rect 376720 3340 376726 3352
rect 407206 3340 407212 3352
rect 407264 3340 407270 3392
rect 422202 3340 422208 3392
rect 422260 3380 422266 3392
rect 468662 3380 468668 3392
rect 422260 3352 468668 3380
rect 422260 3340 422266 3352
rect 468662 3340 468668 3352
rect 468720 3340 468726 3392
rect 484210 3340 484216 3392
rect 484268 3380 484274 3392
rect 553762 3380 553768 3392
rect 484268 3352 553768 3380
rect 484268 3340 484274 3352
rect 553762 3340 553768 3352
rect 553820 3340 553826 3392
rect 182542 3272 182548 3324
rect 182600 3312 182606 3324
rect 212718 3312 212724 3324
rect 182600 3284 212724 3312
rect 182600 3272 182606 3284
rect 212718 3272 212724 3284
rect 212776 3272 212782 3324
rect 229830 3272 229836 3324
rect 229888 3312 229894 3324
rect 233878 3312 233884 3324
rect 229888 3284 233884 3312
rect 229888 3272 229894 3284
rect 233878 3272 233884 3284
rect 233936 3272 233942 3324
rect 234614 3272 234620 3324
rect 234672 3312 234678 3324
rect 238018 3312 238024 3324
rect 234672 3284 238024 3312
rect 234672 3272 234678 3284
rect 238018 3272 238024 3284
rect 238076 3272 238082 3324
rect 246390 3272 246396 3324
rect 246448 3312 246454 3324
rect 246942 3312 246948 3324
rect 246448 3284 246948 3312
rect 246448 3272 246454 3284
rect 246942 3272 246948 3284
rect 247000 3272 247006 3324
rect 249058 3312 249064 3324
rect 248386 3284 249064 3312
rect 184934 3204 184940 3256
rect 184992 3244 184998 3256
rect 214374 3244 214380 3256
rect 184992 3216 214380 3244
rect 184992 3204 184998 3216
rect 214374 3204 214380 3216
rect 214432 3204 214438 3256
rect 223942 3204 223948 3256
rect 224000 3244 224006 3256
rect 224862 3244 224868 3256
rect 224000 3216 224868 3244
rect 224000 3204 224006 3216
rect 224862 3204 224868 3216
rect 224920 3204 224926 3256
rect 241698 3204 241704 3256
rect 241756 3244 241762 3256
rect 242802 3244 242808 3256
rect 241756 3216 242808 3244
rect 241756 3204 241762 3216
rect 242802 3204 242808 3216
rect 242860 3204 242866 3256
rect 242894 3204 242900 3256
rect 242952 3244 242958 3256
rect 248386 3244 248414 3284
rect 249058 3272 249064 3284
rect 249116 3272 249122 3324
rect 252370 3272 252376 3324
rect 252428 3312 252434 3324
rect 255958 3312 255964 3324
rect 252428 3284 255964 3312
rect 252428 3272 252434 3284
rect 255958 3272 255964 3284
rect 256016 3272 256022 3324
rect 271230 3272 271236 3324
rect 271288 3312 271294 3324
rect 271782 3312 271788 3324
rect 271288 3284 271788 3312
rect 271288 3272 271294 3284
rect 271782 3272 271788 3284
rect 271840 3272 271846 3324
rect 287790 3272 287796 3324
rect 287848 3312 287854 3324
rect 288342 3312 288348 3324
rect 287848 3284 288348 3312
rect 287848 3272 287854 3284
rect 288342 3272 288348 3284
rect 288400 3272 288406 3324
rect 307662 3272 307668 3324
rect 307720 3312 307726 3324
rect 311434 3312 311440 3324
rect 307720 3284 311440 3312
rect 307720 3272 307726 3284
rect 311434 3272 311440 3284
rect 311492 3272 311498 3324
rect 325602 3272 325608 3324
rect 325660 3312 325666 3324
rect 336274 3312 336280 3324
rect 325660 3284 336280 3312
rect 325660 3272 325666 3284
rect 336274 3272 336280 3284
rect 336332 3272 336338 3324
rect 348050 3312 348056 3324
rect 340846 3284 348056 3312
rect 242952 3216 248414 3244
rect 242952 3204 242958 3216
rect 324222 3204 324228 3256
rect 324280 3244 324286 3256
rect 333882 3244 333888 3256
rect 324280 3216 333888 3244
rect 324280 3204 324286 3216
rect 333882 3204 333888 3216
rect 333940 3204 333946 3256
rect 186038 3176 186044 3188
rect 149572 3148 180794 3176
rect 181364 3148 186044 3176
rect 149572 3136 149578 3148
rect 34790 3068 34796 3120
rect 34848 3108 34854 3120
rect 34848 3080 45554 3108
rect 34848 3068 34854 3080
rect 45526 3040 45554 3080
rect 50154 3068 50160 3120
rect 50212 3108 50218 3120
rect 53837 3111 53895 3117
rect 53837 3108 53849 3111
rect 50212 3080 53849 3108
rect 50212 3068 50218 3080
rect 53837 3077 53849 3080
rect 53883 3077 53895 3111
rect 53837 3071 53895 3077
rect 64322 3068 64328 3120
rect 64380 3108 64386 3120
rect 126606 3108 126612 3120
rect 64380 3080 126612 3108
rect 64380 3068 64386 3080
rect 126606 3068 126612 3080
rect 126664 3068 126670 3120
rect 180766 3108 180794 3148
rect 186038 3136 186044 3148
rect 186096 3136 186102 3188
rect 189718 3136 189724 3188
rect 189776 3176 189782 3188
rect 217870 3176 217876 3188
rect 189776 3148 217876 3176
rect 189776 3136 189782 3148
rect 217870 3136 217876 3148
rect 217928 3136 217934 3188
rect 265342 3136 265348 3188
rect 265400 3176 265406 3188
rect 269758 3176 269764 3188
rect 265400 3148 269764 3176
rect 265400 3136 265406 3148
rect 269758 3136 269764 3148
rect 269816 3136 269822 3188
rect 284294 3136 284300 3188
rect 284352 3176 284358 3188
rect 286778 3176 286784 3188
rect 284352 3148 286784 3176
rect 284352 3136 284358 3148
rect 286778 3136 286784 3148
rect 286836 3136 286842 3188
rect 311710 3136 311716 3188
rect 311768 3176 311774 3188
rect 317322 3176 317328 3188
rect 311768 3148 317328 3176
rect 311768 3136 311774 3148
rect 317322 3136 317328 3148
rect 317380 3136 317386 3188
rect 340846 3176 340874 3284
rect 348050 3272 348056 3284
rect 348108 3272 348114 3324
rect 351730 3272 351736 3324
rect 351788 3312 351794 3324
rect 356149 3315 356207 3321
rect 351788 3284 356100 3312
rect 351788 3272 351794 3284
rect 352834 3244 352840 3256
rect 336752 3148 340874 3176
rect 344986 3216 352840 3244
rect 188614 3108 188620 3120
rect 180766 3080 188620 3108
rect 188614 3068 188620 3080
rect 188672 3068 188678 3120
rect 193214 3068 193220 3120
rect 193272 3108 193278 3120
rect 213733 3111 213791 3117
rect 213733 3108 213745 3111
rect 193272 3080 213745 3108
rect 193272 3068 193278 3080
rect 213733 3077 213745 3080
rect 213779 3077 213791 3111
rect 213733 3071 213791 3077
rect 239306 3068 239312 3120
rect 239364 3108 239370 3120
rect 246298 3108 246304 3120
rect 239364 3080 246304 3108
rect 239364 3068 239370 3080
rect 246298 3068 246304 3080
rect 246356 3068 246362 3120
rect 281902 3068 281908 3120
rect 281960 3108 281966 3120
rect 285030 3108 285036 3120
rect 281960 3080 285036 3108
rect 281960 3068 281966 3080
rect 285030 3068 285036 3080
rect 285088 3068 285094 3120
rect 336090 3068 336096 3120
rect 336148 3108 336154 3120
rect 336752 3108 336780 3148
rect 336148 3080 336780 3108
rect 336148 3068 336154 3080
rect 338758 3068 338764 3120
rect 338816 3108 338822 3120
rect 344986 3108 345014 3216
rect 352834 3204 352840 3216
rect 352892 3204 352898 3256
rect 352929 3247 352987 3253
rect 352929 3213 352941 3247
rect 352975 3244 352987 3247
rect 355965 3247 356023 3253
rect 355965 3244 355977 3247
rect 352975 3216 355977 3244
rect 352975 3213 352987 3216
rect 352929 3207 352987 3213
rect 355965 3213 355977 3216
rect 356011 3213 356023 3247
rect 356072 3244 356100 3284
rect 356149 3281 356161 3315
rect 356195 3312 356207 3315
rect 369394 3312 369400 3324
rect 356195 3284 369400 3312
rect 356195 3281 356207 3284
rect 356149 3275 356207 3281
rect 369394 3272 369400 3284
rect 369452 3272 369458 3324
rect 380802 3272 380808 3324
rect 380860 3312 380866 3324
rect 411898 3312 411904 3324
rect 380860 3284 411904 3312
rect 380860 3272 380866 3284
rect 411898 3272 411904 3284
rect 411956 3272 411962 3324
rect 415302 3272 415308 3324
rect 415360 3312 415366 3324
rect 460382 3312 460388 3324
rect 415360 3284 460388 3312
rect 415360 3272 415366 3284
rect 460382 3272 460388 3284
rect 460440 3272 460446 3324
rect 481542 3272 481548 3324
rect 481600 3312 481606 3324
rect 481600 3284 543044 3312
rect 481600 3272 481606 3284
rect 371694 3244 371700 3256
rect 356072 3216 371700 3244
rect 355965 3207 356023 3213
rect 371694 3204 371700 3216
rect 371752 3204 371758 3256
rect 375190 3204 375196 3256
rect 375248 3244 375254 3256
rect 404814 3244 404820 3256
rect 375248 3216 404820 3244
rect 375248 3204 375254 3216
rect 404814 3204 404820 3216
rect 404872 3204 404878 3256
rect 416590 3204 416596 3256
rect 416648 3244 416654 3256
rect 461578 3244 461584 3256
rect 416648 3216 461584 3244
rect 416648 3204 416654 3216
rect 461578 3204 461584 3216
rect 461636 3204 461642 3256
rect 478782 3204 478788 3256
rect 478840 3244 478846 3256
rect 542817 3247 542875 3253
rect 542817 3244 542829 3247
rect 478840 3216 542829 3244
rect 478840 3204 478846 3216
rect 542817 3213 542829 3216
rect 542863 3213 542875 3247
rect 542817 3207 542875 3213
rect 350350 3136 350356 3188
rect 350408 3176 350414 3188
rect 370590 3176 370596 3188
rect 350408 3148 370596 3176
rect 350408 3136 350414 3148
rect 370590 3136 370596 3148
rect 370648 3136 370654 3188
rect 378042 3136 378048 3188
rect 378100 3176 378106 3188
rect 408402 3176 408408 3188
rect 378100 3148 408408 3176
rect 378100 3136 378106 3148
rect 408402 3136 408408 3148
rect 408460 3136 408466 3188
rect 412542 3136 412548 3188
rect 412600 3176 412606 3188
rect 456886 3176 456892 3188
rect 412600 3148 456892 3176
rect 412600 3136 412606 3148
rect 456886 3136 456892 3148
rect 456944 3136 456950 3188
rect 476022 3136 476028 3188
rect 476080 3176 476086 3188
rect 543016 3176 543044 3284
rect 544378 3272 544384 3324
rect 544436 3312 544442 3324
rect 545482 3312 545488 3324
rect 544436 3284 545488 3312
rect 544436 3272 544442 3284
rect 545482 3272 545488 3284
rect 545540 3272 545546 3324
rect 547138 3204 547144 3256
rect 547196 3244 547202 3256
rect 559742 3244 559748 3256
rect 547196 3216 559748 3244
rect 547196 3204 547202 3216
rect 559742 3204 559748 3216
rect 559800 3204 559806 3256
rect 550266 3176 550272 3188
rect 476080 3148 538214 3176
rect 543016 3148 550272 3176
rect 476080 3136 476086 3148
rect 338816 3080 345014 3108
rect 338816 3068 338822 3080
rect 348970 3068 348976 3120
rect 349028 3108 349034 3120
rect 355873 3111 355931 3117
rect 355873 3108 355885 3111
rect 349028 3080 355885 3108
rect 349028 3068 349034 3080
rect 355873 3077 355885 3080
rect 355919 3077 355931 3111
rect 355873 3071 355931 3077
rect 355965 3111 356023 3117
rect 355965 3077 355977 3111
rect 356011 3108 356023 3111
rect 368198 3108 368204 3120
rect 356011 3080 368204 3108
rect 356011 3077 356023 3080
rect 355965 3071 356023 3077
rect 368198 3068 368204 3080
rect 368256 3068 368262 3120
rect 372522 3068 372528 3120
rect 372580 3108 372586 3120
rect 401318 3108 401324 3120
rect 372580 3080 401324 3108
rect 372580 3068 372586 3080
rect 401318 3068 401324 3080
rect 401376 3068 401382 3120
rect 411070 3068 411076 3120
rect 411128 3108 411134 3120
rect 454494 3108 454500 3120
rect 411128 3080 454500 3108
rect 411128 3068 411134 3080
rect 454494 3068 454500 3080
rect 454552 3068 454558 3120
rect 470502 3068 470508 3120
rect 470560 3108 470566 3120
rect 536098 3108 536104 3120
rect 470560 3080 536104 3108
rect 470560 3068 470566 3080
rect 536098 3068 536104 3080
rect 536156 3068 536162 3120
rect 538186 3108 538214 3148
rect 550266 3136 550272 3148
rect 550324 3136 550330 3188
rect 543182 3108 543188 3120
rect 538186 3080 543188 3108
rect 543182 3068 543188 3080
rect 543240 3068 543246 3120
rect 57146 3040 57152 3052
rect 45526 3012 57152 3040
rect 57146 3000 57152 3012
rect 57204 3000 57210 3052
rect 60826 3000 60832 3052
rect 60884 3040 60890 3052
rect 124030 3040 124036 3052
rect 60884 3012 124036 3040
rect 60884 3000 60890 3012
rect 124030 3000 124036 3012
rect 124088 3000 124094 3052
rect 190822 3000 190828 3052
rect 190880 3040 190886 3052
rect 191742 3040 191748 3052
rect 190880 3012 191748 3040
rect 190880 3000 190886 3012
rect 191742 3000 191748 3012
rect 191800 3000 191806 3052
rect 199102 3000 199108 3052
rect 199160 3040 199166 3052
rect 220078 3040 220084 3052
rect 199160 3012 220084 3040
rect 199160 3000 199166 3012
rect 220078 3000 220084 3012
rect 220136 3000 220142 3052
rect 261754 3000 261760 3052
rect 261812 3040 261818 3052
rect 266998 3040 267004 3052
rect 261812 3012 267004 3040
rect 261812 3000 261818 3012
rect 266998 3000 267004 3012
rect 267056 3000 267062 3052
rect 274818 3000 274824 3052
rect 274876 3040 274882 3052
rect 276658 3040 276664 3052
rect 274876 3012 276664 3040
rect 274876 3000 274882 3012
rect 276658 3000 276664 3012
rect 276716 3000 276722 3052
rect 283098 3000 283104 3052
rect 283156 3040 283162 3052
rect 284938 3040 284944 3052
rect 283156 3012 284944 3040
rect 283156 3000 283162 3012
rect 284938 3000 284944 3012
rect 284996 3000 285002 3052
rect 310422 3000 310428 3052
rect 310480 3040 310486 3052
rect 316218 3040 316224 3052
rect 310480 3012 316224 3040
rect 310480 3000 310486 3012
rect 316218 3000 316224 3012
rect 316276 3000 316282 3052
rect 316678 3000 316684 3052
rect 316736 3040 316742 3052
rect 323302 3040 323308 3052
rect 316736 3012 323308 3040
rect 316736 3000 316742 3012
rect 323302 3000 323308 3012
rect 323360 3000 323366 3052
rect 335998 3000 336004 3052
rect 336056 3040 336062 3052
rect 343358 3040 343364 3052
rect 336056 3012 343364 3040
rect 336056 3000 336062 3012
rect 343358 3000 343364 3012
rect 343416 3000 343422 3052
rect 347682 3000 347688 3052
rect 347740 3040 347746 3052
rect 367002 3040 367008 3052
rect 347740 3012 367008 3040
rect 347740 3000 347746 3012
rect 367002 3000 367008 3012
rect 367060 3000 367066 3052
rect 394234 3040 394240 3052
rect 367112 3012 394240 3040
rect 27706 2932 27712 2984
rect 27764 2972 27770 2984
rect 35158 2972 35164 2984
rect 27764 2944 35164 2972
rect 27764 2932 27770 2944
rect 35158 2932 35164 2944
rect 35216 2932 35222 2984
rect 73798 2932 73804 2984
rect 73856 2972 73862 2984
rect 74442 2972 74448 2984
rect 73856 2944 74448 2972
rect 73856 2932 73862 2944
rect 74442 2932 74448 2944
rect 74500 2932 74506 2984
rect 76190 2932 76196 2984
rect 76248 2972 76254 2984
rect 77202 2972 77208 2984
rect 76248 2944 77208 2972
rect 76248 2932 76254 2944
rect 77202 2932 77208 2944
rect 77260 2932 77266 2984
rect 129182 2972 129188 2984
rect 77496 2944 129188 2972
rect 67910 2864 67916 2916
rect 67968 2904 67974 2916
rect 77496 2904 77524 2944
rect 129182 2932 129188 2944
rect 129240 2932 129246 2984
rect 213733 2975 213791 2981
rect 213733 2941 213745 2975
rect 213779 2972 213791 2975
rect 220446 2972 220452 2984
rect 213779 2944 220452 2972
rect 213779 2941 213791 2944
rect 213733 2935 213791 2941
rect 220446 2932 220452 2944
rect 220504 2932 220510 2984
rect 343542 2932 343548 2984
rect 343600 2972 343606 2984
rect 361114 2972 361120 2984
rect 343600 2944 361120 2972
rect 343600 2932 343606 2944
rect 361114 2932 361120 2944
rect 361172 2932 361178 2984
rect 366910 2932 366916 2984
rect 366968 2972 366974 2984
rect 367112 2972 367140 3012
rect 394234 3000 394240 3012
rect 394292 3000 394298 3052
rect 413922 3000 413928 3052
rect 413980 3040 413986 3052
rect 458082 3040 458088 3052
rect 413980 3012 458088 3040
rect 413980 3000 413986 3012
rect 458082 3000 458088 3012
rect 458140 3000 458146 3052
rect 466362 3000 466368 3052
rect 466420 3040 466426 3052
rect 529014 3040 529020 3052
rect 466420 3012 529020 3040
rect 466420 3000 466426 3012
rect 529014 3000 529020 3012
rect 529072 3000 529078 3052
rect 542817 3043 542875 3049
rect 542817 3009 542829 3043
rect 542863 3040 542875 3043
rect 546678 3040 546684 3052
rect 542863 3012 546684 3040
rect 542863 3009 542875 3012
rect 542817 3003 542875 3009
rect 546678 3000 546684 3012
rect 546736 3000 546742 3052
rect 366968 2944 367140 2972
rect 366968 2932 366974 2944
rect 372430 2932 372436 2984
rect 372488 2972 372494 2984
rect 400122 2972 400128 2984
rect 372488 2944 400128 2972
rect 372488 2932 372494 2944
rect 400122 2932 400128 2944
rect 400180 2932 400186 2984
rect 405642 2932 405648 2984
rect 405700 2972 405706 2984
rect 447410 2972 447416 2984
rect 405700 2944 447416 2972
rect 405700 2932 405706 2944
rect 447410 2932 447416 2944
rect 447468 2932 447474 2984
rect 460842 2932 460848 2984
rect 460900 2972 460906 2984
rect 521838 2972 521844 2984
rect 460900 2944 521844 2972
rect 460900 2932 460906 2944
rect 521838 2932 521844 2944
rect 521896 2932 521902 2984
rect 134334 2904 134340 2916
rect 67968 2876 77524 2904
rect 77588 2876 134340 2904
rect 67968 2864 67974 2876
rect 74994 2796 75000 2848
rect 75052 2836 75058 2848
rect 77588 2836 77616 2876
rect 134334 2864 134340 2876
rect 134392 2864 134398 2916
rect 192018 2864 192024 2916
rect 192076 2904 192082 2916
rect 219618 2904 219624 2916
rect 192076 2876 219624 2904
rect 192076 2864 192082 2876
rect 219618 2864 219624 2876
rect 219676 2864 219682 2916
rect 344922 2864 344928 2916
rect 344980 2904 344986 2916
rect 362310 2904 362316 2916
rect 344980 2876 362316 2904
rect 344980 2864 344986 2876
rect 362310 2864 362316 2876
rect 362368 2864 362374 2916
rect 369762 2864 369768 2916
rect 369820 2904 369826 2916
rect 396534 2904 396540 2916
rect 369820 2876 396540 2904
rect 369820 2864 369826 2876
rect 396534 2864 396540 2876
rect 396592 2864 396598 2916
rect 411162 2864 411168 2916
rect 411220 2904 411226 2916
rect 453298 2904 453304 2916
rect 411220 2876 453304 2904
rect 411220 2864 411226 2876
rect 453298 2864 453304 2876
rect 453356 2864 453362 2916
rect 455322 2864 455328 2916
rect 455380 2904 455386 2916
rect 514754 2904 514760 2916
rect 455380 2876 514760 2904
rect 455380 2864 455386 2876
rect 514754 2864 514760 2876
rect 514812 2864 514818 2916
rect 75052 2808 77616 2836
rect 75052 2796 75058 2808
rect 80882 2796 80888 2848
rect 80940 2836 80946 2848
rect 81342 2836 81348 2848
rect 80940 2808 81348 2836
rect 80940 2796 80946 2808
rect 81342 2796 81348 2808
rect 81400 2796 81406 2848
rect 82078 2796 82084 2848
rect 82136 2836 82142 2848
rect 139486 2836 139492 2848
rect 82136 2808 139492 2836
rect 82136 2796 82142 2808
rect 139486 2796 139492 2808
rect 139544 2796 139550 2848
rect 186130 2796 186136 2848
rect 186188 2836 186194 2848
rect 215386 2836 215392 2848
rect 186188 2808 215392 2836
rect 186188 2796 186194 2808
rect 215386 2796 215392 2808
rect 215444 2796 215450 2848
rect 340138 2796 340144 2848
rect 340196 2836 340202 2848
rect 354030 2836 354036 2848
rect 340196 2808 354036 2836
rect 340196 2796 340202 2808
rect 354030 2796 354036 2808
rect 354088 2796 354094 2848
rect 365622 2796 365628 2848
rect 365680 2836 365686 2848
rect 390646 2836 390652 2848
rect 365680 2808 390652 2836
rect 365680 2796 365686 2808
rect 390646 2796 390652 2808
rect 390704 2796 390710 2848
rect 408310 2796 408316 2848
rect 408368 2836 408374 2848
rect 450906 2836 450912 2848
rect 408368 2808 450912 2836
rect 408368 2796 408374 2808
rect 450906 2796 450912 2808
rect 450964 2796 450970 2848
rect 452562 2796 452568 2848
rect 452620 2836 452626 2848
rect 511258 2836 511264 2848
rect 452620 2808 511264 2836
rect 452620 2796 452626 2808
rect 511258 2796 511264 2808
rect 511316 2796 511322 2848
rect 448514 2320 448520 2372
rect 448572 2360 448578 2372
rect 449802 2360 449808 2372
rect 448572 2332 449808 2360
rect 448572 2320 448578 2332
rect 449802 2320 449808 2332
rect 449860 2320 449866 2372
<< via1 >>
rect 154120 700952 154172 701004
rect 322940 700952 322992 701004
rect 137836 700884 137888 700936
rect 318800 700884 318852 700936
rect 264888 700816 264940 700868
rect 462320 700816 462372 700868
rect 269028 700748 269080 700800
rect 478512 700748 478564 700800
rect 89168 700680 89220 700732
rect 333980 700680 334032 700732
rect 72976 700612 73028 700664
rect 329840 700612 329892 700664
rect 253848 700544 253900 700596
rect 527180 700544 527232 700596
rect 256608 700476 256660 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 338120 700408 338172 700460
rect 24308 700340 24360 700392
rect 345020 700340 345072 700392
rect 8116 700272 8168 700324
rect 342260 700272 342312 700324
rect 280068 700204 280120 700256
rect 413652 700204 413704 700256
rect 275928 700136 275980 700188
rect 397460 700136 397512 700188
rect 202788 700068 202840 700120
rect 307760 700068 307812 700120
rect 218980 700000 219032 700052
rect 311900 700000 311952 700052
rect 291108 699932 291160 699984
rect 348792 699932 348844 699984
rect 286968 699864 287020 699916
rect 332508 699864 332560 699916
rect 267648 699796 267700 699848
rect 296720 699796 296772 699848
rect 283840 699728 283892 699780
rect 300860 699728 300912 699780
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 242808 696940 242860 696992
rect 580172 696940 580224 696992
rect 245568 683204 245620 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 349160 683136 349212 683188
rect 238668 670760 238720 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 356060 670692 356112 670744
rect 3424 656888 3476 656940
rect 353300 656888 353352 656940
rect 231768 643084 231820 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 360200 632068 360252 632120
rect 234528 630640 234580 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 367100 618264 367152 618316
rect 227628 616836 227680 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 364432 605820 364484 605872
rect 219348 590656 219400 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 371240 579640 371292 579692
rect 223488 576852 223540 576904
rect 580172 576852 580224 576904
rect 175096 569032 175148 569084
rect 556804 569032 556856 569084
rect 152740 568964 152792 569016
rect 547144 568964 547196 569016
rect 130384 568896 130436 568948
rect 543004 568896 543056 568948
rect 7564 568828 7616 568880
rect 423956 568828 424008 568880
rect 119160 568760 119212 568812
rect 540244 568760 540296 568812
rect 111708 568692 111760 568744
rect 560944 568692 560996 568744
rect 100576 568624 100628 568676
rect 558184 568624 558236 568676
rect 14464 568556 14516 568608
rect 502432 568556 502484 568608
rect 227168 568488 227220 568540
rect 227628 568488 227680 568540
rect 230940 568488 230992 568540
rect 231768 568488 231820 568540
rect 242072 568488 242124 568540
rect 242808 568488 242860 568540
rect 253296 568488 253348 568540
rect 253848 568488 253900 568540
rect 264428 568488 264480 568540
rect 264888 568488 264940 568540
rect 268200 568488 268252 568540
rect 269028 568488 269080 568540
rect 279332 568488 279384 568540
rect 280068 568488 280120 568540
rect 290556 568488 290608 568540
rect 291108 568488 291160 568540
rect 293868 568488 293920 568540
rect 299480 568488 299532 568540
rect 235908 568420 235960 568472
rect 305000 568420 305052 568472
rect 282828 568352 282880 568404
rect 364340 568352 364392 568404
rect 171048 568284 171100 568336
rect 316040 568284 316092 568336
rect 271788 568216 271840 568268
rect 429200 568216 429252 568268
rect 106188 568148 106240 568200
rect 327080 568148 327132 568200
rect 260564 568080 260616 568132
rect 494060 568080 494112 568132
rect 249524 568012 249576 568064
rect 558920 568012 558972 568064
rect 61384 567944 61436 567996
rect 386696 567944 386748 567996
rect 189908 567876 189960 567928
rect 525064 567876 525116 567928
rect 178776 567808 178828 567860
rect 522304 567808 522356 567860
rect 57244 567740 57296 567792
rect 409052 567740 409104 567792
rect 167644 567672 167696 567724
rect 520924 567672 520976 567724
rect 156420 567604 156472 567656
rect 519544 567604 519596 567656
rect 145288 567536 145340 567588
rect 518164 567536 518216 567588
rect 51724 567468 51776 567520
rect 431408 567468 431460 567520
rect 133788 567400 133840 567452
rect 515404 567400 515456 567452
rect 4896 567332 4948 567384
rect 446312 567332 446364 567384
rect 17224 567264 17276 567316
rect 468668 567264 468720 567316
rect 4804 567196 4856 567248
rect 457444 567196 457496 567248
rect 204812 567060 204864 567112
rect 507124 567060 507176 567112
rect 193680 566992 193732 567044
rect 505744 566992 505796 567044
rect 79324 566924 79376 566976
rect 405280 566924 405332 566976
rect 65524 566856 65576 566908
rect 394148 566856 394200 566908
rect 43444 566788 43496 566840
rect 383016 566788 383068 566840
rect 75184 566720 75236 566772
rect 416780 566720 416832 566772
rect 53104 566652 53156 566704
rect 397920 566652 397972 566704
rect 197268 566584 197320 566636
rect 548524 566584 548576 566636
rect 76564 566516 76616 566568
rect 438860 566516 438912 566568
rect 170956 566448 171008 566500
rect 533344 566448 533396 566500
rect 54484 566380 54536 566432
rect 420184 566380 420236 566432
rect 3424 566312 3476 566364
rect 379520 566312 379572 566364
rect 68284 566244 68336 566296
rect 461216 566244 461268 566296
rect 126612 566176 126664 566228
rect 526444 566176 526496 566228
rect 148968 566108 149020 566160
rect 551284 566108 551336 566160
rect 104256 566040 104308 566092
rect 508504 566040 508556 566092
rect 58624 565972 58676 566024
rect 472348 565972 472400 566024
rect 32404 565904 32456 565956
rect 454040 565904 454092 565956
rect 50344 565836 50396 565888
rect 494704 565836 494756 565888
rect 71044 565632 71096 565684
rect 375564 565632 375616 565684
rect 208216 565564 208268 565616
rect 537484 565564 537536 565616
rect 77944 565496 77996 565548
rect 427958 565496 428010 565548
rect 182226 565428 182278 565480
rect 536104 565428 536156 565480
rect 211942 565360 211994 565412
rect 580448 565360 580500 565412
rect 160008 565292 160060 565344
rect 530584 565292 530636 565344
rect 72424 565224 72476 565276
rect 449992 565224 450044 565276
rect 201132 565156 201184 565208
rect 580356 565156 580408 565208
rect 3792 565088 3844 565140
rect 390560 565088 390612 565140
rect 137836 565020 137888 565072
rect 529204 565020 529256 565072
rect 47584 564952 47636 565004
rect 442540 564952 442592 565004
rect 186228 564884 186280 564936
rect 580264 564884 580316 564936
rect 115480 564816 115532 564868
rect 511264 564816 511316 564868
rect 3700 564748 3752 564800
rect 401600 564748 401652 564800
rect 3608 564680 3660 564732
rect 412824 564680 412876 564732
rect 435088 564723 435140 564732
rect 435088 564689 435097 564723
rect 435097 564689 435131 564723
rect 435131 564689 435140 564723
rect 435088 564680 435140 564689
rect 69664 564612 69716 564664
rect 483572 564612 483624 564664
rect 108028 564544 108080 564596
rect 491208 564544 491260 564596
rect 538864 564544 538916 564596
rect 3516 564476 3568 564528
rect 3424 564408 3476 564460
rect 3332 554684 3384 554736
rect 71044 554684 71096 554736
rect 537484 538160 537536 538212
rect 580172 538160 580224 538212
rect 3240 528504 3292 528556
rect 43444 528504 43496 528556
rect 507124 511912 507176 511964
rect 580172 511912 580224 511964
rect 3240 502256 3292 502308
rect 61384 502256 61436 502308
rect 548524 485732 548576 485784
rect 580172 485732 580224 485784
rect 3332 476008 3384 476060
rect 65524 476008 65576 476060
rect 505744 458124 505796 458176
rect 580172 458124 580224 458176
rect 3332 449828 3384 449880
rect 53104 449828 53156 449880
rect 3332 423580 3384 423632
rect 79324 423580 79376 423632
rect 525064 419432 525116 419484
rect 580172 419432 580224 419484
rect 536104 405628 536156 405680
rect 580172 405628 580224 405680
rect 3332 398760 3384 398812
rect 57244 398760 57296 398812
rect 556804 379448 556856 379500
rect 580172 379448 580224 379500
rect 3332 372512 3384 372564
rect 75184 372512 75236 372564
rect 522304 365644 522356 365696
rect 580172 365644 580224 365696
rect 3148 358572 3200 358624
rect 7564 358572 7616 358624
rect 533344 353200 533396 353252
rect 580172 353200 580224 353252
rect 3332 346332 3384 346384
rect 54484 346332 54536 346384
rect 555424 325592 555476 325644
rect 580172 325592 580224 325644
rect 3332 320084 3384 320136
rect 77944 320084 77996 320136
rect 520924 313216 520976 313268
rect 580172 313216 580224 313268
rect 530584 299412 530636 299464
rect 580172 299412 580224 299464
rect 3056 293904 3108 293956
rect 51724 293904 51776 293956
rect 547144 273164 547196 273216
rect 580172 273164 580224 273216
rect 3516 267656 3568 267708
rect 76564 267656 76616 267708
rect 519544 259360 519596 259412
rect 580172 259360 580224 259412
rect 2780 254328 2832 254380
rect 4896 254328 4948 254380
rect 551284 245556 551336 245608
rect 580172 245556 580224 245608
rect 3516 241408 3568 241460
rect 47584 241408 47636 241460
rect 544384 233180 544436 233232
rect 579988 233180 580040 233232
rect 518164 219376 518216 219428
rect 580172 219376 580224 219428
rect 3332 215228 3384 215280
rect 72424 215228 72476 215280
rect 529204 206932 529256 206984
rect 579804 206932 579856 206984
rect 2780 202716 2832 202768
rect 4804 202716 4856 202768
rect 543004 193128 543056 193180
rect 580172 193128 580224 193180
rect 3516 188980 3568 189032
rect 32404 188980 32456 189032
rect 515404 179324 515456 179376
rect 580172 179324 580224 179376
rect 526444 166948 526496 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 68284 164160 68336 164212
rect 540244 153144 540296 153196
rect 580172 153144 580224 153196
rect 3516 150356 3568 150408
rect 17224 150356 17276 150408
rect 512644 139340 512696 139392
rect 580172 139340 580224 139392
rect 80060 138388 80112 138440
rect 81026 138388 81078 138440
rect 161572 138388 161624 138440
rect 162814 138388 162866 138440
rect 3516 137912 3568 137964
rect 11704 137912 11756 137964
rect 54484 136552 54536 136604
rect 111984 136552 112036 136604
rect 115296 136552 115348 136604
rect 117964 136552 118016 136604
rect 124128 136552 124180 136604
rect 169668 136552 169720 136604
rect 170496 136552 170548 136604
rect 171416 136552 171468 136604
rect 180708 136552 180760 136604
rect 210976 136552 211028 136604
rect 213828 136552 213880 136604
rect 235080 136552 235132 136604
rect 238024 136552 238076 136604
rect 250628 136552 250680 136604
rect 274548 136552 274600 136604
rect 279056 136552 279108 136604
rect 315304 136552 315356 136604
rect 316684 136552 316736 136604
rect 403992 136552 404044 136604
rect 435364 136552 435416 136604
rect 68284 136484 68336 136536
rect 125784 136484 125836 136536
rect 126244 136484 126296 136536
rect 136088 136484 136140 136536
rect 142804 136484 142856 136536
rect 172244 136484 172296 136536
rect 173808 136484 173860 136536
rect 74448 136416 74500 136468
rect 133512 136416 133564 136468
rect 170404 136416 170456 136468
rect 173992 136416 174044 136468
rect 177856 136484 177908 136536
rect 209320 136484 209372 136536
rect 215208 136484 215260 136536
rect 236000 136484 236052 136536
rect 238668 136484 238720 136536
rect 253204 136484 253256 136536
rect 255964 136484 256016 136536
rect 263508 136484 263560 136536
rect 303252 136484 303304 136536
rect 306564 136484 306616 136536
rect 398748 136484 398800 136536
rect 429752 136484 429804 136536
rect 441068 136484 441120 136536
rect 443644 136484 443696 136536
rect 449624 136484 449676 136536
rect 506480 136484 506532 136536
rect 205824 136416 205876 136468
rect 211068 136416 211120 136468
rect 233424 136416 233476 136468
rect 235908 136416 235960 136468
rect 251456 136416 251508 136468
rect 256608 136416 256660 136468
rect 266084 136416 266136 136468
rect 286968 136416 287020 136468
rect 288532 136416 288584 136468
rect 393688 136416 393740 136468
rect 429936 136416 429988 136468
rect 453948 136416 454000 136468
rect 78496 136348 78548 136400
rect 136916 136348 136968 136400
rect 140780 136348 140832 136400
rect 145564 136348 145616 136400
rect 169576 136348 169628 136400
rect 203248 136348 203300 136400
rect 204904 136348 204956 136400
rect 228272 136348 228324 136400
rect 229008 136348 229060 136400
rect 246304 136348 246356 136400
rect 251088 136348 251140 136400
rect 261852 136348 261904 136400
rect 395436 136348 395488 136400
rect 444472 136348 444524 136400
rect 508596 136416 508648 136468
rect 511356 136348 511408 136400
rect 71688 136280 71740 136332
rect 131764 136280 131816 136332
rect 144184 136280 144236 136332
rect 181720 136280 181772 136332
rect 186964 136280 187016 136332
rect 192024 136280 192076 136332
rect 216220 136280 216272 136332
rect 216588 136280 216640 136332
rect 236828 136280 236880 136332
rect 237288 136280 237340 136332
rect 252376 136280 252428 136332
rect 253848 136280 253900 136332
rect 264428 136280 264480 136332
rect 267648 136280 267700 136332
rect 273904 136280 273956 136332
rect 400588 136280 400640 136332
rect 440240 136280 440292 136332
rect 451372 136280 451424 136332
rect 529204 136280 529256 136332
rect 51724 136212 51776 136264
rect 115388 136212 115440 136264
rect 117228 136212 117280 136264
rect 164516 136212 164568 136264
rect 166908 136212 166960 136264
rect 200672 136212 200724 136264
rect 202788 136212 202840 136264
rect 226524 136212 226576 136264
rect 227628 136212 227680 136264
rect 244556 136212 244608 136264
rect 246948 136212 247000 136264
rect 259276 136212 259328 136264
rect 263508 136212 263560 136264
rect 29644 136144 29696 136196
rect 93032 136144 93084 136196
rect 104164 136144 104216 136196
rect 109408 136144 109460 136196
rect 113088 136144 113140 136196
rect 161940 136144 161992 136196
rect 162768 136144 162820 136196
rect 198096 136144 198148 136196
rect 205548 136144 205600 136196
rect 229100 136144 229152 136196
rect 234528 136144 234580 136196
rect 249800 136144 249852 136196
rect 252468 136144 252520 136196
rect 262680 136144 262732 136196
rect 264244 136144 264296 136196
rect 267004 136144 267056 136196
rect 268752 136212 268804 136264
rect 271328 136144 271380 136196
rect 276664 136144 276716 136196
rect 279884 136144 279936 136196
rect 391112 136144 391164 136196
rect 399484 136144 399536 136196
rect 407488 136144 407540 136196
rect 448520 136212 448572 136264
rect 457444 136212 457496 136264
rect 517520 136212 517572 136264
rect 409144 136144 409196 136196
rect 450452 136144 450504 136196
rect 456524 136144 456576 136196
rect 464252 136144 464304 136196
rect 469496 136144 469548 136196
rect 482376 136144 482428 136196
rect 543004 136144 543056 136196
rect 32404 136076 32456 136128
rect 99012 136076 99064 136128
rect 107568 136076 107620 136128
rect 157616 136076 157668 136128
rect 160008 136076 160060 136128
rect 195520 136076 195572 136128
rect 202696 136076 202748 136128
rect 227352 136076 227404 136128
rect 227536 136076 227588 136128
rect 245476 136076 245528 136128
rect 249708 136076 249760 136128
rect 260932 136076 260984 136128
rect 264888 136076 264940 136128
rect 272156 136076 272208 136128
rect 273904 136076 273956 136128
rect 278228 136076 278280 136128
rect 385960 136076 386012 136128
rect 407764 136076 407816 136128
rect 17224 136008 17276 136060
rect 87880 136008 87932 136060
rect 93768 136008 93820 136060
rect 147312 136008 147364 136060
rect 148968 136008 149020 136060
rect 153108 136008 153160 136060
rect 187608 136008 187660 136060
rect 198648 136008 198700 136060
rect 223948 136008 224000 136060
rect 224868 136008 224920 136060
rect 242900 136008 242952 136060
rect 245568 136008 245620 136060
rect 258356 136008 258408 136060
rect 259368 136008 259420 136060
rect 267832 136008 267884 136060
rect 271788 136008 271840 136060
rect 277308 136008 277360 136060
rect 372988 136008 373040 136060
rect 395344 136008 395396 136060
rect 414388 136008 414440 136060
rect 18604 135940 18656 135992
rect 92204 135940 92256 135992
rect 95056 135940 95108 135992
rect 153016 135940 153068 135992
rect 195336 135940 195388 135992
rect 221372 135940 221424 135992
rect 223488 135940 223540 135992
rect 241980 135940 242032 135992
rect 242808 135940 242860 135992
rect 255780 135940 255832 135992
rect 7564 135872 7616 135924
rect 83556 135872 83608 135924
rect 88248 135872 88300 135924
rect 143816 135872 143868 135924
rect 148968 135872 149020 135924
rect 187792 135872 187844 135924
rect 191748 135872 191800 135924
rect 218796 135872 218848 135924
rect 222200 135872 222252 135924
rect 240324 135872 240376 135924
rect 241428 135872 241480 135924
rect 254952 135872 255004 135924
rect 255228 135872 255280 135924
rect 265256 135940 265308 135992
rect 267004 135940 267056 135992
rect 270408 135940 270460 135992
rect 305828 135940 305880 135992
rect 309232 135940 309284 135992
rect 314476 135940 314528 135992
rect 321652 135940 321704 135992
rect 336004 135940 336056 135992
rect 336648 135940 336700 135992
rect 365260 135940 365312 135992
rect 385684 135940 385736 135992
rect 391848 135940 391900 135992
rect 414664 135940 414716 135992
rect 416964 135940 417016 135992
rect 260748 135872 260800 135924
rect 277308 135872 277360 135924
rect 281632 135872 281684 135924
rect 333428 135872 333480 135924
rect 336096 135872 336148 135924
rect 352380 135872 352432 135924
rect 374092 135872 374144 135924
rect 378048 135872 378100 135924
rect 400864 135872 400916 135924
rect 402336 135872 402388 135924
rect 421564 135872 421616 135924
rect 422116 135940 422168 135992
rect 468484 136076 468536 136128
rect 474648 136076 474700 136128
rect 536104 136076 536156 136128
rect 457536 136008 457588 136060
rect 462596 136008 462648 136060
rect 524420 136008 524472 136060
rect 461584 135940 461636 135992
rect 467748 135940 467800 135992
rect 531320 135940 531372 135992
rect 81348 135804 81400 135856
rect 138664 135804 138716 135856
rect 146944 135804 146996 135856
rect 176568 135804 176620 135856
rect 177948 135804 178000 135856
rect 208400 135804 208452 135856
rect 209688 135804 209740 135856
rect 231676 135804 231728 135856
rect 231768 135804 231820 135856
rect 248052 135804 248104 135856
rect 260656 135804 260708 135856
rect 269580 135804 269632 135856
rect 399668 135804 399720 135856
rect 417424 135804 417476 135856
rect 424692 135804 424744 135856
rect 471244 135872 471296 135924
rect 472900 135872 472952 135924
rect 539600 135872 539652 135924
rect 431960 135804 432012 135856
rect 434996 135804 435048 135856
rect 65524 135736 65576 135788
rect 120540 135736 120592 135788
rect 125508 135736 125560 135788
rect 170588 135736 170640 135788
rect 190276 135736 190328 135788
rect 191196 135736 191248 135788
rect 204996 135736 205048 135788
rect 213184 135736 213236 135788
rect 234252 135736 234304 135788
rect 246304 135736 246356 135788
rect 254032 135736 254084 135788
rect 329932 135736 329984 135788
rect 336004 135736 336056 135788
rect 432420 135736 432472 135788
rect 86868 135668 86920 135720
rect 142068 135668 142120 135720
rect 180064 135668 180116 135720
rect 185216 135668 185268 135720
rect 199384 135668 199436 135720
rect 220084 135668 220136 135720
rect 224776 135668 224828 135720
rect 226248 135668 226300 135720
rect 243728 135668 243780 135720
rect 251824 135668 251876 135720
rect 260104 135668 260156 135720
rect 304908 135668 304960 135720
rect 305644 135668 305696 135720
rect 427268 135668 427320 135720
rect 436652 135668 436704 135720
rect 438492 135668 438544 135720
rect 486424 135804 486476 135856
rect 486700 135736 486752 135788
rect 520924 135804 520976 135856
rect 499488 135736 499540 135788
rect 526444 135736 526496 135788
rect 480628 135668 480680 135720
rect 481548 135668 481600 135720
rect 483204 135668 483256 135720
rect 484216 135668 484268 135720
rect 485872 135668 485924 135720
rect 487068 135668 487120 135720
rect 489276 135668 489328 135720
rect 489828 135668 489880 135720
rect 490104 135668 490156 135720
rect 491208 135668 491260 135720
rect 491852 135668 491904 135720
rect 493876 135668 493928 135720
rect 494428 135668 494480 135720
rect 522304 135668 522356 135720
rect 47584 135600 47636 135652
rect 101680 135600 101732 135652
rect 130384 135600 130436 135652
rect 153292 135600 153344 135652
rect 198004 135600 198056 135652
rect 199844 135600 199896 135652
rect 200764 135600 200816 135652
rect 202420 135600 202472 135652
rect 206928 135600 206980 135652
rect 229928 135600 229980 135652
rect 233148 135600 233200 135652
rect 248880 135600 248932 135652
rect 268936 135600 268988 135652
rect 274732 135600 274784 135652
rect 280804 135600 280856 135652
rect 283380 135600 283432 135652
rect 289820 135600 289872 135652
rect 291108 135600 291160 135652
rect 297180 135600 297232 135652
rect 298100 135600 298152 135652
rect 300676 135600 300728 135652
rect 302240 135600 302292 135652
rect 302424 135600 302476 135652
rect 305000 135600 305052 135652
rect 320456 135600 320508 135652
rect 321468 135600 321520 135652
rect 327356 135600 327408 135652
rect 328368 135600 328420 135652
rect 338580 135600 338632 135652
rect 339408 135600 339460 135652
rect 354956 135600 355008 135652
rect 356704 135600 356756 135652
rect 362684 135600 362736 135652
rect 363604 135600 363656 135652
rect 429844 135600 429896 135652
rect 72424 135532 72476 135584
rect 123208 135532 123260 135584
rect 137284 135532 137336 135584
rect 140412 135532 140464 135584
rect 75184 135464 75236 135516
rect 82728 135464 82780 135516
rect 83464 135464 83516 135516
rect 130016 135464 130068 135516
rect 133144 135464 133196 135516
rect 163688 135532 163740 135584
rect 188344 135532 188396 135584
rect 189448 135532 189500 135584
rect 184848 135464 184900 135516
rect 213552 135532 213604 135584
rect 217968 135532 218020 135584
rect 237748 135532 237800 135584
rect 249064 135532 249116 135584
rect 256700 135532 256752 135584
rect 269764 135532 269816 135584
rect 272984 135532 273036 135584
rect 282184 135532 282236 135584
rect 284208 135532 284260 135584
rect 284944 135532 284996 135584
rect 285956 135532 286008 135584
rect 288348 135532 288400 135584
rect 289360 135532 289412 135584
rect 289728 135532 289780 135584
rect 290280 135532 290332 135584
rect 292580 135532 292632 135584
rect 293684 135532 293736 135584
rect 298008 135532 298060 135584
rect 298744 135532 298796 135584
rect 298928 135532 298980 135584
rect 299572 135532 299624 135584
rect 299848 135532 299900 135584
rect 300768 135532 300820 135584
rect 301504 135532 301556 135584
rect 303620 135532 303672 135584
rect 304080 135532 304132 135584
rect 304908 135532 304960 135584
rect 306656 135532 306708 135584
rect 307668 135532 307720 135584
rect 309324 135532 309376 135584
rect 310336 135532 310388 135584
rect 310980 135532 311032 135584
rect 311716 135532 311768 135584
rect 312728 135532 312780 135584
rect 313188 135532 313240 135584
rect 313556 135532 313608 135584
rect 314568 135532 314620 135584
rect 316132 135532 316184 135584
rect 317328 135532 317380 135584
rect 317880 135532 317932 135584
rect 318708 135532 318760 135584
rect 319628 135532 319680 135584
rect 320824 135532 320876 135584
rect 322204 135532 322256 135584
rect 322848 135532 322900 135584
rect 323032 135532 323084 135584
rect 324228 135532 324280 135584
rect 324780 135532 324832 135584
rect 325608 135532 325660 135584
rect 326528 135532 326580 135584
rect 327724 135532 327776 135584
rect 329104 135532 329156 135584
rect 329748 135532 329800 135584
rect 331680 135532 331732 135584
rect 332416 135532 332468 135584
rect 334256 135532 334308 135584
rect 335176 135532 335228 135584
rect 336832 135532 336884 135584
rect 338764 135532 338816 135584
rect 340328 135532 340380 135584
rect 340788 135532 340840 135584
rect 341156 135532 341208 135584
rect 342168 135532 342220 135584
rect 342904 135532 342956 135584
rect 343548 135532 343600 135584
rect 343732 135532 343784 135584
rect 344928 135532 344980 135584
rect 345480 135532 345532 135584
rect 346308 135532 346360 135584
rect 347136 135532 347188 135584
rect 347688 135532 347740 135584
rect 348056 135532 348108 135584
rect 349068 135532 349120 135584
rect 349804 135532 349856 135584
rect 350448 135532 350500 135584
rect 350632 135532 350684 135584
rect 351736 135532 351788 135584
rect 354036 135532 354088 135584
rect 354588 135532 354640 135584
rect 356612 135532 356664 135584
rect 357348 135532 357400 135584
rect 357532 135532 357584 135584
rect 358636 135532 358688 135584
rect 359188 135532 359240 135584
rect 360108 135532 360160 135584
rect 360936 135532 360988 135584
rect 361488 135532 361540 135584
rect 361856 135532 361908 135584
rect 362868 135532 362920 135584
rect 363512 135532 363564 135584
rect 364248 135532 364300 135584
rect 364432 135532 364484 135584
rect 365628 135532 365680 135584
rect 366088 135532 366140 135584
rect 367008 135532 367060 135584
rect 367836 135532 367888 135584
rect 368388 135532 368440 135584
rect 368664 135532 368716 135584
rect 369768 135532 369820 135584
rect 370412 135532 370464 135584
rect 371148 135532 371200 135584
rect 371332 135532 371384 135584
rect 372436 135532 372488 135584
rect 374736 135532 374788 135584
rect 375288 135532 375340 135584
rect 375564 135532 375616 135584
rect 376576 135532 376628 135584
rect 381636 135532 381688 135584
rect 382188 135532 382240 135584
rect 382464 135532 382516 135584
rect 383568 135532 383620 135584
rect 384212 135532 384264 135584
rect 384948 135532 385000 135584
rect 386788 135532 386840 135584
rect 387616 135532 387668 135584
rect 388536 135532 388588 135584
rect 389088 135532 389140 135584
rect 389364 135532 389416 135584
rect 390468 135532 390520 135584
rect 396264 135532 396316 135584
rect 397368 135532 397420 135584
rect 398012 135532 398064 135584
rect 398748 135532 398800 135584
rect 403164 135532 403216 135584
rect 404268 135532 404320 135584
rect 404912 135532 404964 135584
rect 406384 135532 406436 135584
rect 406568 135532 406620 135584
rect 407028 135532 407080 135584
rect 418620 135532 418672 135584
rect 419448 135532 419500 135584
rect 420368 135532 420420 135584
rect 420828 135532 420880 135584
rect 421196 135532 421248 135584
rect 422208 135532 422260 135584
rect 422944 135532 422996 135584
rect 423588 135532 423640 135584
rect 423864 135532 423916 135584
rect 424968 135532 425020 135584
rect 428096 135532 428148 135584
rect 429108 135532 429160 135584
rect 430672 135532 430724 135584
rect 431776 135532 431828 135584
rect 434168 135532 434220 135584
rect 434628 135532 434680 135584
rect 436744 135532 436796 135584
rect 437388 135532 437440 135584
rect 437572 135532 437624 135584
rect 438768 135532 438820 135584
rect 439320 135532 439372 135584
rect 440148 135532 440200 135584
rect 441896 135532 441948 135584
rect 442908 135532 442960 135584
rect 446220 135532 446272 135584
rect 446956 135532 447008 135584
rect 447968 135532 448020 135584
rect 448428 135532 448480 135584
rect 448796 135532 448848 135584
rect 449808 135532 449860 135584
rect 191104 135464 191156 135516
rect 220728 135464 220780 135516
rect 224224 135464 224276 135516
rect 232504 135464 232556 135516
rect 233884 135464 233936 135516
rect 247224 135464 247276 135516
rect 251916 135464 251968 135516
rect 257528 135464 257580 135516
rect 269028 135464 269080 135516
rect 275560 135464 275612 135516
rect 278688 135464 278740 135516
rect 282460 135464 282512 135516
rect 308404 135464 308456 135516
rect 313372 135464 313424 135516
rect 317052 135464 317104 135516
rect 324504 135464 324556 135516
rect 337660 135464 337712 135516
rect 340144 135464 340196 135516
rect 377312 135464 377364 135516
rect 378048 135464 378100 135516
rect 380808 135464 380860 135516
rect 381544 135464 381596 135516
rect 425520 135464 425572 135516
rect 426348 135464 426400 135516
rect 443552 135464 443604 135516
rect 450544 135464 450596 135516
rect 451188 135464 451240 135516
rect 76932 135396 76984 135448
rect 95608 135396 95660 135448
rect 219348 135396 219400 135448
rect 238576 135396 238628 135448
rect 270408 135396 270460 135448
rect 276480 135396 276532 135448
rect 453120 135600 453172 135652
rect 453948 135600 454000 135652
rect 454868 135600 454920 135652
rect 455328 135600 455380 135652
rect 455696 135600 455748 135652
rect 456708 135600 456760 135652
rect 466920 135600 466972 135652
rect 467748 135600 467800 135652
rect 468576 135600 468628 135652
rect 469128 135600 469180 135652
rect 457444 135464 457496 135516
rect 466000 135464 466052 135516
rect 512644 135600 512696 135652
rect 471152 135532 471204 135584
rect 471888 135532 471940 135584
rect 472072 135532 472124 135584
rect 473268 135532 473320 135584
rect 475476 135532 475528 135584
rect 476028 135532 476080 135584
rect 478052 135532 478104 135584
rect 478788 135532 478840 135584
rect 473820 135464 473872 135516
rect 475384 135396 475436 135448
rect 476396 135464 476448 135516
rect 519544 135532 519596 135584
rect 515404 135464 515456 135516
rect 485044 135396 485096 135448
rect 496176 135396 496228 135448
rect 496728 135396 496780 135448
rect 499580 135396 499632 135448
rect 501328 135396 501380 135448
rect 502156 135396 502208 135448
rect 503076 135396 503128 135448
rect 503628 135396 503680 135448
rect 503904 135396 503956 135448
rect 505008 135396 505060 135448
rect 79324 135328 79376 135380
rect 88708 135328 88760 135380
rect 228364 135328 228416 135380
rect 241152 135328 241204 135380
rect 379888 135328 379940 135380
rect 380808 135328 380860 135380
rect 482284 135328 482336 135380
rect 498752 135328 498804 135380
rect 499488 135328 499540 135380
rect 231124 135260 231176 135312
rect 239404 135260 239456 135312
rect 410064 135260 410116 135312
rect 411168 135260 411220 135312
rect 411812 135260 411864 135312
rect 412456 135260 412508 135312
rect 413468 135260 413520 135312
rect 413928 135260 413980 135312
rect 416044 135260 416096 135312
rect 416688 135260 416740 135312
rect 458272 135260 458324 135312
rect 459376 135260 459428 135312
rect 460020 135260 460072 135312
rect 460848 135260 460900 135312
rect 461676 135260 461728 135312
rect 462228 135260 462280 135312
rect 464344 135260 464396 135312
rect 464988 135260 465040 135312
rect 465172 135260 465224 135312
rect 466368 135260 466420 135312
rect 481456 135260 481508 135312
rect 488632 135260 488684 135312
rect 43444 135124 43496 135176
rect 96436 135124 96488 135176
rect 22008 135056 22060 135108
rect 76932 135056 76984 135108
rect 77208 135056 77260 135108
rect 135168 135056 135220 135108
rect 53748 134988 53800 135040
rect 115296 134988 115348 135040
rect 487528 134988 487580 135040
rect 547144 134988 547196 135040
rect 62028 134920 62080 134972
rect 124864 134920 124916 134972
rect 459100 134920 459152 134972
rect 520280 134920 520332 134972
rect 41328 134852 41380 134904
rect 104164 134852 104216 134904
rect 488632 134852 488684 134904
rect 550640 134852 550692 134904
rect 39396 134784 39448 134836
rect 102508 134784 102560 134836
rect 477224 134784 477276 134836
rect 544384 134784 544436 134836
rect 35164 134716 35216 134768
rect 99932 134716 99984 134768
rect 478972 134716 479024 134768
rect 547880 134716 547932 134768
rect 37188 134648 37240 134700
rect 106832 134648 106884 134700
rect 484124 134648 484176 134700
rect 554780 134648 554832 134700
rect 15844 134580 15896 134632
rect 89536 134580 89588 134632
rect 135168 134580 135220 134632
rect 177396 134580 177448 134632
rect 493876 134580 493928 134632
rect 564532 134580 564584 134632
rect 11704 134512 11756 134564
rect 86132 134512 86184 134564
rect 91008 134512 91060 134564
rect 140780 134512 140832 134564
rect 142068 134512 142120 134564
rect 182548 134512 182600 134564
rect 497004 134512 497056 134564
rect 572812 134512 572864 134564
rect 57244 133152 57296 133204
rect 105084 133152 105136 133204
rect 484952 133152 485004 133204
rect 556252 133152 556304 133204
rect 511264 126896 511316 126948
rect 580172 126896 580224 126948
rect 538864 113092 538916 113144
rect 579804 113092 579856 113144
rect 3148 111732 3200 111784
rect 58624 111732 58676 111784
rect 560944 100648 560996 100700
rect 580172 100648 580224 100700
rect 3516 97928 3568 97980
rect 22744 97928 22796 97980
rect 508504 86912 508556 86964
rect 580172 86912 580224 86964
rect 3516 85484 3568 85536
rect 25504 85484 25556 85536
rect 3516 71680 3568 71732
rect 69664 71680 69716 71732
rect 70308 71000 70360 71052
rect 130936 71000 130988 71052
rect 558184 60664 558236 60716
rect 580172 60664 580224 60716
rect 473268 48968 473320 49020
rect 538220 48968 538272 49020
rect 446956 47540 447008 47592
rect 502340 47540 502392 47592
rect 3424 45500 3476 45552
rect 39304 45500 39356 45552
rect 3148 33056 3200 33108
rect 50344 33056 50396 33108
rect 50436 32376 50488 32428
rect 107660 32376 107712 32428
rect 35256 26868 35308 26920
rect 104256 26868 104308 26920
rect 104808 25508 104860 25560
rect 155868 25508 155920 25560
rect 97908 24080 97960 24132
rect 150716 24080 150768 24132
rect 3424 20612 3476 20664
rect 14464 20612 14516 20664
rect 368388 15852 368440 15904
rect 395252 15852 395304 15904
rect 436008 15852 436060 15904
rect 488816 15852 488868 15904
rect 489828 15852 489880 15904
rect 562048 15852 562100 15904
rect 381544 14424 381596 14476
rect 412640 14424 412692 14476
rect 471888 14424 471940 14476
rect 537208 14424 537260 14476
rect 376576 11704 376628 11756
rect 406016 11704 406068 11756
rect 406384 11704 406436 11756
rect 445760 11704 445812 11756
rect 449808 11704 449860 11756
rect 506572 11704 506624 11756
rect 512644 11704 512696 11756
rect 530124 11704 530176 11756
rect 526444 10276 526496 10328
rect 575848 10276 575900 10328
rect 4068 8916 4120 8968
rect 75184 8916 75236 8968
rect 83280 8916 83332 8968
rect 137284 8916 137336 8968
rect 137652 8916 137704 8968
rect 179972 8916 180024 8968
rect 363604 8916 363656 8968
rect 388260 8916 388312 8968
rect 469128 8916 469180 8968
rect 533712 8916 533764 8968
rect 132960 7692 133012 7744
rect 146944 7692 146996 7744
rect 115204 7624 115256 7676
rect 133144 7624 133196 7676
rect 147128 7624 147180 7676
rect 186872 7624 186924 7676
rect 397276 7624 397328 7676
rect 435548 7624 435600 7676
rect 520924 7624 520976 7676
rect 558552 7624 558604 7676
rect 12348 7556 12400 7608
rect 79324 7556 79376 7608
rect 111616 7556 111668 7608
rect 161020 7556 161072 7608
rect 358636 7556 358688 7608
rect 381176 7556 381228 7608
rect 419356 7556 419408 7608
rect 466276 7556 466328 7608
rect 522304 7556 522356 7608
rect 569132 7556 569184 7608
rect 3424 6808 3476 6860
rect 33784 6808 33836 6860
rect 431776 6604 431828 6656
rect 481732 6604 481784 6656
rect 433248 6536 433300 6588
rect 485228 6536 485280 6588
rect 144736 6468 144788 6520
rect 180064 6468 180116 6520
rect 464344 6468 464396 6520
rect 517152 6468 517204 6520
rect 138848 6400 138900 6452
rect 180892 6400 180944 6452
rect 443644 6400 443696 6452
rect 495900 6400 495952 6452
rect 519544 6400 519596 6452
rect 544292 6400 544344 6452
rect 122380 6332 122432 6384
rect 168840 6332 168892 6384
rect 462228 6332 462280 6384
rect 524236 6332 524288 6384
rect 118792 6264 118844 6316
rect 166264 6264 166316 6316
rect 464988 6264 465040 6316
rect 527824 6264 527876 6316
rect 108120 6196 108172 6248
rect 158444 6196 158496 6248
rect 467748 6196 467800 6248
rect 531320 6196 531372 6248
rect 69112 6128 69164 6180
rect 83464 6128 83516 6180
rect 86868 6128 86920 6180
rect 142988 6128 143040 6180
rect 142436 6060 142488 6112
rect 183468 6128 183520 6180
rect 436744 6128 436796 6180
rect 476948 6128 477000 6180
rect 480076 6128 480128 6180
rect 549076 6128 549128 6180
rect 59636 5448 59688 5500
rect 72424 5448 72476 5500
rect 72608 5448 72660 5500
rect 132684 5448 132736 5500
rect 161296 5448 161348 5500
rect 197268 5448 197320 5500
rect 438768 5448 438820 5500
rect 491024 5448 491076 5500
rect 65616 5380 65668 5432
rect 127440 5380 127492 5432
rect 135260 5380 135312 5432
rect 178316 5380 178368 5432
rect 414664 5380 414716 5432
rect 428464 5380 428516 5432
rect 440056 5380 440108 5432
rect 494704 5380 494756 5432
rect 56048 5312 56100 5364
rect 65524 5312 65576 5364
rect 66720 5312 66772 5364
rect 128360 5312 128412 5364
rect 129372 5312 129424 5364
rect 170404 5312 170456 5364
rect 407764 5312 407816 5364
rect 420184 5312 420236 5364
rect 421564 5312 421616 5364
rect 442632 5312 442684 5364
rect 445668 5312 445720 5364
rect 501788 5312 501840 5364
rect 58440 5244 58492 5296
rect 122288 5244 122340 5296
rect 136456 5244 136508 5296
rect 179144 5244 179196 5296
rect 399484 5244 399536 5296
rect 427268 5244 427320 5296
rect 442816 5244 442868 5296
rect 498200 5244 498252 5296
rect 44272 5176 44324 5228
rect 54484 5176 54536 5228
rect 54944 5176 54996 5228
rect 119712 5176 119764 5228
rect 131764 5176 131816 5228
rect 175740 5176 175792 5228
rect 383476 5176 383528 5228
rect 416688 5176 416740 5228
rect 417424 5176 417476 5228
rect 439136 5176 439188 5228
rect 448428 5176 448480 5228
rect 505376 5176 505428 5228
rect 51356 5108 51408 5160
rect 117136 5108 117188 5160
rect 130568 5108 130620 5160
rect 174820 5108 174872 5160
rect 389088 5108 389140 5160
rect 423772 5108 423824 5160
rect 429844 5108 429896 5160
rect 437940 5108 437992 5160
rect 451188 5108 451240 5160
rect 508872 5108 508924 5160
rect 30104 5040 30156 5092
rect 47584 5040 47636 5092
rect 47860 5040 47912 5092
rect 114560 5040 114612 5092
rect 125876 5040 125928 5092
rect 170496 5040 170548 5092
rect 171968 5040 172020 5092
rect 191104 5040 191156 5092
rect 397368 5040 397420 5092
rect 7656 4972 7708 5024
rect 85304 4972 85356 5024
rect 128176 4972 128228 5024
rect 173072 4972 173124 5024
rect 394608 4972 394660 5024
rect 432052 5040 432104 5092
rect 453948 5040 454000 5092
rect 512460 5040 512512 5092
rect 435364 4972 435416 5024
rect 445024 4972 445076 5024
rect 456708 4972 456760 5024
rect 1676 4904 1728 4956
rect 80060 4904 80112 4956
rect 93952 4904 94004 4956
rect 148140 4904 148192 4956
rect 157800 4904 157852 4956
rect 194692 4904 194744 4956
rect 356704 4904 356756 4956
rect 377680 4904 377732 4956
rect 401508 4904 401560 4956
rect 441528 4904 441580 4956
rect 459376 4904 459428 4956
rect 515404 4972 515456 5024
rect 540796 4972 540848 5024
rect 515956 4904 516008 4956
rect 2872 4836 2924 4888
rect 81808 4836 81860 4888
rect 91560 4836 91612 4888
rect 146392 4836 146444 4888
rect 150624 4836 150676 4888
rect 188344 4836 188396 4888
rect 360016 4836 360068 4888
rect 384764 4836 384816 4888
rect 407028 4836 407080 4888
rect 448612 4836 448664 4888
rect 463608 4836 463660 4888
rect 526628 4836 526680 4888
rect 572 4768 624 4820
rect 80152 4768 80204 4820
rect 84476 4768 84528 4820
rect 141240 4768 141292 4820
rect 143540 4768 143592 4820
rect 184296 4768 184348 4820
rect 371148 4768 371200 4820
rect 398932 4768 398984 4820
rect 400864 4768 400916 4820
rect 409604 4768 409656 4820
rect 412456 4768 412508 4820
rect 455696 4768 455748 4820
rect 460756 4768 460808 4820
rect 523040 4768 523092 4820
rect 536104 4768 536156 4820
rect 541992 4768 542044 4820
rect 543004 4768 543056 4820
rect 552664 4768 552716 4820
rect 63224 4700 63276 4752
rect 68284 4700 68336 4752
rect 79692 4700 79744 4752
rect 137836 4700 137888 4752
rect 154212 4700 154264 4752
rect 186964 4700 187016 4752
rect 434444 4700 434496 4752
rect 475384 4700 475436 4752
rect 499396 4700 499448 4752
rect 508596 4700 508648 4752
rect 510068 4700 510120 4752
rect 519544 4700 519596 4752
rect 77392 4632 77444 4684
rect 126244 4632 126296 4684
rect 126980 4632 127032 4684
rect 142804 4632 142856 4684
rect 164884 4632 164936 4684
rect 198004 4632 198056 4684
rect 457444 4632 457496 4684
rect 480536 4632 480588 4684
rect 486424 4632 486476 4684
rect 492312 4632 492364 4684
rect 101036 4564 101088 4616
rect 130384 4564 130436 4616
rect 168380 4564 168432 4616
rect 200764 4564 200816 4616
rect 140044 4496 140096 4548
rect 144184 4496 144236 4548
rect 450544 4360 450596 4412
rect 452108 4360 452160 4412
rect 26516 4156 26568 4208
rect 32404 4156 32456 4208
rect 48964 4156 49016 4208
rect 51724 4156 51776 4208
rect 87052 4156 87104 4208
rect 94044 4156 94096 4208
rect 41880 4088 41932 4140
rect 110236 4088 110288 4140
rect 385684 4156 385736 4208
rect 391848 4156 391900 4208
rect 395344 4156 395396 4208
rect 402520 4156 402572 4208
rect 429936 4156 429988 4208
rect 430856 4156 430908 4208
rect 431960 4156 432012 4208
rect 433248 4156 433300 4208
rect 457536 4156 457588 4208
rect 459192 4156 459244 4208
rect 461584 4156 461636 4208
rect 462780 4156 462832 4208
rect 468484 4156 468536 4208
rect 469864 4156 469916 4208
rect 471244 4156 471296 4208
rect 473452 4156 473504 4208
rect 482284 4156 482336 4208
rect 484032 4156 484084 4208
rect 485044 4156 485096 4208
rect 487620 4156 487672 4208
rect 506480 4156 506532 4208
rect 507676 4156 507728 4208
rect 511356 4156 511408 4208
rect 513564 4156 513616 4208
rect 529204 4156 529256 4208
rect 534908 4156 534960 4208
rect 112812 4088 112864 4140
rect 31300 4020 31352 4072
rect 39396 4020 39448 4072
rect 43076 4020 43128 4072
rect 23020 3952 23072 4004
rect 43444 3952 43496 4004
rect 46664 3952 46716 4004
rect 109316 4020 109368 4072
rect 159364 4088 159416 4140
rect 175464 4088 175516 4140
rect 207572 4088 207624 4140
rect 285404 4088 285456 4140
rect 287704 4088 287756 4140
rect 296628 4088 296680 4140
rect 297272 4088 297324 4140
rect 304908 4088 304960 4140
rect 307944 4088 307996 4140
rect 335268 4088 335320 4140
rect 350448 4088 350500 4140
rect 353208 4088 353260 4140
rect 375288 4088 375340 4140
rect 382188 4088 382240 4140
rect 410800 4088 410852 4140
rect 419448 4088 419500 4140
rect 465172 4088 465224 4140
rect 487068 4088 487120 4140
rect 557356 4088 557408 4140
rect 167000 4020 167052 4072
rect 179052 4020 179104 4072
rect 111064 3952 111116 4004
rect 114008 3952 114060 4004
rect 161572 3952 161624 4004
rect 174268 3952 174320 4004
rect 206744 3952 206796 4004
rect 35992 3884 36044 3936
rect 100760 3884 100812 3936
rect 102232 3884 102284 3936
rect 149888 3884 149940 3936
rect 5264 3816 5316 3868
rect 7564 3816 7616 3868
rect 39580 3816 39632 3868
rect 108488 3816 108540 3868
rect 110512 3816 110564 3868
rect 160100 3884 160152 3936
rect 170772 3884 170824 3936
rect 204076 3884 204128 3936
rect 167184 3816 167236 3868
rect 311808 4020 311860 4072
rect 318524 4020 318576 4072
rect 322848 4020 322900 4072
rect 332692 4020 332744 4072
rect 342168 4020 342220 4072
rect 358636 4020 358688 4072
rect 360108 4020 360160 4072
rect 383476 4020 383528 4072
rect 324136 3952 324188 4004
rect 335084 3952 335136 4004
rect 336648 3952 336700 4004
rect 351644 3952 351696 4004
rect 357348 3952 357400 4004
rect 379980 3952 380032 4004
rect 383568 3952 383620 4004
rect 415492 4020 415544 4072
rect 420828 4020 420880 4072
rect 467472 4020 467524 4072
rect 491208 4020 491260 4072
rect 563244 4020 563296 4072
rect 414296 3952 414348 4004
rect 418068 3952 418120 4004
rect 463976 3952 464028 4004
rect 488356 3952 488408 4004
rect 560852 3952 560904 4004
rect 305644 3884 305696 3936
rect 309048 3884 309100 3936
rect 328368 3884 328420 3936
rect 339868 3884 339920 3936
rect 340788 3884 340840 3936
rect 357532 3884 357584 3936
rect 362868 3884 362920 3936
rect 210148 3816 210200 3868
rect 18236 3748 18288 3800
rect 29644 3748 29696 3800
rect 32404 3748 32456 3800
rect 28908 3680 28960 3732
rect 105636 3748 105688 3800
rect 105728 3748 105780 3800
rect 156788 3748 156840 3800
rect 160100 3748 160152 3800
rect 196348 3748 196400 3800
rect 103244 3680 103296 3732
rect 103336 3680 103388 3732
rect 155040 3680 155092 3732
rect 163688 3680 163740 3732
rect 198924 3748 198976 3800
rect 209780 3748 209832 3800
rect 224224 3816 224276 3868
rect 313188 3816 313240 3868
rect 319720 3816 319772 3868
rect 321468 3816 321520 3868
rect 330392 3816 330444 3868
rect 331128 3816 331180 3868
rect 344560 3816 344612 3868
rect 346308 3816 346360 3868
rect 364616 3816 364668 3868
rect 367008 3816 367060 3868
rect 384948 3884 385000 3936
rect 417884 3884 417936 3936
rect 424876 3884 424928 3936
rect 472256 3884 472308 3936
rect 492588 3884 492640 3936
rect 566832 3884 566884 3936
rect 387156 3816 387208 3868
rect 390468 3816 390520 3868
rect 424968 3816 425020 3868
rect 426348 3816 426400 3868
rect 474556 3816 474608 3868
rect 493968 3816 494020 3868
rect 568028 3816 568080 3868
rect 230848 3748 230900 3800
rect 327724 3748 327776 3800
rect 338672 3748 338724 3800
rect 339408 3748 339460 3800
rect 355232 3748 355284 3800
rect 355968 3748 356020 3800
rect 378876 3748 378928 3800
rect 379428 3748 379480 3800
rect 384856 3748 384908 3800
rect 418988 3748 419040 3800
rect 423588 3748 423640 3800
rect 471060 3748 471112 3800
rect 491116 3748 491168 3800
rect 564440 3748 564492 3800
rect 196808 3680 196860 3732
rect 24216 3612 24268 3664
rect 97356 3612 97408 3664
rect 97448 3612 97500 3664
rect 97908 3612 97960 3664
rect 98644 3612 98696 3664
rect 151544 3612 151596 3664
rect 156604 3612 156656 3664
rect 193772 3612 193824 3664
rect 195612 3612 195664 3664
rect 199384 3612 199436 3664
rect 200304 3680 200356 3732
rect 225696 3680 225748 3732
rect 314568 3680 314620 3732
rect 320916 3680 320968 3732
rect 321008 3680 321060 3732
rect 329196 3680 329248 3732
rect 329748 3680 329800 3732
rect 223028 3612 223080 3664
rect 318616 3612 318668 3664
rect 325516 3612 325568 3664
rect 337476 3612 337528 3664
rect 339316 3612 339368 3664
rect 342076 3680 342128 3732
rect 359924 3680 359976 3732
rect 361488 3680 361540 3732
rect 385960 3680 386012 3732
rect 387708 3680 387760 3732
rect 25320 3544 25372 3596
rect 98184 3544 98236 3596
rect 99840 3544 99892 3596
rect 154120 3544 154172 3596
rect 155408 3544 155460 3596
rect 17040 3476 17092 3528
rect 18604 3476 18656 3528
rect 19432 3476 19484 3528
rect 9956 3408 10008 3460
rect 85672 3476 85724 3528
rect 86684 3476 86736 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 96252 3476 96304 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 151820 3476 151872 3528
rect 153108 3476 153160 3528
rect 158904 3476 158956 3528
rect 160008 3476 160060 3528
rect 166080 3476 166132 3528
rect 166908 3476 166960 3528
rect 173164 3476 173216 3528
rect 173808 3476 173860 3528
rect 176660 3476 176712 3528
rect 177948 3476 178000 3528
rect 180248 3476 180300 3528
rect 180708 3476 180760 3528
rect 89168 3408 89220 3460
rect 134156 3408 134208 3460
rect 135168 3408 135220 3460
rect 141240 3408 141292 3460
rect 142068 3408 142120 3460
rect 145932 3408 145984 3460
rect 11152 3340 11204 3392
rect 17224 3340 17276 3392
rect 33600 3340 33652 3392
rect 35256 3340 35308 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 45468 3340 45520 3392
rect 106924 3340 106976 3392
rect 107568 3340 107620 3392
rect 113732 3340 113784 3392
rect 116400 3340 116452 3392
rect 117228 3340 117280 3392
rect 121092 3340 121144 3392
rect 167920 3340 167972 3392
rect 52552 3272 52604 3324
rect 53748 3272 53800 3324
rect 116308 3272 116360 3324
rect 117596 3272 117648 3324
rect 165344 3272 165396 3324
rect 8760 3204 8812 3256
rect 11704 3204 11756 3256
rect 38384 3204 38436 3256
rect 50436 3204 50488 3256
rect 118884 3204 118936 3256
rect 119896 3204 119948 3256
rect 123484 3204 123536 3256
rect 124128 3204 124180 3256
rect 124680 3204 124732 3256
rect 125508 3204 125560 3256
rect 144644 3204 144696 3256
rect 152464 3204 152516 3256
rect 13544 3136 13596 3188
rect 15844 3136 15896 3188
rect 53748 3136 53800 3188
rect 57244 3136 57296 3188
rect 121644 3136 121696 3188
rect 149520 3136 149572 3188
rect 183744 3408 183796 3460
rect 184848 3408 184900 3460
rect 201592 3544 201644 3596
rect 207388 3544 207440 3596
rect 221556 3544 221608 3596
rect 228364 3544 228416 3596
rect 247592 3544 247644 3596
rect 251824 3544 251876 3596
rect 267740 3544 267792 3596
rect 268936 3544 268988 3596
rect 318708 3544 318760 3596
rect 326804 3544 326856 3596
rect 328276 3544 328328 3596
rect 340972 3544 341024 3596
rect 342168 3612 342220 3664
rect 356336 3612 356388 3664
rect 358728 3612 358780 3664
rect 382372 3612 382424 3664
rect 387616 3612 387668 3664
rect 421380 3680 421432 3732
rect 429108 3680 429160 3732
rect 478144 3680 478196 3732
rect 495348 3680 495400 3732
rect 570328 3680 570380 3732
rect 422576 3612 422628 3664
rect 426256 3612 426308 3664
rect 475752 3612 475804 3664
rect 499488 3612 499540 3664
rect 575112 3612 575164 3664
rect 344836 3544 344888 3596
rect 363512 3544 363564 3596
rect 364248 3544 364300 3596
rect 389456 3544 389508 3596
rect 393044 3544 393096 3596
rect 393228 3544 393280 3596
rect 429660 3544 429712 3596
rect 431868 3544 431920 3596
rect 482836 3544 482888 3596
rect 496728 3544 496780 3596
rect 571524 3544 571576 3596
rect 188528 3476 188580 3528
rect 192944 3408 192996 3460
rect 194416 3408 194468 3460
rect 195244 3408 195296 3460
rect 197912 3408 197964 3460
rect 198648 3408 198700 3460
rect 201500 3476 201552 3528
rect 202788 3476 202840 3528
rect 203892 3476 203944 3528
rect 204904 3476 204956 3528
rect 205088 3476 205140 3528
rect 205548 3476 205600 3528
rect 206192 3476 206244 3528
rect 206928 3476 206980 3528
rect 208584 3476 208636 3528
rect 209688 3476 209740 3528
rect 212172 3476 212224 3528
rect 213184 3476 213236 3528
rect 213368 3476 213420 3528
rect 213828 3476 213880 3528
rect 214472 3476 214524 3528
rect 215208 3476 215260 3528
rect 215668 3476 215720 3528
rect 216588 3476 216640 3528
rect 216864 3476 216916 3528
rect 217968 3476 218020 3528
rect 218060 3476 218112 3528
rect 219348 3476 219400 3528
rect 222752 3476 222804 3528
rect 223488 3476 223540 3528
rect 225144 3476 225196 3528
rect 226248 3476 226300 3528
rect 226340 3476 226392 3528
rect 227628 3476 227680 3528
rect 231032 3476 231084 3528
rect 231768 3476 231820 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 238116 3476 238168 3528
rect 238668 3476 238720 3528
rect 240508 3476 240560 3528
rect 241428 3476 241480 3528
rect 248788 3476 248840 3528
rect 249708 3476 249760 3528
rect 249984 3476 250036 3528
rect 251088 3476 251140 3528
rect 251180 3476 251232 3528
rect 252468 3476 252520 3528
rect 254676 3476 254728 3528
rect 255228 3476 255280 3528
rect 255872 3476 255924 3528
rect 256608 3476 256660 3528
rect 258264 3476 258316 3528
rect 259368 3476 259420 3528
rect 259460 3476 259512 3528
rect 260748 3476 260800 3528
rect 262956 3476 263008 3528
rect 263508 3476 263560 3528
rect 264152 3476 264204 3528
rect 264888 3476 264940 3528
rect 266544 3476 266596 3528
rect 267648 3476 267700 3528
rect 273628 3476 273680 3528
rect 274548 3476 274600 3528
rect 279516 3476 279568 3528
rect 280804 3476 280856 3528
rect 288992 3476 289044 3528
rect 289728 3476 289780 3528
rect 291384 3476 291436 3528
rect 291936 3476 291988 3528
rect 292580 3476 292632 3528
rect 293684 3476 293736 3528
rect 295340 3476 295392 3528
rect 296076 3476 296128 3528
rect 298744 3476 298796 3528
rect 299664 3476 299716 3528
rect 300768 3476 300820 3528
rect 301964 3476 302016 3528
rect 310336 3476 310388 3528
rect 315028 3476 315080 3528
rect 321376 3476 321428 3528
rect 217048 3408 217100 3460
rect 181444 3340 181496 3392
rect 211896 3340 211948 3392
rect 219256 3340 219308 3392
rect 231124 3408 231176 3460
rect 244096 3408 244148 3460
rect 251916 3408 251968 3460
rect 257068 3408 257120 3460
rect 264244 3408 264296 3460
rect 272432 3408 272484 3460
rect 273904 3408 273956 3460
rect 276020 3408 276072 3460
rect 280160 3408 280212 3460
rect 280712 3408 280764 3460
rect 282184 3408 282236 3460
rect 307576 3408 307628 3460
rect 312636 3408 312688 3460
rect 317328 3408 317380 3460
rect 324412 3408 324464 3460
rect 328000 3476 328052 3528
rect 332416 3476 332468 3528
rect 345756 3476 345808 3528
rect 346216 3476 346268 3528
rect 365812 3476 365864 3528
rect 369676 3476 369728 3528
rect 397736 3476 397788 3528
rect 398748 3476 398800 3528
rect 436744 3476 436796 3528
rect 437388 3476 437440 3528
rect 489920 3476 489972 3528
rect 498016 3476 498068 3528
rect 573916 3476 573968 3528
rect 331588 3408 331640 3460
rect 335176 3408 335228 3460
rect 349252 3408 349304 3460
rect 351828 3408 351880 3460
rect 372896 3408 372948 3460
rect 373908 3408 373960 3460
rect 403624 3408 403676 3460
rect 404268 3408 404320 3460
rect 443828 3408 443880 3460
rect 447048 3408 447100 3460
rect 504180 3408 504232 3460
rect 505008 3408 505060 3460
rect 583392 3408 583444 3460
rect 332508 3340 332560 3392
rect 346952 3340 347004 3392
rect 349068 3340 349120 3392
rect 354588 3340 354640 3392
rect 376484 3340 376536 3392
rect 376668 3340 376720 3392
rect 407212 3340 407264 3392
rect 422208 3340 422260 3392
rect 468668 3340 468720 3392
rect 484216 3340 484268 3392
rect 553768 3340 553820 3392
rect 182548 3272 182600 3324
rect 212724 3272 212776 3324
rect 229836 3272 229888 3324
rect 233884 3272 233936 3324
rect 234620 3272 234672 3324
rect 238024 3272 238076 3324
rect 246396 3272 246448 3324
rect 246948 3272 247000 3324
rect 184940 3204 184992 3256
rect 214380 3204 214432 3256
rect 223948 3204 224000 3256
rect 224868 3204 224920 3256
rect 241704 3204 241756 3256
rect 242808 3204 242860 3256
rect 242900 3204 242952 3256
rect 249064 3272 249116 3324
rect 252376 3272 252428 3324
rect 255964 3272 256016 3324
rect 271236 3272 271288 3324
rect 271788 3272 271840 3324
rect 287796 3272 287848 3324
rect 288348 3272 288400 3324
rect 307668 3272 307720 3324
rect 311440 3272 311492 3324
rect 325608 3272 325660 3324
rect 336280 3272 336332 3324
rect 324228 3204 324280 3256
rect 333888 3204 333940 3256
rect 34796 3068 34848 3120
rect 50160 3068 50212 3120
rect 64328 3068 64380 3120
rect 126612 3068 126664 3120
rect 186044 3136 186096 3188
rect 189724 3136 189776 3188
rect 217876 3136 217928 3188
rect 265348 3136 265400 3188
rect 269764 3136 269816 3188
rect 284300 3136 284352 3188
rect 286784 3136 286836 3188
rect 311716 3136 311768 3188
rect 317328 3136 317380 3188
rect 348056 3272 348108 3324
rect 351736 3272 351788 3324
rect 188620 3068 188672 3120
rect 193220 3068 193272 3120
rect 239312 3068 239364 3120
rect 246304 3068 246356 3120
rect 281908 3068 281960 3120
rect 285036 3068 285088 3120
rect 336096 3068 336148 3120
rect 338764 3068 338816 3120
rect 352840 3204 352892 3256
rect 369400 3272 369452 3324
rect 380808 3272 380860 3324
rect 411904 3272 411956 3324
rect 415308 3272 415360 3324
rect 460388 3272 460440 3324
rect 481548 3272 481600 3324
rect 371700 3204 371752 3256
rect 375196 3204 375248 3256
rect 404820 3204 404872 3256
rect 416596 3204 416648 3256
rect 461584 3204 461636 3256
rect 478788 3204 478840 3256
rect 350356 3136 350408 3188
rect 370596 3136 370648 3188
rect 378048 3136 378100 3188
rect 408408 3136 408460 3188
rect 412548 3136 412600 3188
rect 456892 3136 456944 3188
rect 476028 3136 476080 3188
rect 544384 3272 544436 3324
rect 545488 3272 545540 3324
rect 547144 3204 547196 3256
rect 559748 3204 559800 3256
rect 348976 3068 349028 3120
rect 368204 3068 368256 3120
rect 372528 3068 372580 3120
rect 401324 3068 401376 3120
rect 411076 3068 411128 3120
rect 454500 3068 454552 3120
rect 470508 3068 470560 3120
rect 536104 3068 536156 3120
rect 550272 3136 550324 3188
rect 543188 3068 543240 3120
rect 57152 3000 57204 3052
rect 60832 3000 60884 3052
rect 124036 3000 124088 3052
rect 190828 3000 190880 3052
rect 191748 3000 191800 3052
rect 199108 3000 199160 3052
rect 220084 3000 220136 3052
rect 261760 3000 261812 3052
rect 267004 3000 267056 3052
rect 274824 3000 274876 3052
rect 276664 3000 276716 3052
rect 283104 3000 283156 3052
rect 284944 3000 284996 3052
rect 310428 3000 310480 3052
rect 316224 3000 316276 3052
rect 316684 3000 316736 3052
rect 323308 3000 323360 3052
rect 336004 3000 336056 3052
rect 343364 3000 343416 3052
rect 347688 3000 347740 3052
rect 367008 3000 367060 3052
rect 27712 2932 27764 2984
rect 35164 2932 35216 2984
rect 73804 2932 73856 2984
rect 74448 2932 74500 2984
rect 76196 2932 76248 2984
rect 77208 2932 77260 2984
rect 67916 2864 67968 2916
rect 129188 2932 129240 2984
rect 220452 2932 220504 2984
rect 343548 2932 343600 2984
rect 361120 2932 361172 2984
rect 366916 2932 366968 2984
rect 394240 3000 394292 3052
rect 413928 3000 413980 3052
rect 458088 3000 458140 3052
rect 466368 3000 466420 3052
rect 529020 3000 529072 3052
rect 546684 3000 546736 3052
rect 372436 2932 372488 2984
rect 400128 2932 400180 2984
rect 405648 2932 405700 2984
rect 447416 2932 447468 2984
rect 460848 2932 460900 2984
rect 521844 2932 521896 2984
rect 75000 2796 75052 2848
rect 134340 2864 134392 2916
rect 192024 2864 192076 2916
rect 219624 2864 219676 2916
rect 344928 2864 344980 2916
rect 362316 2864 362368 2916
rect 369768 2864 369820 2916
rect 396540 2864 396592 2916
rect 411168 2864 411220 2916
rect 453304 2864 453356 2916
rect 455328 2864 455380 2916
rect 514760 2864 514812 2916
rect 80888 2796 80940 2848
rect 81348 2796 81400 2848
rect 82084 2796 82136 2848
rect 139492 2796 139544 2848
rect 186136 2796 186188 2848
rect 215392 2796 215444 2848
rect 340144 2796 340196 2848
rect 354036 2796 354088 2848
rect 365628 2796 365680 2848
rect 390652 2796 390704 2848
rect 408316 2796 408368 2848
rect 450912 2796 450964 2848
rect 452568 2796 452620 2848
rect 511264 2796 511316 2848
rect 448520 2320 448572 2372
rect 449808 2320 449860 2372
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700670 73016 703520
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 105464 699718 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 170324 699718 170352 703520
rect 202800 700126 202828 703520
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 218992 700058 219020 703520
rect 218980 700052 219032 700058
rect 218980 699994 219032 700000
rect 235184 699718 235212 703520
rect 264888 700868 264940 700874
rect 264888 700810 264940 700816
rect 253848 700596 253900 700602
rect 253848 700538 253900 700544
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 7564 568880 7616 568886
rect 7564 568822 7616 568828
rect 4896 567384 4948 567390
rect 4896 567326 4948 567332
rect 4804 567248 4856 567254
rect 4804 567190 4856 567196
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 566370 3464 566879
rect 3424 566364 3476 566370
rect 3424 566306 3476 566312
rect 3792 565140 3844 565146
rect 3792 565082 3844 565088
rect 3700 564800 3752 564806
rect 3700 564742 3752 564748
rect 3608 564732 3660 564738
rect 3608 564674 3660 564680
rect 3516 564528 3568 564534
rect 3516 564470 3568 564476
rect 3424 564460 3476 564466
rect 3424 564402 3476 564408
rect 3332 554736 3384 554742
rect 3332 554678 3384 554684
rect 3344 553897 3372 554678
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3240 528556 3292 528562
rect 3240 528498 3292 528504
rect 3252 527921 3280 528498
rect 3238 527912 3294 527921
rect 3238 527847 3294 527856
rect 3240 502308 3292 502314
rect 3240 502250 3292 502256
rect 3252 501809 3280 502250
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3332 476060 3384 476066
rect 3332 476002 3384 476008
rect 3344 475697 3372 476002
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3148 358624 3200 358630
rect 3148 358566 3200 358572
rect 3160 358465 3188 358566
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 2780 254380 2832 254386
rect 2780 254322 2832 254328
rect 2792 254153 2820 254322
rect 2778 254144 2834 254153
rect 2778 254079 2834 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 2780 202768 2832 202774
rect 2780 202710 2832 202716
rect 2792 201929 2820 202710
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 58585 3464 564402
rect 3528 306241 3556 564470
rect 3620 410553 3648 564674
rect 3712 462641 3740 564742
rect 3804 514865 3832 565082
rect 3790 514856 3846 514865
rect 3790 514791 3846 514800
rect 3698 462632 3754 462641
rect 3698 462567 3754 462576
rect 3606 410544 3662 410553
rect 3606 410479 3662 410488
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 4816 202774 4844 567190
rect 4908 254386 4936 567326
rect 7576 358630 7604 568822
rect 100576 568676 100628 568682
rect 100576 568618 100628 568624
rect 14464 568608 14516 568614
rect 14464 568550 14516 568556
rect 11702 563816 11758 563825
rect 11702 563751 11758 563760
rect 7564 358624 7616 358630
rect 7564 358566 7616 358572
rect 4896 254380 4948 254386
rect 4896 254322 4948 254328
rect 4804 202768 4856 202774
rect 4804 202710 4856 202716
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 11716 137970 11744 563751
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 11704 137964 11756 137970
rect 11704 137906 11756 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 7564 135924 7616 135930
rect 7564 135866 7616 135872
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 4956 1728 4962
rect 1676 4898 1728 4904
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4898
rect 2872 4888 2924 4894
rect 2872 4830 2924 4836
rect 2884 480 2912 4830
rect 4080 480 4108 8910
rect 7576 3874 7604 135866
rect 11704 134564 11756 134570
rect 11704 134506 11756 134512
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3868 5316 3874
rect 5264 3810 5316 3816
rect 7564 3868 7616 3874
rect 7564 3810 7616 3816
rect 5276 480 5304 3810
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 8760 3256 8812 3262
rect 8760 3198 8812 3204
rect 8772 480 8800 3198
rect 9968 480 9996 3402
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 480 11192 3334
rect 11716 3262 11744 134506
rect 14476 20670 14504 568550
rect 61384 567996 61436 568002
rect 61384 567938 61436 567944
rect 57244 567792 57296 567798
rect 57244 567734 57296 567740
rect 51724 567520 51776 567526
rect 22742 567488 22798 567497
rect 51724 567462 51776 567468
rect 22742 567423 22798 567432
rect 17224 567316 17276 567322
rect 17224 567258 17276 567264
rect 17236 150414 17264 567258
rect 17224 150408 17276 150414
rect 17224 150350 17276 150356
rect 17224 136060 17276 136066
rect 17224 136002 17276 136008
rect 15844 134632 15896 134638
rect 15844 134574 15896 134580
rect 14464 20664 14516 20670
rect 14464 20606 14516 20612
rect 12348 7608 12400 7614
rect 12348 7550 12400 7556
rect 11704 3256 11756 3262
rect 11704 3198 11756 3204
rect 12360 480 12388 7550
rect 14738 3632 14794 3641
rect 14738 3567 14794 3576
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13556 480 13584 3130
rect 14752 480 14780 3567
rect 15856 3194 15884 134574
rect 17040 3528 17092 3534
rect 15934 3496 15990 3505
rect 17040 3470 17092 3476
rect 15934 3431 15990 3440
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15948 480 15976 3431
rect 17052 480 17080 3470
rect 17236 3398 17264 136002
rect 18604 135992 18656 135998
rect 18604 135934 18656 135940
rect 18236 3800 18288 3806
rect 18236 3742 18288 3748
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 18248 480 18276 3742
rect 18616 3534 18644 135934
rect 22008 135108 22060 135114
rect 22008 135050 22060 135056
rect 22020 6914 22048 135050
rect 22756 97986 22784 567423
rect 43444 566840 43496 566846
rect 43444 566782 43496 566788
rect 32404 565956 32456 565962
rect 32404 565898 32456 565904
rect 25502 563952 25558 563961
rect 25502 563887 25558 563896
rect 22744 97980 22796 97986
rect 22744 97922 22796 97928
rect 25516 85542 25544 563887
rect 32416 189038 32444 565898
rect 39302 564088 39358 564097
rect 39302 564023 39358 564032
rect 33782 563680 33838 563689
rect 33782 563615 33838 563624
rect 32404 189032 32456 189038
rect 32404 188974 32456 188980
rect 29644 136196 29696 136202
rect 29644 136138 29696 136144
rect 25504 85536 25556 85542
rect 25504 85478 25556 85484
rect 21836 6886 22048 6914
rect 20626 3768 20682 3777
rect 20626 3703 20682 3712
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19444 480 19472 3470
rect 20640 480 20668 3703
rect 21836 480 21864 6886
rect 26516 4208 26568 4214
rect 26516 4150 26568 4156
rect 23020 4004 23072 4010
rect 23020 3946 23072 3952
rect 23032 480 23060 3946
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24228 480 24256 3606
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25332 480 25360 3538
rect 26528 480 26556 4150
rect 29656 3806 29684 136138
rect 32404 136128 32456 136134
rect 32404 136070 32456 136076
rect 30104 5092 30156 5098
rect 30104 5034 30156 5040
rect 29644 3800 29696 3806
rect 29644 3742 29696 3748
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 27712 2984 27764 2990
rect 27712 2926 27764 2932
rect 27724 480 27752 2926
rect 28920 480 28948 3674
rect 30116 480 30144 5034
rect 32416 4214 32444 136070
rect 33796 6866 33824 563615
rect 35164 134768 35216 134774
rect 35164 134710 35216 134716
rect 33784 6860 33836 6866
rect 33784 6802 33836 6808
rect 32404 4208 32456 4214
rect 32404 4150 32456 4156
rect 31300 4072 31352 4078
rect 31300 4014 31352 4020
rect 31312 480 31340 4014
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32416 480 32444 3742
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33612 480 33640 3334
rect 34796 3120 34848 3126
rect 34796 3062 34848 3068
rect 34808 480 34836 3062
rect 35176 2990 35204 134710
rect 37188 134700 37240 134706
rect 37188 134642 37240 134648
rect 35256 26920 35308 26926
rect 35256 26862 35308 26868
rect 35268 3398 35296 26862
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 35256 3392 35308 3398
rect 35256 3334 35308 3340
rect 35164 2984 35216 2990
rect 35164 2926 35216 2932
rect 36004 480 36032 3878
rect 37200 480 37228 134642
rect 39316 45558 39344 564023
rect 43456 528562 43484 566782
rect 50344 565888 50396 565894
rect 50344 565830 50396 565836
rect 47584 565004 47636 565010
rect 47584 564946 47636 564952
rect 43444 528556 43496 528562
rect 43444 528498 43496 528504
rect 47596 241466 47624 564946
rect 47584 241460 47636 241466
rect 47584 241402 47636 241408
rect 47584 135652 47636 135658
rect 47584 135594 47636 135600
rect 43444 135176 43496 135182
rect 43444 135118 43496 135124
rect 41328 134904 41380 134910
rect 41328 134846 41380 134852
rect 39396 134836 39448 134842
rect 39396 134778 39448 134784
rect 39304 45552 39356 45558
rect 39304 45494 39356 45500
rect 39408 4078 39436 134778
rect 39396 4072 39448 4078
rect 39396 4014 39448 4020
rect 39580 3868 39632 3874
rect 39580 3810 39632 3816
rect 38384 3256 38436 3262
rect 38384 3198 38436 3204
rect 38396 480 38424 3198
rect 39592 480 39620 3810
rect 41340 3398 41368 134846
rect 41880 4140 41932 4146
rect 41880 4082 41932 4088
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 40696 480 40724 3334
rect 41892 480 41920 4082
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 43088 480 43116 4014
rect 43456 4010 43484 135118
rect 44272 5228 44324 5234
rect 44272 5170 44324 5176
rect 43444 4004 43496 4010
rect 43444 3946 43496 3952
rect 44284 480 44312 5170
rect 47596 5098 47624 135594
rect 50356 33114 50384 565830
rect 51736 293962 51764 567462
rect 53104 566704 53156 566710
rect 53104 566646 53156 566652
rect 53116 449886 53144 566646
rect 54484 566432 54536 566438
rect 54484 566374 54536 566380
rect 53104 449880 53156 449886
rect 53104 449822 53156 449828
rect 54496 346390 54524 566374
rect 57256 398818 57284 567734
rect 58624 566024 58676 566030
rect 58624 565966 58676 565972
rect 57244 398812 57296 398818
rect 57244 398754 57296 398760
rect 54484 346384 54536 346390
rect 54484 346326 54536 346332
rect 51724 293956 51776 293962
rect 51724 293898 51776 293904
rect 54484 136604 54536 136610
rect 54484 136546 54536 136552
rect 51724 136264 51776 136270
rect 51724 136206 51776 136212
rect 50344 33108 50396 33114
rect 50344 33050 50396 33056
rect 50436 32428 50488 32434
rect 50436 32370 50488 32376
rect 47584 5092 47636 5098
rect 47584 5034 47636 5040
rect 47860 5092 47912 5098
rect 47860 5034 47912 5040
rect 46664 4004 46716 4010
rect 46664 3946 46716 3952
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45480 480 45508 3334
rect 46676 480 46704 3946
rect 47872 480 47900 5034
rect 48964 4208 49016 4214
rect 48964 4150 49016 4156
rect 48976 480 49004 4150
rect 50448 3262 50476 32370
rect 51356 5160 51408 5166
rect 51356 5102 51408 5108
rect 50436 3256 50488 3262
rect 50436 3198 50488 3204
rect 50160 3120 50212 3126
rect 50160 3062 50212 3068
rect 50172 480 50200 3062
rect 51368 480 51396 5102
rect 51736 4214 51764 136206
rect 53748 135040 53800 135046
rect 53748 134982 53800 134988
rect 51724 4208 51776 4214
rect 51724 4150 51776 4156
rect 53760 3330 53788 134982
rect 54496 5234 54524 136546
rect 57244 133204 57296 133210
rect 57244 133146 57296 133152
rect 57256 6914 57284 133146
rect 58636 111790 58664 565966
rect 61396 502314 61424 567938
rect 79324 566976 79376 566982
rect 79324 566918 79376 566924
rect 65524 566908 65576 566914
rect 65524 566850 65576 566856
rect 61384 502308 61436 502314
rect 61384 502250 61436 502256
rect 65536 476066 65564 566850
rect 75184 566772 75236 566778
rect 75184 566714 75236 566720
rect 68284 566296 68336 566302
rect 68284 566238 68336 566244
rect 65524 476060 65576 476066
rect 65524 476002 65576 476008
rect 68296 164218 68324 566238
rect 71044 565684 71096 565690
rect 71044 565626 71096 565632
rect 69664 564664 69716 564670
rect 69664 564606 69716 564612
rect 68284 164212 68336 164218
rect 68284 164154 68336 164160
rect 68284 136536 68336 136542
rect 68284 136478 68336 136484
rect 65524 135788 65576 135794
rect 65524 135730 65576 135736
rect 62028 134972 62080 134978
rect 62028 134914 62080 134920
rect 58624 111784 58676 111790
rect 58624 111726 58676 111732
rect 57164 6886 57284 6914
rect 56048 5364 56100 5370
rect 56048 5306 56100 5312
rect 54484 5228 54536 5234
rect 54484 5170 54536 5176
rect 54944 5228 54996 5234
rect 54944 5170 54996 5176
rect 52552 3324 52604 3330
rect 52552 3266 52604 3272
rect 53748 3324 53800 3330
rect 53748 3266 53800 3272
rect 52564 480 52592 3266
rect 53748 3188 53800 3194
rect 53748 3130 53800 3136
rect 53760 480 53788 3130
rect 54956 480 54984 5170
rect 56060 480 56088 5306
rect 57164 3058 57192 6886
rect 59636 5500 59688 5506
rect 59636 5442 59688 5448
rect 58440 5296 58492 5302
rect 58440 5238 58492 5244
rect 57244 3188 57296 3194
rect 57244 3130 57296 3136
rect 57152 3052 57204 3058
rect 57152 2994 57204 3000
rect 57256 480 57284 3130
rect 58452 480 58480 5238
rect 59648 480 59676 5442
rect 60832 3052 60884 3058
rect 60832 2994 60884 3000
rect 60844 480 60872 2994
rect 62040 480 62068 134914
rect 65536 5370 65564 135730
rect 65616 5432 65668 5438
rect 65616 5374 65668 5380
rect 65524 5364 65576 5370
rect 65524 5306 65576 5312
rect 63224 4752 63276 4758
rect 63224 4694 63276 4700
rect 63236 480 63264 4694
rect 64328 3120 64380 3126
rect 64328 3062 64380 3068
rect 64340 480 64368 3062
rect 65628 2802 65656 5374
rect 66720 5364 66772 5370
rect 66720 5306 66772 5312
rect 65536 2774 65656 2802
rect 65536 480 65564 2774
rect 66732 480 66760 5306
rect 68296 4758 68324 136478
rect 69676 71738 69704 564606
rect 71056 554742 71084 565626
rect 72424 565276 72476 565282
rect 72424 565218 72476 565224
rect 71044 554736 71096 554742
rect 71044 554678 71096 554684
rect 72436 215286 72464 565218
rect 75196 372570 75224 566714
rect 76564 566568 76616 566574
rect 76564 566510 76616 566516
rect 75184 372564 75236 372570
rect 75184 372506 75236 372512
rect 76576 267714 76604 566510
rect 77944 565548 77996 565554
rect 77944 565490 77996 565496
rect 77956 320142 77984 565490
rect 79336 423638 79364 566918
rect 100588 565298 100616 568618
rect 106200 568206 106228 699654
rect 152740 569016 152792 569022
rect 152740 568958 152792 568964
rect 130384 568948 130436 568954
rect 130384 568890 130436 568896
rect 119160 568812 119212 568818
rect 119160 568754 119212 568760
rect 111708 568744 111760 568750
rect 111708 568686 111760 568692
rect 106188 568200 106240 568206
rect 106188 568142 106240 568148
rect 104256 566092 104308 566098
rect 104256 566034 104308 566040
rect 104268 565298 104296 566034
rect 111720 565298 111748 568686
rect 119172 565298 119200 568754
rect 122746 567352 122802 567361
rect 122746 567287 122802 567296
rect 122760 565298 122788 567287
rect 126612 566228 126664 566234
rect 126612 566170 126664 566176
rect 126624 565298 126652 566170
rect 130396 565298 130424 568890
rect 145288 567588 145340 567594
rect 145288 567530 145340 567536
rect 133788 567452 133840 567458
rect 133788 567394 133840 567400
rect 133800 565570 133828 567394
rect 100280 565270 100616 565298
rect 103960 565270 104296 565298
rect 111412 565270 111748 565298
rect 118864 565270 119200 565298
rect 122636 565270 122788 565298
rect 126316 565270 126652 565298
rect 130088 565270 130424 565298
rect 133754 565542 133828 565570
rect 133754 565284 133782 565542
rect 145300 565298 145328 567530
rect 148968 566160 149020 566166
rect 148968 566102 149020 566108
rect 148980 565298 149008 566102
rect 152752 565298 152780 568958
rect 171060 568342 171088 699654
rect 231768 643136 231820 643142
rect 231768 643078 231820 643084
rect 227628 616888 227680 616894
rect 227628 616830 227680 616836
rect 219348 590708 219400 590714
rect 219348 590650 219400 590656
rect 175096 569084 175148 569090
rect 175096 569026 175148 569032
rect 171048 568336 171100 568342
rect 171048 568278 171100 568284
rect 167644 567724 167696 567730
rect 167644 567666 167696 567672
rect 156420 567656 156472 567662
rect 156420 567598 156472 567604
rect 156432 565298 156460 567598
rect 160008 565344 160060 565350
rect 144992 565270 145328 565298
rect 148672 565270 149008 565298
rect 152444 565270 152780 565298
rect 156124 565270 156460 565298
rect 159896 565292 160008 565298
rect 167656 565298 167684 567666
rect 170956 566500 171008 566506
rect 170956 566442 171008 566448
rect 159896 565286 160060 565292
rect 159896 565270 160048 565286
rect 167348 565270 167684 565298
rect 170968 565162 170996 566442
rect 175108 565298 175136 569026
rect 189908 567928 189960 567934
rect 189908 567870 189960 567876
rect 178776 567860 178828 567866
rect 178776 567802 178828 567808
rect 178788 565298 178816 567802
rect 182226 565480 182278 565486
rect 182226 565422 182278 565428
rect 174800 565270 175136 565298
rect 178480 565270 178816 565298
rect 182238 565284 182266 565422
rect 189920 565298 189948 567870
rect 204812 567112 204864 567118
rect 204812 567054 204864 567060
rect 193680 567044 193732 567050
rect 193680 566986 193732 566992
rect 193692 565298 193720 566986
rect 197268 566636 197320 566642
rect 197268 566578 197320 566584
rect 197280 565298 197308 566578
rect 204824 565298 204852 567054
rect 208216 565616 208268 565622
rect 208216 565558 208268 565564
rect 189612 565270 189948 565298
rect 193384 565270 193720 565298
rect 197064 565270 197308 565298
rect 204516 565270 204852 565298
rect 201132 565208 201184 565214
rect 170968 565134 171028 565162
rect 200836 565156 201132 565162
rect 200836 565150 201184 565156
rect 208228 565162 208256 565558
rect 211942 565412 211994 565418
rect 211942 565354 211994 565360
rect 211954 565284 211982 565354
rect 219360 565298 219388 590650
rect 223488 576904 223540 576910
rect 223488 576846 223540 576852
rect 223500 565298 223528 576846
rect 227640 568546 227668 616830
rect 231780 568546 231808 643078
rect 234528 630692 234580 630698
rect 234528 630634 234580 630640
rect 227168 568540 227220 568546
rect 227168 568482 227220 568488
rect 227628 568540 227680 568546
rect 227628 568482 227680 568488
rect 230940 568540 230992 568546
rect 230940 568482 230992 568488
rect 231768 568540 231820 568546
rect 231768 568482 231820 568488
rect 227180 565298 227208 568482
rect 230952 565298 230980 568482
rect 234540 565298 234568 630634
rect 235920 568478 235948 699654
rect 242808 696992 242860 696998
rect 242808 696934 242860 696940
rect 238668 670812 238720 670818
rect 238668 670754 238720 670760
rect 235908 568472 235960 568478
rect 235908 568414 235960 568420
rect 238680 567194 238708 670754
rect 242820 568546 242848 696934
rect 245568 683256 245620 683262
rect 245568 683198 245620 683204
rect 242072 568540 242124 568546
rect 242072 568482 242124 568488
rect 242808 568540 242860 568546
rect 242808 568482 242860 568488
rect 238496 567166 238708 567194
rect 238496 565298 238524 567166
rect 242084 565298 242112 568482
rect 245580 565570 245608 683198
rect 253860 568546 253888 700538
rect 256608 700528 256660 700534
rect 256608 700470 256660 700476
rect 253296 568540 253348 568546
rect 253296 568482 253348 568488
rect 253848 568540 253900 568546
rect 253848 568482 253900 568488
rect 249524 568064 249576 568070
rect 249524 568006 249576 568012
rect 219360 565270 219420 565298
rect 223192 565270 223528 565298
rect 226872 565270 227208 565298
rect 230644 565270 230980 565298
rect 234324 565270 234568 565298
rect 238096 565270 238524 565298
rect 241776 565270 242112 565298
rect 245534 565542 245608 565570
rect 245534 565284 245562 565542
rect 249536 565298 249564 568006
rect 253308 565298 253336 568482
rect 249228 565270 249564 565298
rect 253000 565270 253336 565298
rect 256620 565298 256648 700470
rect 264900 568546 264928 700810
rect 267660 699854 267688 703520
rect 269028 700800 269080 700806
rect 269028 700742 269080 700748
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 269040 568546 269068 700742
rect 280068 700256 280120 700262
rect 280068 700198 280120 700204
rect 275928 700188 275980 700194
rect 275928 700130 275980 700136
rect 264428 568540 264480 568546
rect 264428 568482 264480 568488
rect 264888 568540 264940 568546
rect 264888 568482 264940 568488
rect 268200 568540 268252 568546
rect 268200 568482 268252 568488
rect 269028 568540 269080 568546
rect 269028 568482 269080 568488
rect 260564 568132 260616 568138
rect 260564 568074 260616 568080
rect 260576 565298 260604 568074
rect 264440 565298 264468 568482
rect 268212 565298 268240 568482
rect 271788 568268 271840 568274
rect 271788 568210 271840 568216
rect 271800 565298 271828 568210
rect 275940 567194 275968 700130
rect 280080 568546 280108 700198
rect 283852 699786 283880 703520
rect 291108 699984 291160 699990
rect 291108 699926 291160 699932
rect 286968 699916 287020 699922
rect 286968 699858 287020 699864
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 279332 568540 279384 568546
rect 279332 568482 279384 568488
rect 280068 568540 280120 568546
rect 280068 568482 280120 568488
rect 275756 567166 275968 567194
rect 275756 565298 275784 567166
rect 279344 565298 279372 568482
rect 282828 568404 282880 568410
rect 282828 568346 282880 568352
rect 282840 565570 282868 568346
rect 286980 567194 287008 699858
rect 291120 568546 291148 699926
rect 296720 699848 296772 699854
rect 296720 699790 296772 699796
rect 296732 576854 296760 699790
rect 296732 576826 297220 576854
rect 290556 568540 290608 568546
rect 290556 568482 290608 568488
rect 291108 568540 291160 568546
rect 291108 568482 291160 568488
rect 293868 568540 293920 568546
rect 293868 568482 293920 568488
rect 256620 565270 256680 565298
rect 260452 565270 260604 565298
rect 264132 565270 264468 565298
rect 267904 565270 268240 565298
rect 271584 565270 271828 565298
rect 275356 565270 275784 565298
rect 279036 565270 279372 565298
rect 282794 565542 282868 565570
rect 286888 567166 287008 567194
rect 282794 565284 282822 565542
rect 286888 565298 286916 567166
rect 290568 565298 290596 568482
rect 286488 565270 286916 565298
rect 290260 565270 290596 565298
rect 293880 565298 293908 568482
rect 297192 565298 297220 576826
rect 299492 568546 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 322940 701004 322992 701010
rect 322940 700946 322992 700952
rect 318800 700936 318852 700942
rect 318800 700878 318852 700884
rect 307760 700120 307812 700126
rect 307760 700062 307812 700068
rect 300860 699780 300912 699786
rect 300860 699722 300912 699728
rect 300872 576854 300900 699722
rect 307772 576854 307800 700062
rect 311900 700052 311952 700058
rect 311900 699994 311952 700000
rect 311912 576854 311940 699994
rect 318812 576854 318840 700878
rect 322952 576854 322980 700946
rect 329840 700664 329892 700670
rect 329840 700606 329892 700612
rect 329852 576854 329880 700606
rect 332520 699922 332548 703520
rect 333980 700732 334032 700738
rect 333980 700674 334032 700680
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 333992 576854 334020 700674
rect 338120 700460 338172 700466
rect 338120 700402 338172 700408
rect 338132 576854 338160 700402
rect 345020 700392 345072 700398
rect 345020 700334 345072 700340
rect 342260 700324 342312 700330
rect 342260 700266 342312 700272
rect 300872 576826 300992 576854
rect 307772 576826 308444 576854
rect 311912 576826 312124 576854
rect 318812 576826 319576 576854
rect 322952 576826 323348 576854
rect 329852 576826 330800 576854
rect 333992 576826 334480 576854
rect 338132 576826 338252 576854
rect 299480 568540 299532 568546
rect 299480 568482 299532 568488
rect 300964 565298 300992 576826
rect 305000 568472 305052 568478
rect 305000 568414 305052 568420
rect 305012 565298 305040 568414
rect 308416 565298 308444 576826
rect 312096 565298 312124 576826
rect 316040 568336 316092 568342
rect 316040 568278 316092 568284
rect 316052 565298 316080 568278
rect 319548 565298 319576 576826
rect 323320 565298 323348 576826
rect 327080 568200 327132 568206
rect 327080 568142 327132 568148
rect 327092 565298 327120 568142
rect 330772 565298 330800 576826
rect 334452 565298 334480 576826
rect 338224 565298 338252 576826
rect 342272 565298 342300 700266
rect 345032 576854 345060 700334
rect 348804 699990 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 349160 683188 349212 683194
rect 349160 683130 349212 683136
rect 349172 576854 349200 683130
rect 356060 670744 356112 670750
rect 356060 670686 356112 670692
rect 353300 656940 353352 656946
rect 353300 656882 353352 656888
rect 345032 576826 345704 576854
rect 349172 576826 349384 576854
rect 345676 565298 345704 576826
rect 349356 565298 349384 576826
rect 353312 565298 353340 656882
rect 356072 576854 356100 670686
rect 360200 632120 360252 632126
rect 360200 632062 360252 632068
rect 360212 576854 360240 632062
rect 356072 576826 356836 576854
rect 360212 576826 360608 576854
rect 356808 565298 356836 576826
rect 360580 565298 360608 576826
rect 364352 568410 364380 702406
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 367100 618316 367152 618322
rect 367100 618258 367152 618264
rect 364432 605872 364484 605878
rect 364432 605814 364484 605820
rect 364340 568404 364392 568410
rect 364340 568346 364392 568352
rect 364444 565298 364472 605814
rect 367112 576854 367140 618258
rect 371240 579692 371292 579698
rect 371240 579634 371292 579640
rect 371252 576854 371280 579634
rect 367112 576826 368060 576854
rect 371252 576826 371740 576854
rect 368032 565298 368060 576826
rect 371712 565298 371740 576826
rect 423956 568880 424008 568886
rect 423956 568822 424008 568828
rect 386696 567996 386748 568002
rect 386696 567938 386748 567944
rect 383016 566840 383068 566846
rect 383016 566782 383068 566788
rect 379520 566364 379572 566370
rect 379520 566306 379572 566312
rect 375564 565684 375616 565690
rect 375564 565626 375616 565632
rect 375576 565298 375604 565626
rect 379532 565298 379560 566306
rect 383028 565298 383056 566782
rect 386708 565298 386736 567938
rect 409052 567792 409104 567798
rect 409052 567734 409104 567740
rect 405280 566976 405332 566982
rect 405280 566918 405332 566924
rect 394148 566908 394200 566914
rect 394148 566850 394200 566856
rect 394160 565298 394188 566850
rect 397920 566704 397972 566710
rect 397920 566646 397972 566652
rect 397932 565298 397960 566646
rect 405292 565298 405320 566918
rect 409064 565298 409092 567734
rect 416780 566772 416832 566778
rect 416780 566714 416832 566720
rect 416792 565298 416820 566714
rect 420184 566432 420236 566438
rect 420184 566374 420236 566380
rect 420196 565298 420224 566374
rect 423968 565298 423996 568822
rect 429212 568274 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 429200 568268 429252 568274
rect 429200 568210 429252 568216
rect 494072 568138 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 556804 569084 556856 569090
rect 556804 569026 556856 569032
rect 547144 569016 547196 569022
rect 547144 568958 547196 568964
rect 543004 568948 543056 568954
rect 543004 568890 543056 568896
rect 540244 568812 540296 568818
rect 540244 568754 540296 568760
rect 502432 568608 502484 568614
rect 502432 568550 502484 568556
rect 494060 568132 494112 568138
rect 494060 568074 494112 568080
rect 431408 567520 431460 567526
rect 431408 567462 431460 567468
rect 479798 567488 479854 567497
rect 427958 565548 428010 565554
rect 427958 565490 428010 565496
rect 293880 565270 293940 565298
rect 297192 565270 297620 565298
rect 300964 565270 301392 565298
rect 305012 565270 305072 565298
rect 308416 565270 308844 565298
rect 312096 565270 312524 565298
rect 316052 565270 316296 565298
rect 319548 565270 319976 565298
rect 323320 565270 323748 565298
rect 327092 565270 327428 565298
rect 330772 565270 331200 565298
rect 334452 565270 334880 565298
rect 338224 565270 338652 565298
rect 342272 565270 342332 565298
rect 345676 565270 346104 565298
rect 349356 565270 349784 565298
rect 353312 565270 353556 565298
rect 356808 565270 357236 565298
rect 360580 565270 361008 565298
rect 364444 565270 364688 565298
rect 368032 565270 368460 565298
rect 371712 565270 372140 565298
rect 375576 565270 375912 565298
rect 379532 565270 379592 565298
rect 383028 565270 383364 565298
rect 386708 565270 387044 565298
rect 394160 565270 394496 565298
rect 397932 565270 398268 565298
rect 405292 565270 405628 565298
rect 409064 565270 409400 565298
rect 416792 565270 416852 565298
rect 420196 565270 420532 565298
rect 423968 565270 424304 565298
rect 427970 565284 427998 565490
rect 431420 565298 431448 567462
rect 479798 567423 479854 567432
rect 446312 567384 446364 567390
rect 446312 567326 446364 567332
rect 438860 566568 438912 566574
rect 438860 566510 438912 566516
rect 438872 565298 438900 566510
rect 446324 565298 446352 567326
rect 468668 567316 468720 567322
rect 468668 567258 468720 567264
rect 457444 567248 457496 567254
rect 457444 567190 457496 567196
rect 454040 565956 454092 565962
rect 454040 565898 454092 565904
rect 454052 565298 454080 565898
rect 457456 565298 457484 567190
rect 461216 566296 461268 566302
rect 461216 566238 461268 566244
rect 461228 565298 461256 566238
rect 468680 565298 468708 567258
rect 472348 566024 472400 566030
rect 472348 565966 472400 565972
rect 472360 565298 472388 565966
rect 479812 565298 479840 567423
rect 494704 565888 494756 565894
rect 494704 565830 494756 565836
rect 494716 565298 494744 565830
rect 502444 565298 502472 568550
rect 525064 567928 525116 567934
rect 525064 567870 525116 567876
rect 522304 567860 522356 567866
rect 522304 567802 522356 567808
rect 520924 567724 520976 567730
rect 520924 567666 520976 567672
rect 519544 567656 519596 567662
rect 519544 567598 519596 567604
rect 518164 567588 518216 567594
rect 518164 567530 518216 567536
rect 515404 567452 515456 567458
rect 515404 567394 515456 567400
rect 512642 567352 512698 567361
rect 512642 567287 512698 567296
rect 507124 567112 507176 567118
rect 507124 567054 507176 567060
rect 505744 567044 505796 567050
rect 505744 566986 505796 566992
rect 431420 565270 431756 565298
rect 438872 565270 439208 565298
rect 446324 565270 446660 565298
rect 450004 565282 450340 565298
rect 449992 565276 450340 565282
rect 450044 565270 450340 565276
rect 454052 565270 454112 565298
rect 457456 565270 457792 565298
rect 461228 565270 461564 565298
rect 468680 565270 469016 565298
rect 472360 565270 472696 565298
rect 479812 565270 480148 565298
rect 494716 565270 495052 565298
rect 502444 565270 502504 565298
rect 449992 565218 450044 565224
rect 200836 565134 201172 565150
rect 208228 565134 208288 565162
rect 390572 565146 390816 565162
rect 390560 565140 390816 565146
rect 390612 565134 390816 565140
rect 390560 565082 390612 565088
rect 137836 565072 137888 565078
rect 137540 565020 137836 565026
rect 137540 565014 137888 565020
rect 137540 564998 137876 565014
rect 442552 565010 442888 565026
rect 442540 565004 442888 565010
rect 442592 564998 442888 565004
rect 442540 564946 442592 564952
rect 186228 564936 186280 564942
rect 115184 564874 115520 564890
rect 185932 564884 186228 564890
rect 185932 564878 186280 564884
rect 115184 564868 115532 564874
rect 115184 564862 115480 564868
rect 185932 564862 186268 564878
rect 115480 564810 115532 564816
rect 401600 564800 401652 564806
rect 401652 564748 401948 564754
rect 401600 564742 401948 564748
rect 401612 564726 401948 564742
rect 412836 564738 413080 564754
rect 435100 564738 435436 564754
rect 412824 564732 413080 564738
rect 412876 564726 413080 564732
rect 435088 564732 435436 564738
rect 412824 564674 412876 564680
rect 435140 564726 435436 564732
rect 435088 564674 435140 564680
rect 483572 564664 483624 564670
rect 81990 564632 82046 564641
rect 81696 564590 81990 564618
rect 81990 564567 82046 564576
rect 85026 564632 85082 564641
rect 89350 564632 89406 564641
rect 85082 564590 85376 564618
rect 89056 564590 89350 564618
rect 85026 564567 85082 564576
rect 93122 564632 93178 564641
rect 92828 564590 93122 564618
rect 89350 564567 89406 564576
rect 93122 564567 93178 564576
rect 96342 564632 96398 564641
rect 141514 564632 141570 564641
rect 96398 564590 96508 564618
rect 107732 564602 108068 564618
rect 107732 564596 108080 564602
rect 107732 564590 108028 564596
rect 96342 564567 96398 564576
rect 141220 564590 141514 564618
rect 163778 564632 163834 564641
rect 163576 564590 163778 564618
rect 141514 564567 141570 564576
rect 216034 564632 216090 564641
rect 215740 564590 216034 564618
rect 163778 564567 163834 564576
rect 216034 564567 216090 564576
rect 465078 564632 465134 564641
rect 476118 564632 476174 564641
rect 465134 564590 465244 564618
rect 465078 564567 465134 564576
rect 476174 564590 476468 564618
rect 487342 564632 487398 564641
rect 483624 564612 483920 564618
rect 483572 564606 483920 564612
rect 483584 564590 483920 564606
rect 476118 564567 476174 564576
rect 498566 564632 498622 564641
rect 487398 564590 487600 564618
rect 491220 564602 491372 564618
rect 491208 564596 491372 564602
rect 487342 564567 487398 564576
rect 108028 564538 108080 564544
rect 491260 564590 491372 564596
rect 498622 564590 498824 564618
rect 498566 564567 498622 564576
rect 491208 564538 491260 564544
rect 505756 458182 505784 566986
rect 507136 511970 507164 567054
rect 508504 566092 508556 566098
rect 508504 566034 508556 566040
rect 507124 511964 507176 511970
rect 507124 511906 507176 511912
rect 505744 458176 505796 458182
rect 505744 458118 505796 458124
rect 79324 423632 79376 423638
rect 79324 423574 79376 423580
rect 77944 320136 77996 320142
rect 77944 320078 77996 320084
rect 76564 267708 76616 267714
rect 76564 267650 76616 267656
rect 72424 215280 72476 215286
rect 72424 215222 72476 215228
rect 80164 138638 80224 138666
rect 80060 138440 80112 138446
rect 80060 138382 80112 138388
rect 74448 136468 74500 136474
rect 74448 136410 74500 136416
rect 71688 136332 71740 136338
rect 71688 136274 71740 136280
rect 69664 71732 69716 71738
rect 69664 71674 69716 71680
rect 70308 71052 70360 71058
rect 70308 70994 70360 71000
rect 69112 6180 69164 6186
rect 69112 6122 69164 6128
rect 68284 4752 68336 4758
rect 68284 4694 68336 4700
rect 67916 2916 67968 2922
rect 67916 2858 67968 2864
rect 67928 480 67956 2858
rect 69124 480 69152 6122
rect 70320 480 70348 70994
rect 71700 6914 71728 136274
rect 72424 135584 72476 135590
rect 72424 135526 72476 135532
rect 71516 6886 71728 6914
rect 71516 480 71544 6886
rect 72436 5506 72464 135526
rect 72424 5500 72476 5506
rect 72424 5442 72476 5448
rect 72608 5500 72660 5506
rect 72608 5442 72660 5448
rect 72620 480 72648 5442
rect 74460 2990 74488 136410
rect 78496 136400 78548 136406
rect 78496 136342 78548 136348
rect 75184 135516 75236 135522
rect 75184 135458 75236 135464
rect 75196 8974 75224 135458
rect 76932 135448 76984 135454
rect 76932 135390 76984 135396
rect 76944 135114 76972 135390
rect 76932 135108 76984 135114
rect 76932 135050 76984 135056
rect 77208 135108 77260 135114
rect 77208 135050 77260 135056
rect 75184 8968 75236 8974
rect 75184 8910 75236 8916
rect 77220 2990 77248 135050
rect 78508 16574 78536 136342
rect 79324 135380 79376 135386
rect 79324 135322 79376 135328
rect 78508 16546 78628 16574
rect 77392 4684 77444 4690
rect 77392 4626 77444 4632
rect 73804 2984 73856 2990
rect 73804 2926 73856 2932
rect 74448 2984 74500 2990
rect 74448 2926 74500 2932
rect 76196 2984 76248 2990
rect 76196 2926 76248 2932
rect 77208 2984 77260 2990
rect 77208 2926 77260 2932
rect 73816 480 73844 2926
rect 75000 2848 75052 2854
rect 75000 2790 75052 2796
rect 75012 480 75040 2790
rect 76208 480 76236 2926
rect 77404 480 77432 4626
rect 78600 480 78628 16546
rect 79336 7614 79364 135322
rect 79324 7608 79376 7614
rect 79324 7550 79376 7556
rect 80072 4962 80100 138382
rect 80060 4956 80112 4962
rect 80060 4898 80112 4904
rect 80164 4826 80192 138638
rect 81038 138446 81066 138652
rect 81026 138440 81078 138446
rect 81866 138394 81894 138652
rect 82786 138394 82814 138652
rect 83614 138394 83642 138652
rect 84442 138394 84470 138652
rect 85362 138394 85390 138652
rect 86190 138394 86218 138652
rect 81026 138382 81078 138388
rect 81820 138366 81894 138394
rect 82740 138366 82814 138394
rect 83568 138366 83642 138394
rect 84396 138366 84470 138394
rect 85316 138366 85390 138394
rect 86144 138366 86218 138394
rect 87018 138394 87046 138652
rect 87938 138394 87966 138652
rect 88766 138394 88794 138652
rect 89594 138394 89622 138652
rect 90514 138394 90542 138652
rect 91342 138394 91370 138652
rect 92262 138394 92290 138652
rect 93090 138394 93118 138652
rect 87018 138366 87092 138394
rect 81348 135856 81400 135862
rect 81348 135798 81400 135804
rect 80152 4820 80204 4826
rect 80152 4762 80204 4768
rect 79692 4752 79744 4758
rect 79692 4694 79744 4700
rect 79704 480 79732 4694
rect 81360 2854 81388 135798
rect 81820 4894 81848 138366
rect 82740 135522 82768 138366
rect 83568 135930 83596 138366
rect 83556 135924 83608 135930
rect 83556 135866 83608 135872
rect 82728 135516 82780 135522
rect 82728 135458 82780 135464
rect 83464 135516 83516 135522
rect 83464 135458 83516 135464
rect 83280 8968 83332 8974
rect 83280 8910 83332 8916
rect 81808 4888 81860 4894
rect 81808 4830 81860 4836
rect 80888 2848 80940 2854
rect 80888 2790 80940 2796
rect 81348 2848 81400 2854
rect 81348 2790 81400 2796
rect 82084 2848 82136 2854
rect 82084 2790 82136 2796
rect 80900 480 80928 2790
rect 82096 480 82124 2790
rect 83292 480 83320 8910
rect 83476 6186 83504 135458
rect 83464 6180 83516 6186
rect 83464 6122 83516 6128
rect 84396 3369 84424 138366
rect 85316 5030 85344 138366
rect 86144 134570 86172 138366
rect 86868 135720 86920 135726
rect 86868 135662 86920 135668
rect 86132 134564 86184 134570
rect 86132 134506 86184 134512
rect 86880 6914 86908 135662
rect 86696 6886 86908 6914
rect 85304 5024 85356 5030
rect 85304 4966 85356 4972
rect 84476 4820 84528 4826
rect 84476 4762 84528 4768
rect 84382 3360 84438 3369
rect 84382 3295 84438 3304
rect 84488 480 84516 4762
rect 86696 3534 86724 6886
rect 86868 6180 86920 6186
rect 86868 6122 86920 6128
rect 85672 3528 85724 3534
rect 85672 3470 85724 3476
rect 86684 3528 86736 3534
rect 86684 3470 86736 3476
rect 85684 480 85712 3470
rect 86880 480 86908 6122
rect 87064 4214 87092 138366
rect 87892 138366 87966 138394
rect 88720 138366 88794 138394
rect 89548 138366 89622 138394
rect 90468 138366 90542 138394
rect 91296 138366 91370 138394
rect 92216 138366 92290 138394
rect 93044 138366 93118 138394
rect 93918 138394 93946 138652
rect 94838 138394 94866 138652
rect 95666 138394 95694 138652
rect 96494 138394 96522 138652
rect 97414 138394 97442 138652
rect 98242 138394 98270 138652
rect 99070 138394 99098 138652
rect 99990 138394 100018 138652
rect 100818 138394 100846 138652
rect 101738 138394 101766 138652
rect 102566 138394 102594 138652
rect 103394 138394 103422 138652
rect 104314 138394 104342 138652
rect 105142 138394 105170 138652
rect 105970 138394 105998 138652
rect 106890 138394 106918 138652
rect 107718 138394 107746 138652
rect 108546 138394 108574 138652
rect 109466 138394 109494 138652
rect 110294 138394 110322 138652
rect 111122 138394 111150 138652
rect 112042 138394 112070 138652
rect 112870 138394 112898 138652
rect 113790 138394 113818 138652
rect 114618 138394 114646 138652
rect 115446 138394 115474 138652
rect 116366 138394 116394 138652
rect 117194 138394 117222 138652
rect 118022 138394 118050 138652
rect 118942 138394 118970 138652
rect 119770 138394 119798 138652
rect 120598 138394 120626 138652
rect 93918 138366 94084 138394
rect 87892 136066 87920 138366
rect 87880 136060 87932 136066
rect 87880 136002 87932 136008
rect 88248 135924 88300 135930
rect 88248 135866 88300 135872
rect 88260 6914 88288 135866
rect 88720 135386 88748 138366
rect 88708 135380 88760 135386
rect 88708 135322 88760 135328
rect 89548 134638 89576 138366
rect 89536 134632 89588 134638
rect 89536 134574 89588 134580
rect 87984 6886 88288 6914
rect 87052 4208 87104 4214
rect 87052 4150 87104 4156
rect 87984 480 88012 6886
rect 90468 3641 90496 138366
rect 91008 134564 91060 134570
rect 91008 134506 91060 134512
rect 90454 3632 90510 3641
rect 90454 3567 90510 3576
rect 91020 3534 91048 134506
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91296 3505 91324 138366
rect 92216 135998 92244 138366
rect 93044 136202 93072 138366
rect 93032 136196 93084 136202
rect 93032 136138 93084 136144
rect 93768 136060 93820 136066
rect 93768 136002 93820 136008
rect 92204 135992 92256 135998
rect 92204 135934 92256 135940
rect 91560 4888 91612 4894
rect 91560 4830 91612 4836
rect 91008 3470 91060 3476
rect 91282 3496 91338 3505
rect 89168 3460 89220 3466
rect 89168 3402 89220 3408
rect 89180 480 89208 3402
rect 90376 480 90404 3470
rect 91282 3431 91338 3440
rect 91572 480 91600 4830
rect 93780 3534 93808 136002
rect 93952 4956 94004 4962
rect 93952 4898 94004 4904
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 92768 480 92796 3470
rect 93964 480 93992 4898
rect 94056 4214 94084 138366
rect 94792 138366 94866 138394
rect 95620 138366 95694 138394
rect 96448 138366 96522 138394
rect 97368 138366 97442 138394
rect 98196 138366 98270 138394
rect 99024 138366 99098 138394
rect 99944 138366 100018 138394
rect 100772 138366 100846 138394
rect 101692 138366 101766 138394
rect 102520 138366 102594 138394
rect 103348 138366 103422 138394
rect 104268 138366 104342 138394
rect 105096 138366 105170 138394
rect 105924 138366 105998 138394
rect 106844 138366 106918 138394
rect 107672 138366 107746 138394
rect 108500 138366 108574 138394
rect 109420 138366 109494 138394
rect 110248 138366 110322 138394
rect 111076 138366 111150 138394
rect 111996 138366 112070 138394
rect 112824 138366 112898 138394
rect 113744 138366 113818 138394
rect 114572 138366 114646 138394
rect 115400 138366 115474 138394
rect 116320 138366 116394 138394
rect 117148 138366 117222 138394
rect 117976 138366 118050 138394
rect 118896 138366 118970 138394
rect 119724 138366 119798 138394
rect 120552 138366 120626 138394
rect 121518 138394 121546 138652
rect 122346 138394 122374 138652
rect 123266 138394 123294 138652
rect 124094 138394 124122 138652
rect 124922 138394 124950 138652
rect 125842 138394 125870 138652
rect 126670 138394 126698 138652
rect 127498 138394 127526 138652
rect 128418 138394 128446 138652
rect 129246 138394 129274 138652
rect 130074 138394 130102 138652
rect 130994 138394 131022 138652
rect 131822 138394 131850 138652
rect 132742 138394 132770 138652
rect 133570 138394 133598 138652
rect 134398 138394 134426 138652
rect 135318 138394 135346 138652
rect 136146 138394 136174 138652
rect 136974 138394 137002 138652
rect 137894 138394 137922 138652
rect 138722 138394 138750 138652
rect 139550 138394 139578 138652
rect 140470 138394 140498 138652
rect 141298 138394 141326 138652
rect 142126 138394 142154 138652
rect 143046 138394 143074 138652
rect 143874 138394 143902 138652
rect 144794 138394 144822 138652
rect 145622 138394 145650 138652
rect 146450 138394 146478 138652
rect 147370 138394 147398 138652
rect 148198 138394 148226 138652
rect 149026 138394 149054 138652
rect 149946 138394 149974 138652
rect 150774 138394 150802 138652
rect 151602 138394 151630 138652
rect 152522 138394 152550 138652
rect 153350 138394 153378 138652
rect 154270 138394 154298 138652
rect 155098 138394 155126 138652
rect 155926 138394 155954 138652
rect 156846 138394 156874 138652
rect 157674 138394 157702 138652
rect 158502 138394 158530 138652
rect 159422 138394 159450 138652
rect 160250 138394 160278 138652
rect 161078 138394 161106 138652
rect 121518 138366 121684 138394
rect 94044 4208 94096 4214
rect 94044 4150 94096 4156
rect 94792 3777 94820 138366
rect 95056 135992 95108 135998
rect 95056 135934 95108 135940
rect 95068 16574 95096 135934
rect 95620 135454 95648 138366
rect 95608 135448 95660 135454
rect 95608 135390 95660 135396
rect 96448 135182 96476 138366
rect 96436 135176 96488 135182
rect 96436 135118 96488 135124
rect 95068 16546 95188 16574
rect 94778 3768 94834 3777
rect 94778 3703 94834 3712
rect 95160 480 95188 16546
rect 97368 3670 97396 138366
rect 97908 24132 97960 24138
rect 97908 24074 97960 24080
rect 97920 3670 97948 24074
rect 97356 3664 97408 3670
rect 97356 3606 97408 3612
rect 97448 3664 97500 3670
rect 97448 3606 97500 3612
rect 97908 3664 97960 3670
rect 97908 3606 97960 3612
rect 96252 3528 96304 3534
rect 96252 3470 96304 3476
rect 96264 480 96292 3470
rect 97460 480 97488 3606
rect 98196 3602 98224 138366
rect 99024 136134 99052 138366
rect 99012 136128 99064 136134
rect 99012 136070 99064 136076
rect 99944 134774 99972 138366
rect 99932 134768 99984 134774
rect 99932 134710 99984 134716
rect 100772 3942 100800 138366
rect 101692 135658 101720 138366
rect 101680 135652 101732 135658
rect 101680 135594 101732 135600
rect 102520 134842 102548 138366
rect 102508 134836 102560 134842
rect 102508 134778 102560 134784
rect 103348 6914 103376 138366
rect 104164 136196 104216 136202
rect 104164 136138 104216 136144
rect 104176 134910 104204 136138
rect 104164 134904 104216 134910
rect 104164 134846 104216 134852
rect 104268 26926 104296 138366
rect 105096 133210 105124 138366
rect 105084 133204 105136 133210
rect 105084 133146 105136 133152
rect 104256 26920 104308 26926
rect 104256 26862 104308 26868
rect 104808 25560 104860 25566
rect 104808 25502 104860 25508
rect 104820 6914 104848 25502
rect 105924 6914 105952 138366
rect 106844 134706 106872 138366
rect 107568 136128 107620 136134
rect 107568 136070 107620 136076
rect 106832 134700 106884 134706
rect 106832 134642 106884 134648
rect 103256 6886 103376 6914
rect 104544 6886 104848 6914
rect 105648 6886 105952 6914
rect 101036 4616 101088 4622
rect 101036 4558 101088 4564
rect 100760 3936 100812 3942
rect 100760 3878 100812 3884
rect 98644 3664 98696 3670
rect 98644 3606 98696 3612
rect 98184 3596 98236 3602
rect 98184 3538 98236 3544
rect 98656 480 98684 3606
rect 99840 3596 99892 3602
rect 99840 3538 99892 3544
rect 99852 480 99880 3538
rect 101048 480 101076 4558
rect 102232 3936 102284 3942
rect 102232 3878 102284 3884
rect 102244 480 102272 3878
rect 103256 3738 103284 6886
rect 103244 3732 103296 3738
rect 103244 3674 103296 3680
rect 103336 3732 103388 3738
rect 103336 3674 103388 3680
rect 103348 480 103376 3674
rect 104544 480 104572 6886
rect 105648 3806 105676 6886
rect 105636 3800 105688 3806
rect 105636 3742 105688 3748
rect 105728 3800 105780 3806
rect 105728 3742 105780 3748
rect 105740 480 105768 3742
rect 107580 3398 107608 136070
rect 107672 32434 107700 138366
rect 107660 32428 107712 32434
rect 107660 32370 107712 32376
rect 108120 6248 108172 6254
rect 108120 6190 108172 6196
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 107568 3392 107620 3398
rect 107568 3334 107620 3340
rect 106936 480 106964 3334
rect 108132 480 108160 6190
rect 108500 3874 108528 138366
rect 109420 136202 109448 138366
rect 109408 136196 109460 136202
rect 109408 136138 109460 136144
rect 110248 4146 110276 138366
rect 110236 4140 110288 4146
rect 110236 4082 110288 4088
rect 109316 4072 109368 4078
rect 109316 4014 109368 4020
rect 108488 3868 108540 3874
rect 108488 3810 108540 3816
rect 109328 480 109356 4014
rect 111076 4010 111104 138366
rect 111996 136610 112024 138366
rect 111984 136604 112036 136610
rect 111984 136546 112036 136552
rect 111616 7608 111668 7614
rect 111616 7550 111668 7556
rect 111064 4004 111116 4010
rect 111064 3946 111116 3952
rect 110512 3868 110564 3874
rect 110512 3810 110564 3816
rect 110524 480 110552 3810
rect 111628 480 111656 7550
rect 112824 4146 112852 138366
rect 113088 136196 113140 136202
rect 113088 136138 113140 136144
rect 113100 6914 113128 136138
rect 112916 6886 113128 6914
rect 112812 4140 112864 4146
rect 112812 4082 112864 4088
rect 112916 3482 112944 6886
rect 112824 3454 112944 3482
rect 112824 480 112852 3454
rect 113744 3398 113772 138366
rect 114572 5098 114600 138366
rect 115296 136604 115348 136610
rect 115296 136546 115348 136552
rect 115308 135046 115336 136546
rect 115400 136270 115428 138366
rect 115388 136264 115440 136270
rect 115388 136206 115440 136212
rect 115296 135040 115348 135046
rect 115296 134982 115348 134988
rect 115204 7676 115256 7682
rect 115204 7618 115256 7624
rect 114560 5092 114612 5098
rect 114560 5034 114612 5040
rect 114008 4004 114060 4010
rect 114008 3946 114060 3952
rect 113732 3392 113784 3398
rect 113732 3334 113784 3340
rect 114020 480 114048 3946
rect 115216 480 115244 7618
rect 116320 3330 116348 138366
rect 117148 5166 117176 138366
rect 117976 136610 118004 138366
rect 117964 136604 118016 136610
rect 117964 136546 118016 136552
rect 117228 136264 117280 136270
rect 117228 136206 117280 136212
rect 117136 5160 117188 5166
rect 117136 5102 117188 5108
rect 117240 3398 117268 136206
rect 118792 6316 118844 6322
rect 118792 6258 118844 6264
rect 116400 3392 116452 3398
rect 116400 3334 116452 3340
rect 117228 3392 117280 3398
rect 117228 3334 117280 3340
rect 116308 3324 116360 3330
rect 116308 3266 116360 3272
rect 116412 480 116440 3334
rect 117596 3324 117648 3330
rect 117596 3266 117648 3272
rect 117608 480 117636 3266
rect 118804 480 118832 6258
rect 118896 3262 118924 138366
rect 119724 5234 119752 138366
rect 120552 135794 120580 138366
rect 120540 135788 120592 135794
rect 120540 135730 120592 135736
rect 119712 5228 119764 5234
rect 119712 5170 119764 5176
rect 121092 3392 121144 3398
rect 121092 3334 121144 3340
rect 118884 3256 118936 3262
rect 118884 3198 118936 3204
rect 119896 3256 119948 3262
rect 119896 3198 119948 3204
rect 119908 480 119936 3198
rect 121104 480 121132 3334
rect 121656 3194 121684 138366
rect 122300 138366 122374 138394
rect 123220 138366 123294 138394
rect 124048 138366 124122 138394
rect 124876 138366 124950 138394
rect 125796 138366 125870 138394
rect 126624 138366 126698 138394
rect 127452 138366 127526 138394
rect 128372 138366 128446 138394
rect 129200 138366 129274 138394
rect 130028 138366 130102 138394
rect 130948 138366 131022 138394
rect 131776 138366 131850 138394
rect 132696 138366 132770 138394
rect 133524 138366 133598 138394
rect 134352 138366 134426 138394
rect 135272 138366 135346 138394
rect 136100 138366 136174 138394
rect 136928 138366 137002 138394
rect 137848 138366 137922 138394
rect 138676 138366 138750 138394
rect 139504 138366 139578 138394
rect 140424 138366 140498 138394
rect 141252 138366 141326 138394
rect 142080 138366 142154 138394
rect 143000 138366 143074 138394
rect 143828 138366 143902 138394
rect 144748 138366 144822 138394
rect 145576 138366 145650 138394
rect 146404 138366 146478 138394
rect 147324 138366 147398 138394
rect 148152 138366 148226 138394
rect 148980 138366 149054 138394
rect 149900 138366 149974 138394
rect 150728 138366 150802 138394
rect 151556 138366 151630 138394
rect 152476 138366 152550 138394
rect 153304 138366 153378 138394
rect 154224 138366 154298 138394
rect 155052 138366 155126 138394
rect 155880 138366 155954 138394
rect 156800 138366 156874 138394
rect 157628 138366 157702 138394
rect 158456 138366 158530 138394
rect 159376 138366 159450 138394
rect 160112 138366 160278 138394
rect 161032 138366 161106 138394
rect 161572 138440 161624 138446
rect 161998 138394 162026 138652
rect 162826 138446 162854 138652
rect 161572 138382 161624 138388
rect 122300 5302 122328 138366
rect 123220 135590 123248 138366
rect 123208 135584 123260 135590
rect 123208 135526 123260 135532
rect 122380 6384 122432 6390
rect 122380 6326 122432 6332
rect 122288 5296 122340 5302
rect 122288 5238 122340 5244
rect 122392 3210 122420 6326
rect 121644 3188 121696 3194
rect 121644 3130 121696 3136
rect 122300 3182 122420 3210
rect 123484 3256 123536 3262
rect 123484 3198 123536 3204
rect 122300 480 122328 3182
rect 123496 480 123524 3198
rect 124048 3058 124076 138366
rect 124128 136604 124180 136610
rect 124128 136546 124180 136552
rect 124140 3262 124168 136546
rect 124876 134978 124904 138366
rect 125796 136542 125824 138366
rect 125784 136536 125836 136542
rect 125784 136478 125836 136484
rect 126244 136536 126296 136542
rect 126244 136478 126296 136484
rect 125508 135788 125560 135794
rect 125508 135730 125560 135736
rect 124864 134972 124916 134978
rect 124864 134914 124916 134920
rect 125520 3262 125548 135730
rect 125876 5092 125928 5098
rect 125876 5034 125928 5040
rect 124128 3256 124180 3262
rect 124128 3198 124180 3204
rect 124680 3256 124732 3262
rect 124680 3198 124732 3204
rect 125508 3256 125560 3262
rect 125508 3198 125560 3204
rect 124036 3052 124088 3058
rect 124036 2994 124088 3000
rect 124692 480 124720 3198
rect 125888 480 125916 5034
rect 126256 4690 126284 136478
rect 126244 4684 126296 4690
rect 126244 4626 126296 4632
rect 126624 3126 126652 138366
rect 127452 5438 127480 138366
rect 127440 5432 127492 5438
rect 127440 5374 127492 5380
rect 128372 5370 128400 138366
rect 128360 5364 128412 5370
rect 128360 5306 128412 5312
rect 128176 5024 128228 5030
rect 128176 4966 128228 4972
rect 126980 4684 127032 4690
rect 126980 4626 127032 4632
rect 126612 3120 126664 3126
rect 126612 3062 126664 3068
rect 126992 480 127020 4626
rect 128188 480 128216 4966
rect 129200 2990 129228 138366
rect 130028 135522 130056 138366
rect 130384 135652 130436 135658
rect 130384 135594 130436 135600
rect 130016 135516 130068 135522
rect 130016 135458 130068 135464
rect 129372 5364 129424 5370
rect 129372 5306 129424 5312
rect 129188 2984 129240 2990
rect 129188 2926 129240 2932
rect 129384 480 129412 5306
rect 130396 4622 130424 135594
rect 130948 71058 130976 138366
rect 131776 136338 131804 138366
rect 131764 136332 131816 136338
rect 131764 136274 131816 136280
rect 130936 71052 130988 71058
rect 130936 70994 130988 71000
rect 132696 5506 132724 138366
rect 133524 136474 133552 138366
rect 133512 136468 133564 136474
rect 133512 136410 133564 136416
rect 133144 135516 133196 135522
rect 133144 135458 133196 135464
rect 132960 7744 133012 7750
rect 132960 7686 133012 7692
rect 132684 5500 132736 5506
rect 132684 5442 132736 5448
rect 131764 5228 131816 5234
rect 131764 5170 131816 5176
rect 130568 5160 130620 5166
rect 130568 5102 130620 5108
rect 130384 4616 130436 4622
rect 130384 4558 130436 4564
rect 130580 480 130608 5102
rect 131776 480 131804 5170
rect 132972 480 133000 7686
rect 133156 7682 133184 135458
rect 133144 7676 133196 7682
rect 133144 7618 133196 7624
rect 134156 3460 134208 3466
rect 134156 3402 134208 3408
rect 134168 480 134196 3402
rect 134352 2922 134380 138366
rect 135272 135266 135300 138366
rect 136100 136542 136128 138366
rect 136088 136536 136140 136542
rect 136088 136478 136140 136484
rect 136928 136406 136956 138366
rect 136916 136400 136968 136406
rect 136916 136342 136968 136348
rect 137284 135584 137336 135590
rect 137284 135526 137336 135532
rect 135180 135238 135300 135266
rect 135180 135114 135208 135238
rect 135168 135108 135220 135114
rect 135168 135050 135220 135056
rect 135168 134632 135220 134638
rect 135168 134574 135220 134580
rect 135180 3466 135208 134574
rect 137296 8974 137324 135526
rect 137284 8968 137336 8974
rect 137284 8910 137336 8916
rect 137652 8968 137704 8974
rect 137652 8910 137704 8916
rect 135260 5432 135312 5438
rect 135260 5374 135312 5380
rect 135168 3460 135220 3466
rect 135168 3402 135220 3408
rect 134340 2916 134392 2922
rect 134340 2858 134392 2864
rect 135272 480 135300 5374
rect 136456 5296 136508 5302
rect 136456 5238 136508 5244
rect 136468 480 136496 5238
rect 137664 480 137692 8910
rect 137848 4758 137876 138366
rect 138676 135862 138704 138366
rect 138664 135856 138716 135862
rect 138664 135798 138716 135804
rect 138848 6452 138900 6458
rect 138848 6394 138900 6400
rect 137836 4752 137888 4758
rect 137836 4694 137888 4700
rect 138860 480 138888 6394
rect 139504 2854 139532 138366
rect 140424 135590 140452 138366
rect 140780 136400 140832 136406
rect 140780 136342 140832 136348
rect 140412 135584 140464 135590
rect 140412 135526 140464 135532
rect 140792 134570 140820 136342
rect 140780 134564 140832 134570
rect 140780 134506 140832 134512
rect 141252 4826 141280 138366
rect 142080 135726 142108 138366
rect 142804 136536 142856 136542
rect 142804 136478 142856 136484
rect 142068 135720 142120 135726
rect 142068 135662 142120 135668
rect 142068 134564 142120 134570
rect 142068 134506 142120 134512
rect 141240 4820 141292 4826
rect 141240 4762 141292 4768
rect 140044 4548 140096 4554
rect 140044 4490 140096 4496
rect 139492 2848 139544 2854
rect 139492 2790 139544 2796
rect 140056 480 140084 4490
rect 142080 3466 142108 134506
rect 142436 6112 142488 6118
rect 142436 6054 142488 6060
rect 141240 3460 141292 3466
rect 141240 3402 141292 3408
rect 142068 3460 142120 3466
rect 142068 3402 142120 3408
rect 141252 480 141280 3402
rect 142448 480 142476 6054
rect 142816 4690 142844 136478
rect 143000 6186 143028 138366
rect 143828 135930 143856 138366
rect 144184 136332 144236 136338
rect 144184 136274 144236 136280
rect 143816 135924 143868 135930
rect 143816 135866 143868 135872
rect 142988 6180 143040 6186
rect 142988 6122 143040 6128
rect 143540 4820 143592 4826
rect 143540 4762 143592 4768
rect 142804 4684 142856 4690
rect 142804 4626 142856 4632
rect 143552 480 143580 4762
rect 144196 4554 144224 136274
rect 144748 6914 144776 138366
rect 145576 136406 145604 138366
rect 145564 136400 145616 136406
rect 145564 136342 145616 136348
rect 144656 6886 144776 6914
rect 144184 4548 144236 4554
rect 144184 4490 144236 4496
rect 144656 3262 144684 6886
rect 144736 6520 144788 6526
rect 144736 6462 144788 6468
rect 144644 3256 144696 3262
rect 144644 3198 144696 3204
rect 144748 480 144776 6462
rect 146404 4894 146432 138366
rect 147324 136066 147352 138366
rect 147312 136060 147364 136066
rect 147312 136002 147364 136008
rect 146944 135856 146996 135862
rect 146944 135798 146996 135804
rect 146956 7750 146984 135798
rect 146944 7744 146996 7750
rect 146944 7686 146996 7692
rect 147128 7676 147180 7682
rect 147128 7618 147180 7624
rect 146392 4888 146444 4894
rect 146392 4830 146444 4836
rect 145932 3460 145984 3466
rect 145932 3402 145984 3408
rect 145944 480 145972 3402
rect 147140 480 147168 7618
rect 148152 4962 148180 138366
rect 148980 136066 149008 138366
rect 148968 136060 149020 136066
rect 148968 136002 149020 136008
rect 148968 135924 149020 135930
rect 148968 135866 149020 135872
rect 148140 4956 148192 4962
rect 148140 4898 148192 4904
rect 148980 3534 149008 135866
rect 149900 3942 149928 138366
rect 150728 24138 150756 138366
rect 150716 24132 150768 24138
rect 150716 24074 150768 24080
rect 150624 4888 150676 4894
rect 150624 4830 150676 4836
rect 149888 3936 149940 3942
rect 149888 3878 149940 3884
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 148336 480 148364 3470
rect 149520 3188 149572 3194
rect 149520 3130 149572 3136
rect 149532 480 149560 3130
rect 150636 480 150664 4830
rect 151556 3670 151584 138366
rect 151544 3664 151596 3670
rect 151544 3606 151596 3612
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 151832 480 151860 3470
rect 152476 3262 152504 138366
rect 153108 136060 153160 136066
rect 153108 136002 153160 136008
rect 153016 135992 153068 135998
rect 153016 135934 153068 135940
rect 152464 3256 152516 3262
rect 152464 3198 152516 3204
rect 153028 480 153056 135934
rect 153120 3534 153148 136002
rect 153304 135658 153332 138366
rect 153292 135652 153344 135658
rect 153292 135594 153344 135600
rect 154224 6914 154252 138366
rect 154132 6886 154252 6914
rect 154132 3602 154160 6886
rect 154212 4752 154264 4758
rect 154212 4694 154264 4700
rect 154120 3596 154172 3602
rect 154120 3538 154172 3544
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 154224 480 154252 4694
rect 155052 3738 155080 138366
rect 155880 25566 155908 138366
rect 155868 25560 155920 25566
rect 155868 25502 155920 25508
rect 156800 3806 156828 138366
rect 157628 136134 157656 138366
rect 157616 136128 157668 136134
rect 157616 136070 157668 136076
rect 158456 6254 158484 138366
rect 158444 6248 158496 6254
rect 158444 6190 158496 6196
rect 157800 4956 157852 4962
rect 157800 4898 157852 4904
rect 156788 3800 156840 3806
rect 156788 3742 156840 3748
rect 155040 3732 155092 3738
rect 155040 3674 155092 3680
rect 156604 3664 156656 3670
rect 156604 3606 156656 3612
rect 155408 3596 155460 3602
rect 155408 3538 155460 3544
rect 155420 480 155448 3538
rect 156616 480 156644 3606
rect 157812 480 157840 4898
rect 159376 4146 159404 138366
rect 160008 136128 160060 136134
rect 160008 136070 160060 136076
rect 159364 4140 159416 4146
rect 159364 4082 159416 4088
rect 160020 3534 160048 136070
rect 160112 3942 160140 138366
rect 161032 7614 161060 138366
rect 161020 7608 161072 7614
rect 161020 7550 161072 7556
rect 161296 5500 161348 5506
rect 161296 5442 161348 5448
rect 160100 3936 160152 3942
rect 160100 3878 160152 3884
rect 160100 3800 160152 3806
rect 160100 3742 160152 3748
rect 158904 3528 158956 3534
rect 158904 3470 158956 3476
rect 160008 3528 160060 3534
rect 160008 3470 160060 3476
rect 158916 480 158944 3470
rect 160112 480 160140 3742
rect 161308 480 161336 5442
rect 161584 4010 161612 138382
rect 161952 138366 162026 138394
rect 162814 138440 162866 138446
rect 163746 138394 163774 138652
rect 164574 138394 164602 138652
rect 165402 138394 165430 138652
rect 166322 138394 166350 138652
rect 167150 138394 167178 138652
rect 167978 138394 168006 138652
rect 168898 138394 168926 138652
rect 169726 138394 169754 138652
rect 162814 138382 162866 138388
rect 163700 138366 163774 138394
rect 164528 138366 164602 138394
rect 165356 138366 165430 138394
rect 166276 138366 166350 138394
rect 167012 138366 167178 138394
rect 167932 138366 168006 138394
rect 168852 138366 168926 138394
rect 169680 138366 169754 138394
rect 170554 138394 170582 138652
rect 171474 138394 171502 138652
rect 172302 138394 172330 138652
rect 173130 138394 173158 138652
rect 174050 138394 174078 138652
rect 174878 138394 174906 138652
rect 175798 138394 175826 138652
rect 176626 138394 176654 138652
rect 177454 138394 177482 138652
rect 178374 138394 178402 138652
rect 179202 138394 179230 138652
rect 180030 138394 180058 138652
rect 180950 138394 180978 138652
rect 181778 138394 181806 138652
rect 182606 138394 182634 138652
rect 183526 138394 183554 138652
rect 184354 138394 184382 138652
rect 185274 138394 185302 138652
rect 186102 138394 186130 138652
rect 186930 138394 186958 138652
rect 187850 138394 187878 138652
rect 188678 138394 188706 138652
rect 189506 138394 189534 138652
rect 190426 138394 190454 138652
rect 191254 138394 191282 138652
rect 192082 138394 192110 138652
rect 193002 138394 193030 138652
rect 193830 138394 193858 138652
rect 194750 138394 194778 138652
rect 195578 138394 195606 138652
rect 196406 138394 196434 138652
rect 197326 138394 197354 138652
rect 198154 138394 198182 138652
rect 198982 138394 199010 138652
rect 199902 138394 199930 138652
rect 200730 138394 200758 138652
rect 201558 138394 201586 138652
rect 202478 138394 202506 138652
rect 203306 138394 203334 138652
rect 204134 138394 204162 138652
rect 205054 138394 205082 138652
rect 205882 138394 205910 138652
rect 206802 138394 206830 138652
rect 207630 138394 207658 138652
rect 208458 138394 208486 138652
rect 209378 138394 209406 138652
rect 210206 138394 210234 138652
rect 211034 138394 211062 138652
rect 211954 138394 211982 138652
rect 212782 138394 212810 138652
rect 213610 138394 213638 138652
rect 214530 138394 214558 138652
rect 170554 138366 170628 138394
rect 161952 136202 161980 138366
rect 161940 136196 161992 136202
rect 161940 136138 161992 136144
rect 162768 136196 162820 136202
rect 162768 136138 162820 136144
rect 162780 6914 162808 136138
rect 163700 135590 163728 138366
rect 164528 136270 164556 138366
rect 164516 136264 164568 136270
rect 164516 136206 164568 136212
rect 163688 135584 163740 135590
rect 163688 135526 163740 135532
rect 162504 6886 162808 6914
rect 161572 4004 161624 4010
rect 161572 3946 161624 3952
rect 162504 480 162532 6886
rect 164884 4684 164936 4690
rect 164884 4626 164936 4632
rect 163688 3732 163740 3738
rect 163688 3674 163740 3680
rect 163700 480 163728 3674
rect 164896 480 164924 4626
rect 165356 3330 165384 138366
rect 166276 6322 166304 138366
rect 166908 136264 166960 136270
rect 166908 136206 166960 136212
rect 166264 6316 166316 6322
rect 166264 6258 166316 6264
rect 166920 3534 166948 136206
rect 167012 4078 167040 138366
rect 167000 4072 167052 4078
rect 167000 4014 167052 4020
rect 167184 3868 167236 3874
rect 167184 3810 167236 3816
rect 166080 3528 166132 3534
rect 166080 3470 166132 3476
rect 166908 3528 166960 3534
rect 166908 3470 166960 3476
rect 165344 3324 165396 3330
rect 165344 3266 165396 3272
rect 166092 480 166120 3470
rect 167196 480 167224 3810
rect 167932 3398 167960 138366
rect 168852 6390 168880 138366
rect 169680 136610 169708 138366
rect 169668 136604 169720 136610
rect 169668 136546 169720 136552
rect 170496 136604 170548 136610
rect 170496 136546 170548 136552
rect 170404 136468 170456 136474
rect 170404 136410 170456 136416
rect 169576 136400 169628 136406
rect 169576 136342 169628 136348
rect 168840 6384 168892 6390
rect 168840 6326 168892 6332
rect 168380 4616 168432 4622
rect 168380 4558 168432 4564
rect 167920 3392 167972 3398
rect 167920 3334 167972 3340
rect 168392 480 168420 4558
rect 169588 480 169616 136342
rect 170416 5370 170444 136410
rect 170404 5364 170456 5370
rect 170404 5306 170456 5312
rect 170508 5098 170536 136546
rect 170600 135794 170628 138366
rect 171428 138366 171502 138394
rect 172256 138366 172330 138394
rect 173084 138366 173158 138394
rect 174004 138366 174078 138394
rect 174832 138366 174906 138394
rect 175752 138366 175826 138394
rect 176580 138366 176654 138394
rect 177408 138366 177482 138394
rect 178328 138366 178402 138394
rect 179156 138366 179230 138394
rect 179984 138366 180058 138394
rect 180904 138366 180978 138394
rect 181732 138366 181806 138394
rect 182560 138366 182634 138394
rect 183480 138366 183554 138394
rect 184308 138366 184382 138394
rect 185228 138366 185302 138394
rect 186056 138366 186130 138394
rect 186884 138366 186958 138394
rect 187804 138366 187878 138394
rect 188632 138366 188706 138394
rect 189460 138366 189534 138394
rect 190288 138366 190454 138394
rect 191208 138366 191282 138394
rect 192036 138366 192110 138394
rect 192956 138366 193030 138394
rect 193784 138366 193858 138394
rect 194704 138366 194778 138394
rect 195532 138366 195606 138394
rect 196360 138366 196434 138394
rect 197280 138366 197354 138394
rect 198108 138366 198182 138394
rect 198936 138366 199010 138394
rect 199856 138366 199930 138394
rect 200684 138366 200758 138394
rect 201512 138366 201586 138394
rect 202432 138366 202506 138394
rect 203260 138366 203334 138394
rect 204088 138366 204162 138394
rect 205008 138366 205082 138394
rect 205836 138366 205910 138394
rect 206756 138366 206830 138394
rect 207584 138366 207658 138394
rect 208412 138366 208486 138394
rect 209332 138366 209406 138394
rect 210160 138366 210234 138394
rect 210988 138366 211062 138394
rect 211908 138366 211982 138394
rect 212736 138366 212810 138394
rect 213564 138366 213638 138394
rect 214484 138366 214558 138394
rect 215358 138394 215386 138652
rect 216278 138394 216306 138652
rect 217106 138394 217134 138652
rect 217934 138394 217962 138652
rect 218854 138394 218882 138652
rect 219682 138394 219710 138652
rect 220510 138394 220538 138652
rect 221430 138394 221458 138652
rect 222258 138394 222286 138652
rect 223086 138394 223114 138652
rect 224006 138394 224034 138652
rect 224834 138394 224862 138652
rect 225754 138394 225782 138652
rect 226582 138394 226610 138652
rect 227410 138394 227438 138652
rect 228330 138394 228358 138652
rect 229158 138394 229186 138652
rect 229986 138394 230014 138652
rect 230906 138394 230934 138652
rect 231734 138394 231762 138652
rect 232562 138394 232590 138652
rect 233482 138394 233510 138652
rect 234310 138394 234338 138652
rect 235138 138394 235166 138652
rect 236058 138394 236086 138652
rect 236886 138394 236914 138652
rect 237806 138394 237834 138652
rect 238634 138394 238662 138652
rect 239462 138394 239490 138652
rect 240382 138394 240410 138652
rect 241210 138394 241238 138652
rect 242038 138394 242066 138652
rect 242958 138394 242986 138652
rect 243786 138394 243814 138652
rect 244614 138394 244642 138652
rect 245534 138394 245562 138652
rect 246362 138394 246390 138652
rect 247282 138394 247310 138652
rect 248110 138394 248138 138652
rect 248938 138394 248966 138652
rect 249858 138394 249886 138652
rect 250686 138394 250714 138652
rect 251514 138394 251542 138652
rect 252434 138394 252462 138652
rect 253262 138394 253290 138652
rect 254090 138394 254118 138652
rect 255010 138394 255038 138652
rect 255838 138394 255866 138652
rect 256758 138394 256786 138652
rect 257586 138394 257614 138652
rect 258414 138394 258442 138652
rect 259334 138394 259362 138652
rect 260162 138394 260190 138652
rect 260990 138394 261018 138652
rect 261910 138394 261938 138652
rect 262738 138394 262766 138652
rect 263566 138394 263594 138652
rect 264486 138394 264514 138652
rect 265314 138394 265342 138652
rect 266142 138394 266170 138652
rect 267062 138394 267090 138652
rect 267890 138394 267918 138652
rect 268810 138394 268838 138652
rect 269638 138394 269666 138652
rect 270466 138394 270494 138652
rect 271386 138394 271414 138652
rect 272214 138394 272242 138652
rect 273042 138394 273070 138652
rect 273962 138394 273990 138652
rect 274790 138394 274818 138652
rect 275618 138394 275646 138652
rect 276538 138394 276566 138652
rect 277366 138394 277394 138652
rect 278286 138394 278314 138652
rect 279114 138394 279142 138652
rect 279942 138394 279970 138652
rect 280862 138394 280890 138652
rect 281690 138394 281718 138652
rect 282518 138394 282546 138652
rect 283438 138394 283466 138652
rect 284266 138394 284294 138652
rect 285094 138394 285122 138652
rect 286014 138394 286042 138652
rect 286842 138394 286870 138652
rect 287762 138394 287790 138652
rect 288590 138394 288618 138652
rect 289418 138394 289446 138652
rect 290338 138394 290366 138652
rect 291166 138394 291194 138652
rect 291994 138394 292022 138652
rect 292914 138394 292942 138652
rect 293742 138394 293770 138652
rect 294570 138394 294598 138652
rect 295490 138394 295518 138652
rect 215358 138366 215432 138394
rect 171428 136610 171456 138366
rect 171416 136604 171468 136610
rect 171416 136546 171468 136552
rect 172256 136542 172284 138366
rect 172244 136536 172296 136542
rect 172244 136478 172296 136484
rect 170588 135788 170640 135794
rect 170588 135730 170640 135736
rect 170496 5092 170548 5098
rect 170496 5034 170548 5040
rect 171968 5092 172020 5098
rect 171968 5034 172020 5040
rect 170772 3936 170824 3942
rect 170772 3878 170824 3884
rect 170784 480 170812 3878
rect 171980 480 172008 5034
rect 173084 5030 173112 138366
rect 173808 136536 173860 136542
rect 173808 136478 173860 136484
rect 173072 5024 173124 5030
rect 173072 4966 173124 4972
rect 173820 3534 173848 136478
rect 174004 136474 174032 138366
rect 173992 136468 174044 136474
rect 173992 136410 174044 136416
rect 174832 5166 174860 138366
rect 175752 5234 175780 138366
rect 176580 135862 176608 138366
rect 176568 135856 176620 135862
rect 176568 135798 176620 135804
rect 177408 134638 177436 138366
rect 177856 136536 177908 136542
rect 177856 136478 177908 136484
rect 177396 134632 177448 134638
rect 177396 134574 177448 134580
rect 175740 5228 175792 5234
rect 175740 5170 175792 5176
rect 174820 5160 174872 5166
rect 174820 5102 174872 5108
rect 175464 4140 175516 4146
rect 175464 4082 175516 4088
rect 174268 4004 174320 4010
rect 174268 3946 174320 3952
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 173176 480 173204 3470
rect 174280 480 174308 3946
rect 175476 480 175504 4082
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 176672 480 176700 3470
rect 177868 480 177896 136478
rect 177948 135856 178000 135862
rect 177948 135798 178000 135804
rect 177960 3534 177988 135798
rect 178328 5438 178356 138366
rect 178316 5432 178368 5438
rect 178316 5374 178368 5380
rect 179156 5302 179184 138366
rect 179984 8974 180012 138366
rect 180708 136604 180760 136610
rect 180708 136546 180760 136552
rect 180064 135720 180116 135726
rect 180064 135662 180116 135668
rect 179972 8968 180024 8974
rect 179972 8910 180024 8916
rect 180076 6526 180104 135662
rect 180064 6520 180116 6526
rect 180064 6462 180116 6468
rect 179144 5296 179196 5302
rect 179144 5238 179196 5244
rect 179052 4072 179104 4078
rect 179052 4014 179104 4020
rect 177948 3528 178000 3534
rect 177948 3470 178000 3476
rect 179064 480 179092 4014
rect 180720 3534 180748 136546
rect 180904 6458 180932 138366
rect 181732 136338 181760 138366
rect 181720 136332 181772 136338
rect 181720 136274 181772 136280
rect 182560 134570 182588 138366
rect 182548 134564 182600 134570
rect 182548 134506 182600 134512
rect 180892 6452 180944 6458
rect 180892 6394 180944 6400
rect 183480 6186 183508 138366
rect 183468 6180 183520 6186
rect 183468 6122 183520 6128
rect 184308 4826 184336 138366
rect 185228 135726 185256 138366
rect 185216 135720 185268 135726
rect 185216 135662 185268 135668
rect 184848 135516 184900 135522
rect 184848 135458 184900 135464
rect 184296 4820 184348 4826
rect 184296 4762 184348 4768
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 180260 480 180288 3470
rect 184860 3466 184888 135458
rect 183744 3460 183796 3466
rect 183744 3402 183796 3408
rect 184848 3460 184900 3466
rect 184848 3402 184900 3408
rect 181444 3392 181496 3398
rect 181444 3334 181496 3340
rect 181456 480 181484 3334
rect 182548 3324 182600 3330
rect 182548 3266 182600 3272
rect 182560 480 182588 3266
rect 183756 480 183784 3402
rect 184940 3256 184992 3262
rect 184940 3198 184992 3204
rect 184952 480 184980 3198
rect 186056 3194 186084 138366
rect 186884 7682 186912 138366
rect 186964 136332 187016 136338
rect 186964 136274 187016 136280
rect 186872 7676 186924 7682
rect 186872 7618 186924 7624
rect 186976 4758 187004 136274
rect 187608 136060 187660 136066
rect 187608 136002 187660 136008
rect 187620 6914 187648 136002
rect 187804 135930 187832 138366
rect 187792 135924 187844 135930
rect 187792 135866 187844 135872
rect 188344 135584 188396 135590
rect 188344 135526 188396 135532
rect 187344 6886 187648 6914
rect 186964 4752 187016 4758
rect 186964 4694 187016 4700
rect 186044 3188 186096 3194
rect 186044 3130 186096 3136
rect 186136 2848 186188 2854
rect 186136 2790 186188 2796
rect 186148 480 186176 2790
rect 187344 480 187372 6886
rect 188356 4894 188384 135526
rect 188344 4888 188396 4894
rect 188344 4830 188396 4836
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 188540 480 188568 3470
rect 188632 3126 188660 138366
rect 189460 135590 189488 138366
rect 190288 135794 190316 138366
rect 191208 135794 191236 138366
rect 192036 136338 192064 138366
rect 192024 136332 192076 136338
rect 192024 136274 192076 136280
rect 191748 135924 191800 135930
rect 191748 135866 191800 135872
rect 190276 135788 190328 135794
rect 190276 135730 190328 135736
rect 191196 135788 191248 135794
rect 191196 135730 191248 135736
rect 189448 135584 189500 135590
rect 189448 135526 189500 135532
rect 191104 135516 191156 135522
rect 191104 135458 191156 135464
rect 191116 5098 191144 135458
rect 191104 5092 191156 5098
rect 191104 5034 191156 5040
rect 189724 3188 189776 3194
rect 189724 3130 189776 3136
rect 188620 3120 188672 3126
rect 188620 3062 188672 3068
rect 189736 480 189764 3130
rect 191760 3058 191788 135866
rect 192956 3466 192984 138366
rect 193784 3670 193812 138366
rect 194704 4962 194732 138366
rect 195532 136134 195560 138366
rect 195520 136128 195572 136134
rect 195520 136070 195572 136076
rect 195336 135992 195388 135998
rect 195336 135934 195388 135940
rect 195348 122834 195376 135934
rect 195256 122806 195376 122834
rect 194692 4956 194744 4962
rect 194692 4898 194744 4904
rect 193772 3664 193824 3670
rect 193772 3606 193824 3612
rect 195256 3466 195284 122806
rect 196360 3806 196388 138366
rect 197280 5506 197308 138366
rect 198108 136202 198136 138366
rect 198096 136196 198148 136202
rect 198096 136138 198148 136144
rect 198648 136060 198700 136066
rect 198648 136002 198700 136008
rect 198004 135652 198056 135658
rect 198004 135594 198056 135600
rect 197268 5500 197320 5506
rect 197268 5442 197320 5448
rect 198016 4690 198044 135594
rect 198004 4684 198056 4690
rect 198004 4626 198056 4632
rect 196348 3800 196400 3806
rect 196348 3742 196400 3748
rect 196808 3732 196860 3738
rect 196808 3674 196860 3680
rect 195612 3664 195664 3670
rect 195612 3606 195664 3612
rect 192944 3460 192996 3466
rect 192944 3402 192996 3408
rect 194416 3460 194468 3466
rect 194416 3402 194468 3408
rect 195244 3460 195296 3466
rect 195244 3402 195296 3408
rect 193220 3120 193272 3126
rect 193220 3062 193272 3068
rect 190828 3052 190880 3058
rect 190828 2994 190880 3000
rect 191748 3052 191800 3058
rect 191748 2994 191800 3000
rect 190840 480 190868 2994
rect 192024 2916 192076 2922
rect 192024 2858 192076 2864
rect 192036 480 192064 2858
rect 193232 480 193260 3062
rect 194428 480 194456 3402
rect 195624 480 195652 3606
rect 196820 480 196848 3674
rect 198660 3466 198688 136002
rect 198936 3806 198964 138366
rect 199384 135720 199436 135726
rect 199384 135662 199436 135668
rect 198924 3800 198976 3806
rect 198924 3742 198976 3748
rect 199396 3670 199424 135662
rect 199856 135658 199884 138366
rect 200684 136270 200712 138366
rect 200672 136264 200724 136270
rect 200672 136206 200724 136212
rect 199844 135652 199896 135658
rect 199844 135594 199896 135600
rect 200764 135652 200816 135658
rect 200764 135594 200816 135600
rect 200776 4622 200804 135594
rect 201512 16574 201540 138366
rect 202432 135658 202460 138366
rect 203260 136406 203288 138366
rect 203248 136400 203300 136406
rect 203248 136342 203300 136348
rect 202788 136264 202840 136270
rect 202788 136206 202840 136212
rect 202696 136128 202748 136134
rect 202696 136070 202748 136076
rect 202420 135652 202472 135658
rect 202420 135594 202472 135600
rect 201512 16546 201632 16574
rect 200764 4616 200816 4622
rect 200764 4558 200816 4564
rect 200304 3732 200356 3738
rect 200304 3674 200356 3680
rect 199384 3664 199436 3670
rect 199384 3606 199436 3612
rect 197912 3460 197964 3466
rect 197912 3402 197964 3408
rect 198648 3460 198700 3466
rect 198648 3402 198700 3408
rect 197924 480 197952 3402
rect 199108 3052 199160 3058
rect 199108 2994 199160 3000
rect 199120 480 199148 2994
rect 200316 480 200344 3674
rect 201604 3602 201632 16546
rect 201592 3596 201644 3602
rect 201592 3538 201644 3544
rect 201500 3528 201552 3534
rect 201500 3470 201552 3476
rect 201512 480 201540 3470
rect 202708 480 202736 136070
rect 202800 3534 202828 136206
rect 204088 3942 204116 138366
rect 204904 136400 204956 136406
rect 204904 136342 204956 136348
rect 204076 3936 204128 3942
rect 204076 3878 204128 3884
rect 204916 3534 204944 136342
rect 205008 135794 205036 138366
rect 205836 136474 205864 138366
rect 205824 136468 205876 136474
rect 205824 136410 205876 136416
rect 205548 136196 205600 136202
rect 205548 136138 205600 136144
rect 204996 135788 205048 135794
rect 204996 135730 205048 135736
rect 205560 3534 205588 136138
rect 206756 4010 206784 138366
rect 206928 135652 206980 135658
rect 206928 135594 206980 135600
rect 206744 4004 206796 4010
rect 206744 3946 206796 3952
rect 206940 3534 206968 135594
rect 207584 4146 207612 138366
rect 208412 135862 208440 138366
rect 209332 136542 209360 138366
rect 209320 136536 209372 136542
rect 209320 136478 209372 136484
rect 208400 135856 208452 135862
rect 208400 135798 208452 135804
rect 209688 135856 209740 135862
rect 209688 135798 209740 135804
rect 207572 4140 207624 4146
rect 207572 4082 207624 4088
rect 207388 3596 207440 3602
rect 207388 3538 207440 3544
rect 202788 3528 202840 3534
rect 202788 3470 202840 3476
rect 203892 3528 203944 3534
rect 203892 3470 203944 3476
rect 204904 3528 204956 3534
rect 204904 3470 204956 3476
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 206192 3528 206244 3534
rect 206192 3470 206244 3476
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 203904 480 203932 3470
rect 205100 480 205128 3470
rect 206204 480 206232 3470
rect 207400 480 207428 3538
rect 209700 3534 209728 135798
rect 210160 3874 210188 138366
rect 210988 136610 211016 138366
rect 210976 136604 211028 136610
rect 210976 136546 211028 136552
rect 211068 136468 211120 136474
rect 211068 136410 211120 136416
rect 211080 6914 211108 136410
rect 210988 6886 211108 6914
rect 210148 3868 210200 3874
rect 210148 3810 210200 3816
rect 209780 3800 209832 3806
rect 209780 3742 209832 3748
rect 208584 3528 208636 3534
rect 208584 3470 208636 3476
rect 209688 3528 209740 3534
rect 209688 3470 209740 3476
rect 208596 480 208624 3470
rect 209792 480 209820 3742
rect 210988 480 211016 6886
rect 211908 3398 211936 138366
rect 212172 3528 212224 3534
rect 212172 3470 212224 3476
rect 211896 3392 211948 3398
rect 211896 3334 211948 3340
rect 212184 480 212212 3470
rect 212736 3330 212764 138366
rect 213184 135788 213236 135794
rect 213184 135730 213236 135736
rect 213196 3534 213224 135730
rect 213564 135590 213592 138366
rect 213828 136604 213880 136610
rect 213828 136546 213880 136552
rect 213552 135584 213604 135590
rect 213552 135526 213604 135532
rect 213840 3534 213868 136546
rect 214484 6914 214512 138366
rect 215208 136536 215260 136542
rect 215208 136478 215260 136484
rect 214392 6886 214512 6914
rect 213184 3528 213236 3534
rect 213184 3470 213236 3476
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213828 3528 213880 3534
rect 213828 3470 213880 3476
rect 212724 3324 212776 3330
rect 212724 3266 212776 3272
rect 213380 480 213408 3470
rect 214392 3262 214420 6886
rect 215220 3534 215248 136478
rect 214472 3528 214524 3534
rect 214472 3470 214524 3476
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 214380 3256 214432 3262
rect 214380 3198 214432 3204
rect 214484 480 214512 3470
rect 215404 2854 215432 138366
rect 216232 138366 216306 138394
rect 217060 138366 217134 138394
rect 217888 138366 217962 138394
rect 218808 138366 218882 138394
rect 219636 138366 219710 138394
rect 220464 138366 220538 138394
rect 221384 138366 221458 138394
rect 222212 138366 222286 138394
rect 223040 138366 223114 138394
rect 223960 138366 224034 138394
rect 224788 138366 224862 138394
rect 225708 138366 225782 138394
rect 226536 138366 226610 138394
rect 227364 138366 227438 138394
rect 228284 138366 228358 138394
rect 229112 138366 229186 138394
rect 229940 138366 230014 138394
rect 230860 138366 230934 138394
rect 231688 138366 231762 138394
rect 232516 138366 232590 138394
rect 233436 138366 233510 138394
rect 234264 138366 234338 138394
rect 235092 138366 235166 138394
rect 236012 138366 236086 138394
rect 236840 138366 236914 138394
rect 237760 138366 237834 138394
rect 238588 138366 238662 138394
rect 239416 138366 239490 138394
rect 240336 138366 240410 138394
rect 241164 138366 241238 138394
rect 241992 138366 242066 138394
rect 242912 138366 242986 138394
rect 243740 138366 243814 138394
rect 244568 138366 244642 138394
rect 245488 138366 245562 138394
rect 246316 138366 246390 138394
rect 247236 138366 247310 138394
rect 248064 138366 248138 138394
rect 248892 138366 248966 138394
rect 249812 138366 249886 138394
rect 250640 138366 250714 138394
rect 251468 138366 251542 138394
rect 252388 138366 252462 138394
rect 253216 138366 253290 138394
rect 254044 138366 254118 138394
rect 254964 138366 255038 138394
rect 255792 138366 255866 138394
rect 256712 138366 256786 138394
rect 257540 138366 257614 138394
rect 258368 138366 258442 138394
rect 259288 138366 259362 138394
rect 260116 138366 260190 138394
rect 260944 138366 261018 138394
rect 261864 138366 261938 138394
rect 262692 138366 262766 138394
rect 263520 138366 263594 138394
rect 264440 138366 264514 138394
rect 265268 138366 265342 138394
rect 266096 138366 266170 138394
rect 267016 138366 267090 138394
rect 267844 138366 267918 138394
rect 268764 138366 268838 138394
rect 269592 138366 269666 138394
rect 270420 138366 270494 138394
rect 271340 138366 271414 138394
rect 272168 138366 272242 138394
rect 272996 138366 273070 138394
rect 273916 138366 273990 138394
rect 274744 138366 274818 138394
rect 275572 138366 275646 138394
rect 276492 138366 276566 138394
rect 277320 138366 277394 138394
rect 278240 138366 278314 138394
rect 279068 138366 279142 138394
rect 279896 138366 279970 138394
rect 280172 138366 280890 138394
rect 281644 138366 281718 138394
rect 282472 138366 282546 138394
rect 283392 138366 283466 138394
rect 284220 138366 284294 138394
rect 285048 138366 285122 138394
rect 285968 138366 286042 138394
rect 286796 138366 286870 138394
rect 287716 138366 287790 138394
rect 288544 138366 288618 138394
rect 289372 138366 289446 138394
rect 290292 138366 290366 138394
rect 291120 138366 291194 138394
rect 291948 138366 292022 138394
rect 292868 138366 292942 138394
rect 293696 138366 293770 138394
rect 294524 138366 294598 138394
rect 295352 138366 295518 138394
rect 296318 138394 296346 138652
rect 297146 138394 297174 138652
rect 298066 138394 298094 138652
rect 296318 138366 296668 138394
rect 297146 138366 297220 138394
rect 216232 136338 216260 138366
rect 216220 136332 216272 136338
rect 216220 136274 216272 136280
rect 216588 136332 216640 136338
rect 216588 136274 216640 136280
rect 216600 3534 216628 136274
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 216864 3528 216916 3534
rect 216864 3470 216916 3476
rect 215392 2848 215444 2854
rect 215392 2790 215444 2796
rect 215680 480 215708 3470
rect 216876 480 216904 3470
rect 217060 3466 217088 138366
rect 217048 3460 217100 3466
rect 217048 3402 217100 3408
rect 217888 3194 217916 138366
rect 218808 135930 218836 138366
rect 218796 135924 218848 135930
rect 218796 135866 218848 135872
rect 217968 135584 218020 135590
rect 217968 135526 218020 135532
rect 217980 3534 218008 135526
rect 219348 135448 219400 135454
rect 219348 135390 219400 135396
rect 219360 3534 219388 135390
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 219348 3528 219400 3534
rect 219348 3470 219400 3476
rect 217876 3188 217928 3194
rect 217876 3130 217928 3136
rect 218072 480 218100 3470
rect 219256 3392 219308 3398
rect 219256 3334 219308 3340
rect 219268 480 219296 3334
rect 219636 2922 219664 138366
rect 220084 135720 220136 135726
rect 220084 135662 220136 135668
rect 220096 3058 220124 135662
rect 220084 3052 220136 3058
rect 220084 2994 220136 3000
rect 220464 2990 220492 138366
rect 221384 135998 221412 138366
rect 221372 135992 221424 135998
rect 221372 135934 221424 135940
rect 222212 135930 222240 138366
rect 222200 135924 222252 135930
rect 222200 135866 222252 135872
rect 220728 135516 220780 135522
rect 220728 135458 220780 135464
rect 220740 6914 220768 135458
rect 220556 6886 220768 6914
rect 220452 2984 220504 2990
rect 220452 2926 220504 2932
rect 219624 2916 219676 2922
rect 219624 2858 219676 2864
rect 220556 2802 220584 6886
rect 223040 3670 223068 138366
rect 223960 136066 223988 138366
rect 223948 136060 224000 136066
rect 223948 136002 224000 136008
rect 223488 135992 223540 135998
rect 223488 135934 223540 135940
rect 223028 3664 223080 3670
rect 223028 3606 223080 3612
rect 221556 3596 221608 3602
rect 221556 3538 221608 3544
rect 220464 2774 220584 2802
rect 220464 480 220492 2774
rect 221568 480 221596 3538
rect 223500 3534 223528 135934
rect 224788 135726 224816 138366
rect 224868 136060 224920 136066
rect 224868 136002 224920 136008
rect 224776 135720 224828 135726
rect 224776 135662 224828 135668
rect 224224 135516 224276 135522
rect 224224 135458 224276 135464
rect 224236 3874 224264 135458
rect 224224 3868 224276 3874
rect 224224 3810 224276 3816
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 222764 480 222792 3470
rect 224880 3262 224908 136002
rect 225708 3738 225736 138366
rect 226536 136270 226564 138366
rect 226524 136264 226576 136270
rect 226524 136206 226576 136212
rect 227364 136134 227392 138366
rect 228284 136406 228312 138366
rect 228272 136400 228324 136406
rect 228272 136342 228324 136348
rect 229008 136400 229060 136406
rect 229008 136342 229060 136348
rect 227628 136264 227680 136270
rect 227628 136206 227680 136212
rect 227352 136128 227404 136134
rect 227352 136070 227404 136076
rect 227536 136128 227588 136134
rect 227536 136070 227588 136076
rect 226248 135720 226300 135726
rect 226248 135662 226300 135668
rect 225696 3732 225748 3738
rect 225696 3674 225748 3680
rect 226260 3534 226288 135662
rect 225144 3528 225196 3534
rect 225144 3470 225196 3476
rect 226248 3528 226300 3534
rect 226248 3470 226300 3476
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 223948 3256 224000 3262
rect 223948 3198 224000 3204
rect 224868 3256 224920 3262
rect 224868 3198 224920 3204
rect 223960 480 223988 3198
rect 225156 480 225184 3470
rect 226352 480 226380 3470
rect 227548 480 227576 136070
rect 227640 3534 227668 136206
rect 228364 135380 228416 135386
rect 228364 135322 228416 135328
rect 228376 3602 228404 135322
rect 229020 6914 229048 136342
rect 229112 136202 229140 138366
rect 229100 136196 229152 136202
rect 229100 136138 229152 136144
rect 229940 135658 229968 138366
rect 229928 135652 229980 135658
rect 229928 135594 229980 135600
rect 228744 6886 229048 6914
rect 228364 3596 228416 3602
rect 228364 3538 228416 3544
rect 227628 3528 227680 3534
rect 227628 3470 227680 3476
rect 228744 480 228772 6886
rect 230860 3806 230888 138366
rect 231688 135862 231716 138366
rect 231676 135856 231728 135862
rect 231676 135798 231728 135804
rect 231768 135856 231820 135862
rect 231768 135798 231820 135804
rect 231124 135312 231176 135318
rect 231124 135254 231176 135260
rect 230848 3800 230900 3806
rect 230848 3742 230900 3748
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 229836 3324 229888 3330
rect 229836 3266 229888 3272
rect 229848 480 229876 3266
rect 231044 480 231072 3470
rect 231136 3466 231164 135254
rect 231780 3534 231808 135798
rect 232516 135522 232544 138366
rect 233436 136474 233464 138366
rect 233424 136468 233476 136474
rect 233424 136410 233476 136416
rect 234264 135794 234292 138366
rect 235092 136610 235120 138366
rect 235080 136604 235132 136610
rect 235080 136546 235132 136552
rect 236012 136542 236040 138366
rect 236000 136536 236052 136542
rect 236000 136478 236052 136484
rect 235908 136468 235960 136474
rect 235908 136410 235960 136416
rect 234528 136196 234580 136202
rect 234528 136138 234580 136144
rect 234252 135788 234304 135794
rect 234252 135730 234304 135736
rect 233148 135652 233200 135658
rect 233148 135594 233200 135600
rect 232504 135516 232556 135522
rect 232504 135458 232556 135464
rect 233160 3534 233188 135594
rect 233884 135516 233936 135522
rect 233884 135458 233936 135464
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 231124 3460 231176 3466
rect 231124 3402 231176 3408
rect 232240 480 232268 3470
rect 233436 480 233464 3470
rect 233896 3330 233924 135458
rect 234540 3534 234568 136138
rect 235920 6914 235948 136410
rect 236840 136338 236868 138366
rect 236828 136332 236880 136338
rect 236828 136274 236880 136280
rect 237288 136332 237340 136338
rect 237288 136274 237340 136280
rect 237300 6914 237328 136274
rect 237760 135590 237788 138366
rect 238024 136604 238076 136610
rect 238024 136546 238076 136552
rect 237748 135584 237800 135590
rect 237748 135526 237800 135532
rect 235828 6886 235948 6914
rect 237024 6886 237328 6914
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 233884 3324 233936 3330
rect 233884 3266 233936 3272
rect 234620 3324 234672 3330
rect 234620 3266 234672 3272
rect 234632 480 234660 3266
rect 235828 480 235856 6886
rect 237024 480 237052 6886
rect 238036 3330 238064 136546
rect 238588 135454 238616 138366
rect 238668 136536 238720 136542
rect 238668 136478 238720 136484
rect 238576 135448 238628 135454
rect 238576 135390 238628 135396
rect 238680 3534 238708 136478
rect 239416 135318 239444 138366
rect 240336 135930 240364 138366
rect 240324 135924 240376 135930
rect 240324 135866 240376 135872
rect 241164 135386 241192 138366
rect 241992 135998 242020 138366
rect 242912 136066 242940 138366
rect 242900 136060 242952 136066
rect 242900 136002 242952 136008
rect 241980 135992 242032 135998
rect 241980 135934 242032 135940
rect 242808 135992 242860 135998
rect 242808 135934 242860 135940
rect 241428 135924 241480 135930
rect 241428 135866 241480 135872
rect 241152 135380 241204 135386
rect 241152 135322 241204 135328
rect 239404 135312 239456 135318
rect 239404 135254 239456 135260
rect 241440 3534 241468 135866
rect 238116 3528 238168 3534
rect 238116 3470 238168 3476
rect 238668 3528 238720 3534
rect 238668 3470 238720 3476
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 238024 3324 238076 3330
rect 238024 3266 238076 3272
rect 238128 480 238156 3470
rect 239312 3120 239364 3126
rect 239312 3062 239364 3068
rect 239324 480 239352 3062
rect 240520 480 240548 3470
rect 242820 3262 242848 135934
rect 243740 135726 243768 138366
rect 244568 136270 244596 138366
rect 244556 136264 244608 136270
rect 244556 136206 244608 136212
rect 245488 136134 245516 138366
rect 246316 136406 246344 138366
rect 246304 136400 246356 136406
rect 246304 136342 246356 136348
rect 246948 136264 247000 136270
rect 246948 136206 247000 136212
rect 245476 136128 245528 136134
rect 245476 136070 245528 136076
rect 245568 136060 245620 136066
rect 245568 136002 245620 136008
rect 243728 135720 243780 135726
rect 243728 135662 243780 135668
rect 244096 3460 244148 3466
rect 244096 3402 244148 3408
rect 241704 3256 241756 3262
rect 241704 3198 241756 3204
rect 242808 3256 242860 3262
rect 242808 3198 242860 3204
rect 242900 3256 242952 3262
rect 242900 3198 242952 3204
rect 241716 480 241744 3198
rect 242912 480 242940 3198
rect 244108 480 244136 3402
rect 245212 598 245424 626
rect 245212 480 245240 598
rect 245396 490 245424 598
rect 245580 490 245608 136002
rect 246304 135788 246356 135794
rect 246304 135730 246356 135736
rect 246316 3126 246344 135730
rect 246960 3330 246988 136206
rect 247236 135522 247264 138366
rect 248064 135862 248092 138366
rect 248052 135856 248104 135862
rect 248052 135798 248104 135804
rect 248892 135658 248920 138366
rect 249812 136202 249840 138366
rect 250640 136610 250668 138366
rect 250628 136604 250680 136610
rect 250628 136546 250680 136552
rect 251468 136474 251496 138366
rect 251456 136468 251508 136474
rect 251456 136410 251508 136416
rect 251088 136400 251140 136406
rect 251088 136342 251140 136348
rect 249800 136196 249852 136202
rect 249800 136138 249852 136144
rect 249708 136128 249760 136134
rect 249708 136070 249760 136076
rect 248880 135652 248932 135658
rect 248880 135594 248932 135600
rect 249064 135584 249116 135590
rect 249064 135526 249116 135532
rect 247224 135516 247276 135522
rect 247224 135458 247276 135464
rect 247592 3596 247644 3602
rect 247592 3538 247644 3544
rect 246396 3324 246448 3330
rect 246396 3266 246448 3272
rect 246948 3324 247000 3330
rect 246948 3266 247000 3272
rect 246304 3120 246356 3126
rect 246304 3062 246356 3068
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245396 462 245608 490
rect 246408 480 246436 3266
rect 247604 480 247632 3538
rect 248788 3528 248840 3534
rect 248788 3470 248840 3476
rect 248800 480 248828 3470
rect 249076 3330 249104 135526
rect 249720 3534 249748 136070
rect 251100 3534 251128 136342
rect 252388 136338 252416 138366
rect 253216 136542 253244 138366
rect 253204 136536 253256 136542
rect 253204 136478 253256 136484
rect 252376 136332 252428 136338
rect 252376 136274 252428 136280
rect 253848 136332 253900 136338
rect 253848 136274 253900 136280
rect 252468 136196 252520 136202
rect 252468 136138 252520 136144
rect 251824 135720 251876 135726
rect 251824 135662 251876 135668
rect 251836 3602 251864 135662
rect 251916 135516 251968 135522
rect 251916 135458 251968 135464
rect 251824 3596 251876 3602
rect 251824 3538 251876 3544
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 249064 3324 249116 3330
rect 249064 3266 249116 3272
rect 249996 480 250024 3470
rect 251192 480 251220 3470
rect 251928 3466 251956 135458
rect 252480 3534 252508 136138
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 251916 3460 251968 3466
rect 251916 3402 251968 3408
rect 252376 3324 252428 3330
rect 252376 3266 252428 3272
rect 252388 480 252416 3266
rect 253492 598 253704 626
rect 253492 480 253520 598
rect 253676 490 253704 598
rect 253860 490 253888 136274
rect 254044 135794 254072 138366
rect 254964 135930 254992 138366
rect 255792 135998 255820 138366
rect 255964 136536 256016 136542
rect 255964 136478 256016 136484
rect 255780 135992 255832 135998
rect 255780 135934 255832 135940
rect 254952 135924 255004 135930
rect 254952 135866 255004 135872
rect 255228 135924 255280 135930
rect 255228 135866 255280 135872
rect 254032 135788 254084 135794
rect 254032 135730 254084 135736
rect 255240 3534 255268 135866
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 255228 3528 255280 3534
rect 255228 3470 255280 3476
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 253676 462 253888 490
rect 254688 480 254716 3470
rect 255884 480 255912 3470
rect 255976 3330 256004 136478
rect 256608 136468 256660 136474
rect 256608 136410 256660 136416
rect 256620 3534 256648 136410
rect 256712 135590 256740 138366
rect 256700 135584 256752 135590
rect 256700 135526 256752 135532
rect 257540 135522 257568 138366
rect 258368 136066 258396 138366
rect 259288 136270 259316 138366
rect 259276 136264 259328 136270
rect 259276 136206 259328 136212
rect 258356 136060 258408 136066
rect 258356 136002 258408 136008
rect 259368 136060 259420 136066
rect 259368 136002 259420 136008
rect 257528 135516 257580 135522
rect 257528 135458 257580 135464
rect 259380 3534 259408 136002
rect 260116 135726 260144 138366
rect 260944 136134 260972 138366
rect 261864 136406 261892 138366
rect 261852 136400 261904 136406
rect 261852 136342 261904 136348
rect 262692 136202 262720 138366
rect 263520 136542 263548 138366
rect 263508 136536 263560 136542
rect 263508 136478 263560 136484
rect 264440 136338 264468 138366
rect 264428 136332 264480 136338
rect 264428 136274 264480 136280
rect 263508 136264 263560 136270
rect 263508 136206 263560 136212
rect 262680 136196 262732 136202
rect 262680 136138 262732 136144
rect 260932 136128 260984 136134
rect 260932 136070 260984 136076
rect 260748 135924 260800 135930
rect 260748 135866 260800 135872
rect 260656 135856 260708 135862
rect 260656 135798 260708 135804
rect 260104 135720 260156 135726
rect 260104 135662 260156 135668
rect 256608 3528 256660 3534
rect 256608 3470 256660 3476
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 257068 3460 257120 3466
rect 257068 3402 257120 3408
rect 255964 3324 256016 3330
rect 255964 3266 256016 3272
rect 257080 480 257108 3402
rect 258276 480 258304 3470
rect 259472 480 259500 3470
rect 260668 480 260696 135798
rect 260760 3534 260788 135866
rect 263520 3534 263548 136206
rect 264244 136196 264296 136202
rect 264244 136138 264296 136144
rect 260748 3528 260800 3534
rect 260748 3470 260800 3476
rect 262956 3528 263008 3534
rect 262956 3470 263008 3476
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 261760 3052 261812 3058
rect 261760 2994 261812 3000
rect 261772 480 261800 2994
rect 262968 480 262996 3470
rect 264164 480 264192 3470
rect 264256 3466 264284 136138
rect 264888 136128 264940 136134
rect 264888 136070 264940 136076
rect 264900 3534 264928 136070
rect 265268 135998 265296 138366
rect 266096 136474 266124 138366
rect 266084 136468 266136 136474
rect 266084 136410 266136 136416
rect 267016 136202 267044 138366
rect 267648 136332 267700 136338
rect 267648 136274 267700 136280
rect 267004 136196 267056 136202
rect 267004 136138 267056 136144
rect 265256 135992 265308 135998
rect 265256 135934 265308 135940
rect 267004 135992 267056 135998
rect 267004 135934 267056 135940
rect 264888 3528 264940 3534
rect 264888 3470 264940 3476
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 264244 3460 264296 3466
rect 264244 3402 264296 3408
rect 265348 3188 265400 3194
rect 265348 3130 265400 3136
rect 265360 480 265388 3130
rect 266556 480 266584 3470
rect 267016 3058 267044 135934
rect 267660 3534 267688 136274
rect 267844 136066 267872 138366
rect 268764 136270 268792 138366
rect 268752 136264 268804 136270
rect 268752 136206 268804 136212
rect 267832 136060 267884 136066
rect 267832 136002 267884 136008
rect 269592 135862 269620 138366
rect 270420 135998 270448 138366
rect 271340 136202 271368 138366
rect 271328 136196 271380 136202
rect 271328 136138 271380 136144
rect 272168 136134 272196 138366
rect 272156 136128 272208 136134
rect 272156 136070 272208 136076
rect 271788 136060 271840 136066
rect 271788 136002 271840 136008
rect 270408 135992 270460 135998
rect 270408 135934 270460 135940
rect 269580 135856 269632 135862
rect 269580 135798 269632 135804
rect 268936 135652 268988 135658
rect 268936 135594 268988 135600
rect 268948 3602 268976 135594
rect 269764 135584 269816 135590
rect 269764 135526 269816 135532
rect 269028 135516 269080 135522
rect 269028 135458 269080 135464
rect 267740 3596 267792 3602
rect 267740 3538 267792 3544
rect 268936 3596 268988 3602
rect 268936 3538 268988 3544
rect 267648 3528 267700 3534
rect 267648 3470 267700 3476
rect 267004 3052 267056 3058
rect 267004 2994 267056 3000
rect 267752 480 267780 3538
rect 269040 3482 269068 135458
rect 268856 3454 269068 3482
rect 268856 480 268884 3454
rect 269776 3194 269804 135526
rect 270408 135448 270460 135454
rect 270408 135390 270460 135396
rect 269764 3188 269816 3194
rect 269764 3130 269816 3136
rect 270052 598 270264 626
rect 270052 480 270080 598
rect 270236 490 270264 598
rect 270420 490 270448 135390
rect 271800 3330 271828 136002
rect 272996 135590 273024 138366
rect 273916 136338 273944 138366
rect 274548 136604 274600 136610
rect 274548 136546 274600 136552
rect 273904 136332 273956 136338
rect 273904 136274 273956 136280
rect 273904 136128 273956 136134
rect 273904 136070 273956 136076
rect 272984 135584 273036 135590
rect 272984 135526 273036 135532
rect 273628 3528 273680 3534
rect 273628 3470 273680 3476
rect 272432 3460 272484 3466
rect 272432 3402 272484 3408
rect 271236 3324 271288 3330
rect 271236 3266 271288 3272
rect 271788 3324 271840 3330
rect 271788 3266 271840 3272
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270236 462 270448 490
rect 271248 480 271276 3266
rect 272444 480 272472 3402
rect 273640 480 273668 3470
rect 273916 3466 273944 136070
rect 274560 3534 274588 136546
rect 274744 135658 274772 138366
rect 274732 135652 274784 135658
rect 274732 135594 274784 135600
rect 275572 135522 275600 138366
rect 275560 135516 275612 135522
rect 275560 135458 275612 135464
rect 276492 135454 276520 138366
rect 276664 136196 276716 136202
rect 276664 136138 276716 136144
rect 276480 135448 276532 135454
rect 276480 135390 276532 135396
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 273904 3460 273956 3466
rect 273904 3402 273956 3408
rect 276020 3460 276072 3466
rect 276020 3402 276072 3408
rect 274824 3052 274876 3058
rect 274824 2994 274876 3000
rect 274836 480 274864 2994
rect 276032 480 276060 3402
rect 276676 3058 276704 136138
rect 277320 136066 277348 138366
rect 278240 136134 278268 138366
rect 279068 136610 279096 138366
rect 279056 136604 279108 136610
rect 279056 136546 279108 136552
rect 279896 136202 279924 138366
rect 279884 136196 279936 136202
rect 279884 136138 279936 136144
rect 278228 136128 278280 136134
rect 278228 136070 278280 136076
rect 277308 136060 277360 136066
rect 277308 136002 277360 136008
rect 277308 135924 277360 135930
rect 277308 135866 277360 135872
rect 277320 6914 277348 135866
rect 278688 135516 278740 135522
rect 278688 135458 278740 135464
rect 277136 6886 277348 6914
rect 276664 3052 276716 3058
rect 276664 2994 276716 3000
rect 277136 480 277164 6886
rect 278332 598 278544 626
rect 278332 480 278360 598
rect 278516 490 278544 598
rect 278700 490 278728 135458
rect 279516 3528 279568 3534
rect 279516 3470 279568 3476
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 278516 462 278728 490
rect 279528 480 279556 3470
rect 280172 3466 280200 138366
rect 281644 135930 281672 138366
rect 281632 135924 281684 135930
rect 281632 135866 281684 135872
rect 280804 135652 280856 135658
rect 280804 135594 280856 135600
rect 280816 3534 280844 135594
rect 282184 135584 282236 135590
rect 282184 135526 282236 135532
rect 280804 3528 280856 3534
rect 280804 3470 280856 3476
rect 282196 3466 282224 135526
rect 282472 135522 282500 138366
rect 283392 135658 283420 138366
rect 283380 135652 283432 135658
rect 283380 135594 283432 135600
rect 284220 135590 284248 138366
rect 284208 135584 284260 135590
rect 284208 135526 284260 135532
rect 284944 135584 284996 135590
rect 284944 135526 284996 135532
rect 282460 135516 282512 135522
rect 282460 135458 282512 135464
rect 280160 3460 280212 3466
rect 280160 3402 280212 3408
rect 280712 3460 280764 3466
rect 280712 3402 280764 3408
rect 282184 3460 282236 3466
rect 282184 3402 282236 3408
rect 280724 480 280752 3402
rect 284300 3188 284352 3194
rect 284300 3130 284352 3136
rect 281908 3120 281960 3126
rect 281908 3062 281960 3068
rect 281920 480 281948 3062
rect 283104 3052 283156 3058
rect 283104 2994 283156 3000
rect 283116 480 283144 2994
rect 284312 480 284340 3130
rect 284956 3058 284984 135526
rect 285048 3126 285076 138366
rect 285968 135590 285996 138366
rect 285956 135584 286008 135590
rect 285956 135526 286008 135532
rect 285404 4140 285456 4146
rect 285404 4082 285456 4088
rect 285036 3120 285088 3126
rect 285036 3062 285088 3068
rect 284944 3052 284996 3058
rect 284944 2994 284996 3000
rect 285416 480 285444 4082
rect 286796 3194 286824 138366
rect 286968 136468 287020 136474
rect 286968 136410 287020 136416
rect 286784 3188 286836 3194
rect 286784 3130 286836 3136
rect 286612 598 286824 626
rect 286612 480 286640 598
rect 286796 490 286824 598
rect 286980 490 287008 136410
rect 287716 4146 287744 138366
rect 288544 136474 288572 138366
rect 288532 136468 288584 136474
rect 288532 136410 288584 136416
rect 289372 135590 289400 138366
rect 289820 135652 289872 135658
rect 289820 135594 289872 135600
rect 288348 135584 288400 135590
rect 288348 135526 288400 135532
rect 289360 135584 289412 135590
rect 289360 135526 289412 135532
rect 289728 135584 289780 135590
rect 289728 135526 289780 135532
rect 287704 4140 287756 4146
rect 287704 4082 287756 4088
rect 288360 3330 288388 135526
rect 289740 3534 289768 135526
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 287796 3324 287848 3330
rect 287796 3266 287848 3272
rect 288348 3324 288400 3330
rect 288348 3266 288400 3272
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 286796 462 287008 490
rect 287808 480 287836 3266
rect 289004 480 289032 3470
rect 289832 490 289860 135594
rect 290292 135590 290320 138366
rect 291120 135658 291148 138366
rect 291108 135652 291160 135658
rect 291108 135594 291160 135600
rect 290280 135584 290332 135590
rect 290280 135526 290332 135532
rect 291948 3534 291976 138366
rect 292580 135584 292632 135590
rect 292580 135526 292632 135532
rect 292592 3534 292620 135526
rect 292868 6914 292896 138366
rect 293696 135590 293724 138366
rect 293684 135584 293736 135590
rect 293684 135526 293736 135532
rect 294524 16574 294552 138366
rect 294524 16546 294920 16574
rect 292684 6886 292896 6914
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 291936 3528 291988 3534
rect 291936 3470 291988 3476
rect 292580 3528 292632 3534
rect 292580 3470 292632 3476
rect 290016 598 290228 626
rect 290016 490 290044 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 462 290044 490
rect 290200 480 290228 598
rect 291396 480 291424 3470
rect 292684 3346 292712 6886
rect 293684 3528 293736 3534
rect 293684 3470 293736 3476
rect 292592 3318 292712 3346
rect 292592 480 292620 3318
rect 293696 480 293724 3470
rect 294892 480 294920 16546
rect 295352 3534 295380 138366
rect 296640 4146 296668 138366
rect 297192 135658 297220 138366
rect 298020 138366 298094 138394
rect 298894 138394 298922 138652
rect 299814 138394 299842 138652
rect 300642 138394 300670 138652
rect 301470 138394 301498 138652
rect 302390 138394 302418 138652
rect 303218 138394 303246 138652
rect 304046 138394 304074 138652
rect 304966 138394 304994 138652
rect 298894 138366 298968 138394
rect 299814 138366 299888 138394
rect 300642 138366 300716 138394
rect 301470 138366 301544 138394
rect 302390 138366 302464 138394
rect 303218 138366 303292 138394
rect 304046 138366 304120 138394
rect 297180 135652 297232 135658
rect 297180 135594 297232 135600
rect 298020 135590 298048 138366
rect 298100 135652 298152 135658
rect 298100 135594 298152 135600
rect 298008 135584 298060 135590
rect 298008 135526 298060 135532
rect 296628 4140 296680 4146
rect 296628 4082 296680 4088
rect 297272 4140 297324 4146
rect 297272 4082 297324 4088
rect 295340 3528 295392 3534
rect 295340 3470 295392 3476
rect 296076 3528 296128 3534
rect 296076 3470 296128 3476
rect 296088 480 296116 3470
rect 297284 480 297312 4082
rect 298112 490 298140 135594
rect 298940 135590 298968 138366
rect 299860 135590 299888 138366
rect 300688 135658 300716 138366
rect 300676 135652 300728 135658
rect 300676 135594 300728 135600
rect 301516 135590 301544 138366
rect 302436 135658 302464 138366
rect 303264 136542 303292 138366
rect 303252 136536 303304 136542
rect 303252 136478 303304 136484
rect 302240 135652 302292 135658
rect 302240 135594 302292 135600
rect 302424 135652 302476 135658
rect 302424 135594 302476 135600
rect 298744 135584 298796 135590
rect 298744 135526 298796 135532
rect 298928 135584 298980 135590
rect 298928 135526 298980 135532
rect 299572 135584 299624 135590
rect 299572 135526 299624 135532
rect 299848 135584 299900 135590
rect 299848 135526 299900 135532
rect 300768 135584 300820 135590
rect 300768 135526 300820 135532
rect 301504 135584 301556 135590
rect 301504 135526 301556 135532
rect 298756 3534 298784 135526
rect 299584 16574 299612 135526
rect 299584 16546 300716 16574
rect 298744 3528 298796 3534
rect 298744 3470 298796 3476
rect 299664 3528 299716 3534
rect 299664 3470 299716 3476
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3470
rect 300688 3346 300716 16546
rect 300780 3534 300808 135526
rect 302252 16574 302280 135594
rect 304092 135590 304120 138366
rect 304920 138366 304994 138394
rect 305794 138394 305822 138652
rect 306622 138394 306650 138652
rect 307542 138394 307570 138652
rect 308370 138394 308398 138652
rect 309290 138394 309318 138652
rect 310118 138394 310146 138652
rect 310946 138394 310974 138652
rect 311866 138394 311894 138652
rect 305794 138366 305868 138394
rect 306622 138366 306696 138394
rect 307542 138366 307616 138394
rect 308370 138366 308444 138394
rect 309290 138366 309364 138394
rect 310118 138366 310468 138394
rect 310946 138366 311020 138394
rect 304920 135726 304948 138366
rect 305840 135998 305868 138366
rect 306564 136536 306616 136542
rect 306564 136478 306616 136484
rect 305828 135992 305880 135998
rect 305828 135934 305880 135940
rect 304908 135720 304960 135726
rect 304908 135662 304960 135668
rect 305644 135720 305696 135726
rect 305644 135662 305696 135668
rect 305000 135652 305052 135658
rect 305000 135594 305052 135600
rect 303620 135584 303672 135590
rect 303620 135526 303672 135532
rect 304080 135584 304132 135590
rect 304080 135526 304132 135532
rect 304908 135584 304960 135590
rect 304908 135526 304960 135532
rect 303632 16574 303660 135526
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 301964 3528 302016 3534
rect 301964 3470 302016 3476
rect 300688 3318 300808 3346
rect 300780 480 300808 3318
rect 301976 480 302004 3470
rect 303172 480 303200 16546
rect 303908 490 303936 16546
rect 304920 4146 304948 135526
rect 305012 16574 305040 135594
rect 305012 16546 305592 16574
rect 304908 4140 304960 4146
rect 304908 4082 304960 4088
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 16546
rect 305656 3942 305684 135662
rect 306576 16574 306604 136478
rect 306668 135590 306696 138366
rect 306656 135584 306708 135590
rect 306656 135526 306708 135532
rect 306576 16546 306788 16574
rect 305644 3936 305696 3942
rect 305644 3878 305696 3884
rect 306760 480 306788 16546
rect 307588 3466 307616 138366
rect 307668 135584 307720 135590
rect 307668 135526 307720 135532
rect 307576 3460 307628 3466
rect 307576 3402 307628 3408
rect 307680 3330 307708 135526
rect 308416 135522 308444 138366
rect 309232 135992 309284 135998
rect 309232 135934 309284 135940
rect 308404 135516 308456 135522
rect 308404 135458 308456 135464
rect 309244 132494 309272 135934
rect 309336 135590 309364 138366
rect 309324 135584 309376 135590
rect 309324 135526 309376 135532
rect 310336 135584 310388 135590
rect 310336 135526 310388 135532
rect 309244 132466 309364 132494
rect 309336 16574 309364 132466
rect 309336 16546 309824 16574
rect 307944 4140 307996 4146
rect 307944 4082 307996 4088
rect 307668 3324 307720 3330
rect 307668 3266 307720 3272
rect 307956 480 307984 4082
rect 309048 3936 309100 3942
rect 309048 3878 309100 3884
rect 309060 480 309088 3878
rect 309796 490 309824 16546
rect 310348 3534 310376 135526
rect 310336 3528 310388 3534
rect 310336 3470 310388 3476
rect 310440 3058 310468 138366
rect 310992 135590 311020 138366
rect 311820 138366 311894 138394
rect 312694 138394 312722 138652
rect 313522 138394 313550 138652
rect 314442 138394 314470 138652
rect 315270 138394 315298 138652
rect 316098 138394 316126 138652
rect 317018 138394 317046 138652
rect 317846 138394 317874 138652
rect 318766 138394 318794 138652
rect 312694 138366 312768 138394
rect 313522 138366 313596 138394
rect 314442 138366 314516 138394
rect 315270 138366 315344 138394
rect 316098 138366 316172 138394
rect 317018 138366 317092 138394
rect 317846 138366 317920 138394
rect 310980 135584 311032 135590
rect 310980 135526 311032 135532
rect 311716 135584 311768 135590
rect 311716 135526 311768 135532
rect 311440 3324 311492 3330
rect 311440 3266 311492 3272
rect 310428 3052 310480 3058
rect 310428 2994 310480 3000
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 3266
rect 311728 3194 311756 135526
rect 311820 4078 311848 138366
rect 312740 135590 312768 138366
rect 313568 135590 313596 138366
rect 314488 135998 314516 138366
rect 315316 136610 315344 138366
rect 315304 136604 315356 136610
rect 315304 136546 315356 136552
rect 314476 135992 314528 135998
rect 314476 135934 314528 135940
rect 316144 135590 316172 138366
rect 316684 136604 316736 136610
rect 316684 136546 316736 136552
rect 312728 135584 312780 135590
rect 312728 135526 312780 135532
rect 313188 135584 313240 135590
rect 313188 135526 313240 135532
rect 313556 135584 313608 135590
rect 313556 135526 313608 135532
rect 314568 135584 314620 135590
rect 314568 135526 314620 135532
rect 316132 135584 316184 135590
rect 316132 135526 316184 135532
rect 311808 4072 311860 4078
rect 311808 4014 311860 4020
rect 313200 3874 313228 135526
rect 313372 135516 313424 135522
rect 313372 135458 313424 135464
rect 313384 16574 313412 135458
rect 313384 16546 313872 16574
rect 313188 3868 313240 3874
rect 313188 3810 313240 3816
rect 312636 3460 312688 3466
rect 312636 3402 312688 3408
rect 311716 3188 311768 3194
rect 311716 3130 311768 3136
rect 312648 480 312676 3402
rect 313844 480 313872 16546
rect 314580 3738 314608 135526
rect 314568 3732 314620 3738
rect 314568 3674 314620 3680
rect 315028 3528 315080 3534
rect 315028 3470 315080 3476
rect 315040 480 315068 3470
rect 316696 3058 316724 136546
rect 317064 135522 317092 138366
rect 317892 135590 317920 138366
rect 318628 138366 318794 138394
rect 319594 138394 319622 138652
rect 320422 138394 320450 138652
rect 321342 138394 321370 138652
rect 322170 138394 322198 138652
rect 322998 138394 323026 138652
rect 323918 138394 323946 138652
rect 324746 138394 324774 138652
rect 325574 138394 325602 138652
rect 319594 138366 319668 138394
rect 320422 138366 320496 138394
rect 321342 138366 321416 138394
rect 322170 138366 322244 138394
rect 322998 138366 323072 138394
rect 323918 138366 324176 138394
rect 324746 138366 324820 138394
rect 317328 135584 317380 135590
rect 317328 135526 317380 135532
rect 317880 135584 317932 135590
rect 317880 135526 317932 135532
rect 317052 135516 317104 135522
rect 317052 135458 317104 135464
rect 317340 3466 317368 135526
rect 318524 4072 318576 4078
rect 318524 4014 318576 4020
rect 317328 3460 317380 3466
rect 317328 3402 317380 3408
rect 317328 3188 317380 3194
rect 317328 3130 317380 3136
rect 316224 3052 316276 3058
rect 316224 2994 316276 3000
rect 316684 3052 316736 3058
rect 316684 2994 316736 3000
rect 316236 480 316264 2994
rect 317340 480 317368 3130
rect 318536 480 318564 4014
rect 318628 3670 318656 138366
rect 319640 135590 319668 138366
rect 320468 135658 320496 138366
rect 320456 135652 320508 135658
rect 320456 135594 320508 135600
rect 318708 135584 318760 135590
rect 318708 135526 318760 135532
rect 319628 135584 319680 135590
rect 319628 135526 319680 135532
rect 320824 135584 320876 135590
rect 320824 135526 320876 135532
rect 318616 3664 318668 3670
rect 318616 3606 318668 3612
rect 318720 3602 318748 135526
rect 320836 16574 320864 135526
rect 320836 16546 321048 16574
rect 319720 3868 319772 3874
rect 319720 3810 319772 3816
rect 318708 3596 318760 3602
rect 318708 3538 318760 3544
rect 319732 480 319760 3810
rect 321020 3738 321048 16546
rect 320916 3732 320968 3738
rect 320916 3674 320968 3680
rect 321008 3732 321060 3738
rect 321008 3674 321060 3680
rect 320928 480 320956 3674
rect 321388 3534 321416 138366
rect 321652 135992 321704 135998
rect 321652 135934 321704 135940
rect 321468 135652 321520 135658
rect 321468 135594 321520 135600
rect 321480 3874 321508 135594
rect 321664 16574 321692 135934
rect 322216 135590 322244 138366
rect 323044 135590 323072 138366
rect 322204 135584 322256 135590
rect 322204 135526 322256 135532
rect 322848 135584 322900 135590
rect 322848 135526 322900 135532
rect 323032 135584 323084 135590
rect 323032 135526 323084 135532
rect 321664 16546 322152 16574
rect 321468 3868 321520 3874
rect 321468 3810 321520 3816
rect 321376 3528 321428 3534
rect 321376 3470 321428 3476
rect 322124 480 322152 16546
rect 322860 4078 322888 135526
rect 322848 4072 322900 4078
rect 322848 4014 322900 4020
rect 324148 4010 324176 138366
rect 324792 135590 324820 138366
rect 325528 138366 325602 138394
rect 326494 138394 326522 138652
rect 327322 138394 327350 138652
rect 328150 138394 328178 138652
rect 329070 138394 329098 138652
rect 329898 138394 329926 138652
rect 330818 138394 330846 138652
rect 331646 138394 331674 138652
rect 332474 138394 332502 138652
rect 333394 138394 333422 138652
rect 334222 138394 334250 138652
rect 335050 138394 335078 138652
rect 335970 138394 335998 138652
rect 336798 138394 336826 138652
rect 337626 138394 337654 138652
rect 338546 138394 338574 138652
rect 339374 138394 339402 138652
rect 326494 138366 326568 138394
rect 327322 138366 327396 138394
rect 328150 138366 328316 138394
rect 329070 138366 329144 138394
rect 329898 138366 329972 138394
rect 330818 138366 331168 138394
rect 331646 138366 331720 138394
rect 332474 138366 332548 138394
rect 333394 138366 333468 138394
rect 334222 138366 334296 138394
rect 335050 138366 335308 138394
rect 335970 138366 336044 138394
rect 336798 138366 336872 138394
rect 337626 138366 337700 138394
rect 338546 138366 338620 138394
rect 324228 135584 324280 135590
rect 324228 135526 324280 135532
rect 324780 135584 324832 135590
rect 324780 135526 324832 135532
rect 324136 4004 324188 4010
rect 324136 3946 324188 3952
rect 324240 3262 324268 135526
rect 324504 135516 324556 135522
rect 324504 135458 324556 135464
rect 324516 16574 324544 135458
rect 324516 16546 325464 16574
rect 324412 3460 324464 3466
rect 324412 3402 324464 3408
rect 324228 3256 324280 3262
rect 324228 3198 324280 3204
rect 323308 3052 323360 3058
rect 323308 2994 323360 3000
rect 323320 480 323348 2994
rect 324424 480 324452 3402
rect 325436 3210 325464 16546
rect 325528 3670 325556 138366
rect 326540 135590 326568 138366
rect 327368 135658 327396 138366
rect 327356 135652 327408 135658
rect 327356 135594 327408 135600
rect 325608 135584 325660 135590
rect 325608 135526 325660 135532
rect 326528 135584 326580 135590
rect 326528 135526 326580 135532
rect 327724 135584 327776 135590
rect 327724 135526 327776 135532
rect 325516 3664 325568 3670
rect 325516 3606 325568 3612
rect 325620 3330 325648 135526
rect 327736 3806 327764 135526
rect 327724 3800 327776 3806
rect 327724 3742 327776 3748
rect 328288 3602 328316 138366
rect 328368 135652 328420 135658
rect 328368 135594 328420 135600
rect 328380 3942 328408 135594
rect 329116 135590 329144 138366
rect 329944 135794 329972 138366
rect 329932 135788 329984 135794
rect 329932 135730 329984 135736
rect 329104 135584 329156 135590
rect 329104 135526 329156 135532
rect 329748 135584 329800 135590
rect 329748 135526 329800 135532
rect 328368 3936 328420 3942
rect 328368 3878 328420 3884
rect 329760 3738 329788 135526
rect 331140 3874 331168 138366
rect 331692 135590 331720 138366
rect 331680 135584 331732 135590
rect 331680 135526 331732 135532
rect 332416 135584 332468 135590
rect 332416 135526 332468 135532
rect 330392 3868 330444 3874
rect 330392 3810 330444 3816
rect 331128 3868 331180 3874
rect 331128 3810 331180 3816
rect 329196 3732 329248 3738
rect 329196 3674 329248 3680
rect 329748 3732 329800 3738
rect 329748 3674 329800 3680
rect 326804 3596 326856 3602
rect 326804 3538 326856 3544
rect 328276 3596 328328 3602
rect 328276 3538 328328 3544
rect 325608 3324 325660 3330
rect 325608 3266 325660 3272
rect 325436 3182 325648 3210
rect 325620 480 325648 3182
rect 326816 480 326844 3538
rect 328000 3528 328052 3534
rect 328000 3470 328052 3476
rect 328012 480 328040 3470
rect 329208 480 329236 3674
rect 330404 480 330432 3810
rect 332428 3534 332456 135526
rect 332416 3528 332468 3534
rect 332416 3470 332468 3476
rect 331588 3460 331640 3466
rect 331588 3402 331640 3408
rect 331600 480 331628 3402
rect 332520 3398 332548 138366
rect 333440 135930 333468 138366
rect 333428 135924 333480 135930
rect 333428 135866 333480 135872
rect 334268 135590 334296 138366
rect 334256 135584 334308 135590
rect 334256 135526 334308 135532
rect 335176 135584 335228 135590
rect 335176 135526 335228 135532
rect 332692 4072 332744 4078
rect 332692 4014 332744 4020
rect 332508 3392 332560 3398
rect 332508 3334 332560 3340
rect 332704 480 332732 4014
rect 335084 4004 335136 4010
rect 335084 3946 335136 3952
rect 333888 3256 333940 3262
rect 333888 3198 333940 3204
rect 333900 480 333928 3198
rect 335096 480 335124 3946
rect 335188 3466 335216 135526
rect 335280 4146 335308 138366
rect 336016 135998 336044 138366
rect 336004 135992 336056 135998
rect 336004 135934 336056 135940
rect 336648 135992 336700 135998
rect 336648 135934 336700 135940
rect 336096 135924 336148 135930
rect 336096 135866 336148 135872
rect 336004 135788 336056 135794
rect 336004 135730 336056 135736
rect 335268 4140 335320 4146
rect 335268 4082 335320 4088
rect 335176 3460 335228 3466
rect 335176 3402 335228 3408
rect 336016 3058 336044 135730
rect 336108 3126 336136 135866
rect 336660 4010 336688 135934
rect 336844 135590 336872 138366
rect 336832 135584 336884 135590
rect 336832 135526 336884 135532
rect 337672 135522 337700 138366
rect 338592 135658 338620 138366
rect 339328 138366 339402 138394
rect 340294 138394 340322 138652
rect 341122 138394 341150 138652
rect 341950 138394 341978 138652
rect 342870 138394 342898 138652
rect 343698 138394 343726 138652
rect 344526 138394 344554 138652
rect 345446 138394 345474 138652
rect 346274 138394 346302 138652
rect 340294 138366 340368 138394
rect 341122 138366 341196 138394
rect 341950 138366 342116 138394
rect 342870 138366 342944 138394
rect 343698 138366 343772 138394
rect 344526 138366 344876 138394
rect 345446 138366 345520 138394
rect 338580 135652 338632 135658
rect 338580 135594 338632 135600
rect 338764 135584 338816 135590
rect 338764 135526 338816 135532
rect 337660 135516 337712 135522
rect 337660 135458 337712 135464
rect 336648 4004 336700 4010
rect 336648 3946 336700 3952
rect 338672 3800 338724 3806
rect 338672 3742 338724 3748
rect 337476 3664 337528 3670
rect 337476 3606 337528 3612
rect 336280 3324 336332 3330
rect 336280 3266 336332 3272
rect 336096 3120 336148 3126
rect 336096 3062 336148 3068
rect 336004 3052 336056 3058
rect 336004 2994 336056 3000
rect 336292 480 336320 3266
rect 337488 480 337516 3606
rect 338684 480 338712 3742
rect 338776 3126 338804 135526
rect 339328 3670 339356 138366
rect 339408 135652 339460 135658
rect 339408 135594 339460 135600
rect 339420 3806 339448 135594
rect 340340 135590 340368 138366
rect 341168 135590 341196 138366
rect 340328 135584 340380 135590
rect 340328 135526 340380 135532
rect 340788 135584 340840 135590
rect 340788 135526 340840 135532
rect 341156 135584 341208 135590
rect 341156 135526 341208 135532
rect 340144 135516 340196 135522
rect 340144 135458 340196 135464
rect 339868 3936 339920 3942
rect 339868 3878 339920 3884
rect 339408 3800 339460 3806
rect 339408 3742 339460 3748
rect 339316 3664 339368 3670
rect 339316 3606 339368 3612
rect 338764 3120 338816 3126
rect 338764 3062 338816 3068
rect 339880 480 339908 3878
rect 340156 2854 340184 135458
rect 340800 3942 340828 135526
rect 340788 3936 340840 3942
rect 340788 3878 340840 3884
rect 342088 3738 342116 138366
rect 342916 135590 342944 138366
rect 343744 135590 343772 138366
rect 342168 135584 342220 135590
rect 342168 135526 342220 135532
rect 342904 135584 342956 135590
rect 342904 135526 342956 135532
rect 343548 135584 343600 135590
rect 343548 135526 343600 135532
rect 343732 135584 343784 135590
rect 343732 135526 343784 135532
rect 342180 4078 342208 135526
rect 342168 4072 342220 4078
rect 342168 4014 342220 4020
rect 342076 3732 342128 3738
rect 342076 3674 342128 3680
rect 342168 3664 342220 3670
rect 342168 3606 342220 3612
rect 340972 3596 341024 3602
rect 340972 3538 341024 3544
rect 340144 2848 340196 2854
rect 340144 2790 340196 2796
rect 340984 480 341012 3538
rect 342180 480 342208 3606
rect 343364 3052 343416 3058
rect 343364 2994 343416 3000
rect 343376 480 343404 2994
rect 343560 2990 343588 135526
rect 344560 3868 344612 3874
rect 344560 3810 344612 3816
rect 343548 2984 343600 2990
rect 343548 2926 343600 2932
rect 344572 480 344600 3810
rect 344848 3602 344876 138366
rect 345492 135590 345520 138366
rect 346228 138366 346302 138394
rect 347102 138394 347130 138652
rect 348022 138394 348050 138652
rect 348850 138394 348878 138652
rect 349770 138394 349798 138652
rect 350598 138394 350626 138652
rect 351426 138394 351454 138652
rect 352346 138394 352374 138652
rect 353174 138394 353202 138652
rect 354002 138394 354030 138652
rect 354922 138394 354950 138652
rect 355750 138394 355778 138652
rect 356578 138394 356606 138652
rect 357498 138394 357526 138652
rect 358326 138394 358354 138652
rect 359154 138394 359182 138652
rect 360074 138394 360102 138652
rect 347102 138366 347176 138394
rect 348022 138366 348096 138394
rect 348850 138366 349016 138394
rect 349770 138366 349844 138394
rect 350598 138366 350672 138394
rect 351426 138366 351868 138394
rect 352346 138366 352420 138394
rect 353174 138366 353248 138394
rect 354002 138366 354076 138394
rect 354922 138366 354996 138394
rect 355750 138366 356008 138394
rect 356578 138366 356652 138394
rect 357498 138366 357572 138394
rect 358326 138366 358768 138394
rect 359154 138366 359228 138394
rect 344928 135584 344980 135590
rect 344928 135526 344980 135532
rect 345480 135584 345532 135590
rect 345480 135526 345532 135532
rect 344836 3596 344888 3602
rect 344836 3538 344888 3544
rect 344940 2922 344968 135526
rect 346228 3534 346256 138366
rect 347148 135590 347176 138366
rect 348068 135590 348096 138366
rect 346308 135584 346360 135590
rect 346308 135526 346360 135532
rect 347136 135584 347188 135590
rect 347136 135526 347188 135532
rect 347688 135584 347740 135590
rect 347688 135526 347740 135532
rect 348056 135584 348108 135590
rect 348056 135526 348108 135532
rect 346320 3874 346348 135526
rect 346308 3868 346360 3874
rect 346308 3810 346360 3816
rect 345756 3528 345808 3534
rect 345756 3470 345808 3476
rect 346216 3528 346268 3534
rect 346216 3470 346268 3476
rect 344928 2916 344980 2922
rect 344928 2858 344980 2864
rect 345768 480 345796 3470
rect 346952 3392 347004 3398
rect 346952 3334 347004 3340
rect 346964 480 346992 3334
rect 347700 3058 347728 135526
rect 348056 3324 348108 3330
rect 348056 3266 348108 3272
rect 347688 3052 347740 3058
rect 347688 2994 347740 3000
rect 348068 480 348096 3266
rect 348988 3126 349016 138366
rect 349816 135590 349844 138366
rect 350644 135590 350672 138366
rect 349068 135584 349120 135590
rect 349068 135526 349120 135532
rect 349804 135584 349856 135590
rect 349804 135526 349856 135532
rect 350448 135584 350500 135590
rect 350448 135526 350500 135532
rect 350632 135584 350684 135590
rect 350632 135526 350684 135532
rect 351736 135584 351788 135590
rect 351736 135526 351788 135532
rect 349080 3398 349108 135526
rect 350460 6914 350488 135526
rect 350368 6886 350488 6914
rect 349252 3460 349304 3466
rect 349252 3402 349304 3408
rect 349068 3392 349120 3398
rect 349068 3334 349120 3340
rect 348976 3120 349028 3126
rect 348976 3062 349028 3068
rect 349264 480 349292 3402
rect 350368 3194 350396 6886
rect 350448 4140 350500 4146
rect 350448 4082 350500 4088
rect 350356 3188 350408 3194
rect 350356 3130 350408 3136
rect 350460 480 350488 4082
rect 351644 4004 351696 4010
rect 351644 3946 351696 3952
rect 351656 480 351684 3946
rect 351748 3330 351776 135526
rect 351840 3466 351868 138366
rect 352392 135930 352420 138366
rect 352380 135924 352432 135930
rect 352380 135866 352432 135872
rect 353220 4146 353248 138366
rect 354048 135590 354076 138366
rect 354968 135658 354996 138366
rect 354956 135652 355008 135658
rect 354956 135594 355008 135600
rect 354036 135584 354088 135590
rect 354036 135526 354088 135532
rect 354588 135584 354640 135590
rect 354588 135526 354640 135532
rect 353208 4140 353260 4146
rect 353208 4082 353260 4088
rect 351828 3460 351880 3466
rect 351828 3402 351880 3408
rect 354600 3398 354628 135526
rect 355980 3806 356008 138366
rect 356624 135590 356652 138366
rect 356704 135652 356756 135658
rect 356704 135594 356756 135600
rect 356612 135584 356664 135590
rect 356612 135526 356664 135532
rect 356716 4962 356744 135594
rect 357544 135590 357572 138366
rect 357348 135584 357400 135590
rect 357348 135526 357400 135532
rect 357532 135584 357584 135590
rect 357532 135526 357584 135532
rect 358636 135584 358688 135590
rect 358636 135526 358688 135532
rect 356704 4956 356756 4962
rect 356704 4898 356756 4904
rect 357360 4010 357388 135526
rect 358648 7614 358676 135526
rect 358636 7608 358688 7614
rect 358636 7550 358688 7556
rect 358636 4072 358688 4078
rect 358636 4014 358688 4020
rect 357348 4004 357400 4010
rect 357348 3946 357400 3952
rect 357532 3936 357584 3942
rect 357532 3878 357584 3884
rect 355232 3800 355284 3806
rect 355232 3742 355284 3748
rect 355968 3800 356020 3806
rect 355968 3742 356020 3748
rect 354588 3392 354640 3398
rect 354588 3334 354640 3340
rect 351736 3324 351788 3330
rect 351736 3266 351788 3272
rect 352840 3256 352892 3262
rect 352840 3198 352892 3204
rect 352852 480 352880 3198
rect 354036 2848 354088 2854
rect 354036 2790 354088 2796
rect 354048 480 354076 2790
rect 355244 480 355272 3742
rect 356336 3664 356388 3670
rect 356336 3606 356388 3612
rect 356348 480 356376 3606
rect 357544 480 357572 3878
rect 358648 1578 358676 4014
rect 358740 3670 358768 138366
rect 359200 135590 359228 138366
rect 360028 138366 360102 138394
rect 360902 138394 360930 138652
rect 361822 138394 361850 138652
rect 362650 138394 362678 138652
rect 363478 138394 363506 138652
rect 364398 138394 364426 138652
rect 365226 138394 365254 138652
rect 366054 138394 366082 138652
rect 366974 138394 367002 138652
rect 360902 138366 360976 138394
rect 361822 138366 361896 138394
rect 362650 138366 362724 138394
rect 363478 138366 363552 138394
rect 364398 138366 364472 138394
rect 365226 138366 365300 138394
rect 366054 138366 366128 138394
rect 359188 135584 359240 135590
rect 359188 135526 359240 135532
rect 360028 4894 360056 138366
rect 360948 135590 360976 138366
rect 361868 135590 361896 138366
rect 362696 135658 362724 138366
rect 362684 135652 362736 135658
rect 362684 135594 362736 135600
rect 363524 135590 363552 138366
rect 363604 135652 363656 135658
rect 363604 135594 363656 135600
rect 360108 135584 360160 135590
rect 360108 135526 360160 135532
rect 360936 135584 360988 135590
rect 360936 135526 360988 135532
rect 361488 135584 361540 135590
rect 361488 135526 361540 135532
rect 361856 135584 361908 135590
rect 361856 135526 361908 135532
rect 362868 135584 362920 135590
rect 362868 135526 362920 135532
rect 363512 135584 363564 135590
rect 363512 135526 363564 135532
rect 360016 4888 360068 4894
rect 360016 4830 360068 4836
rect 360120 4078 360148 135526
rect 360108 4072 360160 4078
rect 360108 4014 360160 4020
rect 361500 3738 361528 135526
rect 362880 3942 362908 135526
rect 363616 8974 363644 135594
rect 364444 135590 364472 138366
rect 365272 135998 365300 138366
rect 365260 135992 365312 135998
rect 365260 135934 365312 135940
rect 366100 135590 366128 138366
rect 366928 138366 367002 138394
rect 367802 138394 367830 138652
rect 368630 138394 368658 138652
rect 369550 138394 369578 138652
rect 370378 138394 370406 138652
rect 371298 138394 371326 138652
rect 372126 138394 372154 138652
rect 372954 138394 372982 138652
rect 373874 138394 373902 138652
rect 374702 138394 374730 138652
rect 375530 138394 375558 138652
rect 376450 138394 376478 138652
rect 377278 138394 377306 138652
rect 378106 138394 378134 138652
rect 367802 138366 367876 138394
rect 368630 138366 368704 138394
rect 369550 138366 369716 138394
rect 370378 138366 370452 138394
rect 371298 138366 371372 138394
rect 372126 138366 372568 138394
rect 372954 138366 373028 138394
rect 373874 138366 373948 138394
rect 374702 138366 374776 138394
rect 375530 138366 375604 138394
rect 376450 138366 376708 138394
rect 377278 138366 377352 138394
rect 364248 135584 364300 135590
rect 364248 135526 364300 135532
rect 364432 135584 364484 135590
rect 364432 135526 364484 135532
rect 365628 135584 365680 135590
rect 365628 135526 365680 135532
rect 366088 135584 366140 135590
rect 366088 135526 366140 135532
rect 363604 8968 363656 8974
rect 363604 8910 363656 8916
rect 362868 3936 362920 3942
rect 362868 3878 362920 3884
rect 359924 3732 359976 3738
rect 359924 3674 359976 3680
rect 361488 3732 361540 3738
rect 361488 3674 361540 3680
rect 358728 3664 358780 3670
rect 358728 3606 358780 3612
rect 358648 1550 358768 1578
rect 358740 480 358768 1550
rect 359936 480 359964 3674
rect 364260 3602 364288 135526
rect 364616 3868 364668 3874
rect 364616 3810 364668 3816
rect 363512 3596 363564 3602
rect 363512 3538 363564 3544
rect 364248 3596 364300 3602
rect 364248 3538 364300 3544
rect 361120 2984 361172 2990
rect 361120 2926 361172 2932
rect 361132 480 361160 2926
rect 362316 2916 362368 2922
rect 362316 2858 362368 2864
rect 362328 480 362356 2858
rect 363524 480 363552 3538
rect 364628 480 364656 3810
rect 365640 2854 365668 135526
rect 365812 3528 365864 3534
rect 365812 3470 365864 3476
rect 365628 2848 365680 2854
rect 365628 2790 365680 2796
rect 365824 480 365852 3470
rect 366928 2990 366956 138366
rect 367848 135590 367876 138366
rect 368676 135590 368704 138366
rect 367008 135584 367060 135590
rect 367008 135526 367060 135532
rect 367836 135584 367888 135590
rect 367836 135526 367888 135532
rect 368388 135584 368440 135590
rect 368388 135526 368440 135532
rect 368664 135584 368716 135590
rect 368664 135526 368716 135532
rect 367020 3874 367048 135526
rect 368400 15910 368428 135526
rect 368388 15904 368440 15910
rect 368388 15846 368440 15852
rect 367008 3868 367060 3874
rect 367008 3810 367060 3816
rect 369688 3534 369716 138366
rect 370424 135590 370452 138366
rect 371344 135590 371372 138366
rect 369768 135584 369820 135590
rect 369768 135526 369820 135532
rect 370412 135584 370464 135590
rect 370412 135526 370464 135532
rect 371148 135584 371200 135590
rect 371148 135526 371200 135532
rect 371332 135584 371384 135590
rect 371332 135526 371384 135532
rect 372436 135584 372488 135590
rect 372436 135526 372488 135532
rect 369676 3528 369728 3534
rect 369676 3470 369728 3476
rect 369400 3324 369452 3330
rect 369400 3266 369452 3272
rect 368204 3120 368256 3126
rect 368204 3062 368256 3068
rect 367008 3052 367060 3058
rect 367008 2994 367060 3000
rect 366916 2984 366968 2990
rect 366916 2926 366968 2932
rect 367020 480 367048 2994
rect 368216 480 368244 3062
rect 369412 480 369440 3266
rect 369780 2922 369808 135526
rect 371160 4826 371188 135526
rect 371148 4820 371200 4826
rect 371148 4762 371200 4768
rect 371700 3256 371752 3262
rect 371700 3198 371752 3204
rect 370596 3188 370648 3194
rect 370596 3130 370648 3136
rect 369768 2916 369820 2922
rect 369768 2858 369820 2864
rect 370608 480 370636 3130
rect 371712 480 371740 3198
rect 372448 2990 372476 135526
rect 372540 3126 372568 138366
rect 373000 136066 373028 138366
rect 372988 136060 373040 136066
rect 372988 136002 373040 136008
rect 373920 3466 373948 138366
rect 374092 135924 374144 135930
rect 374092 135866 374144 135872
rect 372896 3460 372948 3466
rect 372896 3402 372948 3408
rect 373908 3460 373960 3466
rect 373908 3402 373960 3408
rect 372528 3120 372580 3126
rect 372528 3062 372580 3068
rect 372436 2984 372488 2990
rect 372436 2926 372488 2932
rect 372908 480 372936 3402
rect 374104 480 374132 135866
rect 374748 135590 374776 138366
rect 375576 135590 375604 138366
rect 374736 135584 374788 135590
rect 374736 135526 374788 135532
rect 375288 135584 375340 135590
rect 375288 135526 375340 135532
rect 375564 135584 375616 135590
rect 375564 135526 375616 135532
rect 376576 135584 376628 135590
rect 376576 135526 376628 135532
rect 375300 6914 375328 135526
rect 376588 11762 376616 135526
rect 376576 11756 376628 11762
rect 376576 11698 376628 11704
rect 375208 6886 375328 6914
rect 375208 3262 375236 6886
rect 375288 4140 375340 4146
rect 375288 4082 375340 4088
rect 375196 3256 375248 3262
rect 375196 3198 375248 3204
rect 375300 480 375328 4082
rect 376680 3398 376708 138366
rect 377324 135522 377352 138366
rect 378060 138366 378134 138394
rect 379026 138394 379054 138652
rect 379854 138394 379882 138652
rect 380774 138394 380802 138652
rect 381602 138394 381630 138652
rect 382430 138394 382458 138652
rect 383350 138394 383378 138652
rect 384178 138394 384206 138652
rect 385006 138394 385034 138652
rect 379026 138366 379468 138394
rect 379854 138366 379928 138394
rect 380774 138366 380848 138394
rect 381602 138366 381676 138394
rect 382430 138366 382504 138394
rect 383350 138366 383516 138394
rect 384178 138366 384252 138394
rect 378060 135930 378088 138366
rect 378048 135924 378100 135930
rect 378048 135866 378100 135872
rect 377312 135516 377364 135522
rect 377312 135458 377364 135464
rect 378048 135516 378100 135522
rect 378048 135458 378100 135464
rect 377680 4956 377732 4962
rect 377680 4898 377732 4904
rect 376484 3392 376536 3398
rect 376484 3334 376536 3340
rect 376668 3392 376720 3398
rect 376668 3334 376720 3340
rect 376496 480 376524 3334
rect 377692 480 377720 4898
rect 378060 3194 378088 135458
rect 379440 3806 379468 138366
rect 379900 135386 379928 138366
rect 380820 135522 380848 138366
rect 381648 135590 381676 138366
rect 382476 135590 382504 138366
rect 381636 135584 381688 135590
rect 381636 135526 381688 135532
rect 382188 135584 382240 135590
rect 382188 135526 382240 135532
rect 382464 135584 382516 135590
rect 382464 135526 382516 135532
rect 380808 135516 380860 135522
rect 380808 135458 380860 135464
rect 381544 135516 381596 135522
rect 381544 135458 381596 135464
rect 379888 135380 379940 135386
rect 379888 135322 379940 135328
rect 380808 135380 380860 135386
rect 380808 135322 380860 135328
rect 379980 4004 380032 4010
rect 379980 3946 380032 3952
rect 378876 3800 378928 3806
rect 378876 3742 378928 3748
rect 379428 3800 379480 3806
rect 379428 3742 379480 3748
rect 378048 3188 378100 3194
rect 378048 3130 378100 3136
rect 378888 480 378916 3742
rect 379992 480 380020 3946
rect 380820 3330 380848 135322
rect 381556 14482 381584 135458
rect 381544 14476 381596 14482
rect 381544 14418 381596 14424
rect 381176 7608 381228 7614
rect 381176 7550 381228 7556
rect 380808 3324 380860 3330
rect 380808 3266 380860 3272
rect 381188 480 381216 7550
rect 382200 4146 382228 135526
rect 383488 5234 383516 138366
rect 384224 135590 384252 138366
rect 384868 138366 385034 138394
rect 385926 138394 385954 138652
rect 386754 138394 386782 138652
rect 387582 138394 387610 138652
rect 388502 138394 388530 138652
rect 389330 138394 389358 138652
rect 390158 138394 390186 138652
rect 391078 138394 391106 138652
rect 391906 138394 391934 138652
rect 385926 138366 386000 138394
rect 386754 138366 386828 138394
rect 387582 138366 387748 138394
rect 388502 138366 388576 138394
rect 389330 138366 389404 138394
rect 390158 138366 390416 138394
rect 391078 138366 391152 138394
rect 383568 135584 383620 135590
rect 383568 135526 383620 135532
rect 384212 135584 384264 135590
rect 384212 135526 384264 135532
rect 383476 5228 383528 5234
rect 383476 5170 383528 5176
rect 382188 4140 382240 4146
rect 382188 4082 382240 4088
rect 383476 4072 383528 4078
rect 383476 4014 383528 4020
rect 382372 3664 382424 3670
rect 382372 3606 382424 3612
rect 382384 480 382412 3606
rect 383488 2122 383516 4014
rect 383580 4010 383608 135526
rect 384764 4888 384816 4894
rect 384764 4830 384816 4836
rect 383568 4004 383620 4010
rect 383568 3946 383620 3952
rect 383488 2094 383608 2122
rect 383580 480 383608 2094
rect 384776 480 384804 4830
rect 384868 3806 384896 138366
rect 385972 136134 386000 138366
rect 385960 136128 386012 136134
rect 385960 136070 386012 136076
rect 385684 135992 385736 135998
rect 385684 135934 385736 135940
rect 384948 135584 385000 135590
rect 384948 135526 385000 135532
rect 384960 3942 384988 135526
rect 385696 4214 385724 135934
rect 386800 135590 386828 138366
rect 386788 135584 386840 135590
rect 386788 135526 386840 135532
rect 387616 135584 387668 135590
rect 387616 135526 387668 135532
rect 385684 4208 385736 4214
rect 385684 4150 385736 4156
rect 384948 3936 385000 3942
rect 384948 3878 385000 3884
rect 387156 3868 387208 3874
rect 387156 3810 387208 3816
rect 384856 3800 384908 3806
rect 384856 3742 384908 3748
rect 385960 3732 386012 3738
rect 385960 3674 386012 3680
rect 385972 480 386000 3674
rect 387168 480 387196 3810
rect 387628 3670 387656 135526
rect 387720 3738 387748 138366
rect 388548 135590 388576 138366
rect 389376 135590 389404 138366
rect 388536 135584 388588 135590
rect 388536 135526 388588 135532
rect 389088 135584 389140 135590
rect 389088 135526 389140 135532
rect 389364 135584 389416 135590
rect 389364 135526 389416 135532
rect 388260 8968 388312 8974
rect 388260 8910 388312 8916
rect 387708 3732 387760 3738
rect 387708 3674 387760 3680
rect 387616 3664 387668 3670
rect 387616 3606 387668 3612
rect 388272 480 388300 8910
rect 389100 5166 389128 135526
rect 389088 5160 389140 5166
rect 389088 5102 389140 5108
rect 389456 3596 389508 3602
rect 389456 3538 389508 3544
rect 389468 480 389496 3538
rect 390388 3369 390416 138366
rect 391124 136202 391152 138366
rect 391860 138366 391934 138394
rect 392826 138394 392854 138652
rect 393654 138394 393682 138652
rect 394482 138394 394510 138652
rect 395402 138394 395430 138652
rect 396230 138394 396258 138652
rect 397058 138394 397086 138652
rect 397978 138394 398006 138652
rect 398806 138394 398834 138652
rect 392826 138366 393268 138394
rect 393654 138366 393728 138394
rect 394482 138366 394648 138394
rect 395402 138366 395476 138394
rect 396230 138366 396304 138394
rect 397058 138366 397316 138394
rect 397978 138366 398052 138394
rect 391112 136196 391164 136202
rect 391112 136138 391164 136144
rect 391860 135998 391888 138366
rect 391848 135992 391900 135998
rect 391848 135934 391900 135940
rect 390468 135584 390520 135590
rect 390468 135526 390520 135532
rect 390480 3874 390508 135526
rect 391848 4208 391900 4214
rect 391848 4150 391900 4156
rect 390468 3868 390520 3874
rect 390468 3810 390520 3816
rect 390374 3360 390430 3369
rect 390374 3295 390430 3304
rect 390652 2848 390704 2854
rect 390652 2790 390704 2796
rect 390664 480 390692 2790
rect 391860 480 391888 4150
rect 393240 3602 393268 138366
rect 393700 136474 393728 138366
rect 393688 136468 393740 136474
rect 393688 136410 393740 136416
rect 394620 5030 394648 138366
rect 395448 136406 395476 138366
rect 395436 136400 395488 136406
rect 395436 136342 395488 136348
rect 395344 136060 395396 136066
rect 395344 136002 395396 136008
rect 395252 15904 395304 15910
rect 395252 15846 395304 15852
rect 394608 5024 394660 5030
rect 394608 4966 394660 4972
rect 393044 3596 393096 3602
rect 393044 3538 393096 3544
rect 393228 3596 393280 3602
rect 393228 3538 393280 3544
rect 393056 480 393084 3538
rect 395264 3482 395292 15846
rect 395356 4214 395384 136002
rect 396276 135590 396304 138366
rect 396264 135584 396316 135590
rect 396264 135526 396316 135532
rect 397288 7682 397316 138366
rect 398024 135590 398052 138366
rect 398760 138366 398834 138394
rect 399634 138394 399662 138652
rect 400554 138394 400582 138652
rect 401382 138394 401410 138652
rect 402302 138394 402330 138652
rect 403130 138394 403158 138652
rect 403958 138394 403986 138652
rect 404878 138394 404906 138652
rect 405706 138394 405734 138652
rect 399634 138366 399708 138394
rect 400554 138366 400628 138394
rect 401382 138366 401548 138394
rect 402302 138366 402376 138394
rect 403130 138366 403204 138394
rect 403958 138366 404032 138394
rect 404878 138366 404952 138394
rect 398760 136542 398788 138366
rect 398748 136536 398800 136542
rect 398748 136478 398800 136484
rect 399484 136196 399536 136202
rect 399484 136138 399536 136144
rect 397368 135584 397420 135590
rect 397368 135526 397420 135532
rect 398012 135584 398064 135590
rect 398012 135526 398064 135532
rect 398748 135584 398800 135590
rect 398748 135526 398800 135532
rect 397276 7676 397328 7682
rect 397276 7618 397328 7624
rect 397380 5098 397408 135526
rect 397368 5092 397420 5098
rect 397368 5034 397420 5040
rect 395344 4208 395396 4214
rect 395344 4150 395396 4156
rect 398760 3534 398788 135526
rect 399496 5302 399524 136138
rect 399680 135862 399708 138366
rect 400600 136338 400628 138366
rect 400588 136332 400640 136338
rect 400588 136274 400640 136280
rect 400864 135924 400916 135930
rect 400864 135866 400916 135872
rect 399668 135856 399720 135862
rect 399668 135798 399720 135804
rect 399484 5296 399536 5302
rect 399484 5238 399536 5244
rect 400876 4826 400904 135866
rect 401520 4962 401548 138366
rect 402348 135930 402376 138366
rect 402336 135924 402388 135930
rect 402336 135866 402388 135872
rect 403176 135590 403204 138366
rect 404004 136610 404032 138366
rect 403992 136604 404044 136610
rect 403992 136546 404044 136552
rect 404924 135590 404952 138366
rect 405660 138366 405734 138394
rect 406534 138394 406562 138652
rect 407454 138394 407482 138652
rect 408282 138394 408310 138652
rect 409110 138394 409138 138652
rect 410030 138394 410058 138652
rect 410858 138394 410886 138652
rect 411778 138394 411806 138652
rect 412606 138394 412634 138652
rect 406534 138366 406608 138394
rect 407454 138366 407528 138394
rect 408282 138366 408448 138394
rect 409110 138366 409184 138394
rect 410030 138366 410104 138394
rect 410858 138366 411116 138394
rect 411778 138366 411852 138394
rect 403164 135584 403216 135590
rect 403164 135526 403216 135532
rect 404268 135584 404320 135590
rect 404268 135526 404320 135532
rect 404912 135584 404964 135590
rect 404912 135526 404964 135532
rect 401508 4956 401560 4962
rect 401508 4898 401560 4904
rect 398932 4820 398984 4826
rect 398932 4762 398984 4768
rect 400864 4820 400916 4826
rect 400864 4762 400916 4768
rect 397736 3528 397788 3534
rect 395264 3454 395384 3482
rect 397736 3470 397788 3476
rect 398748 3528 398800 3534
rect 398748 3470 398800 3476
rect 394240 3052 394292 3058
rect 394240 2994 394292 3000
rect 394252 480 394280 2994
rect 395356 480 395384 3454
rect 396540 2916 396592 2922
rect 396540 2858 396592 2864
rect 396552 480 396580 2858
rect 397748 480 397776 3470
rect 398944 480 398972 4762
rect 402520 4208 402572 4214
rect 402520 4150 402572 4156
rect 401324 3120 401376 3126
rect 401324 3062 401376 3068
rect 400128 2984 400180 2990
rect 400128 2926 400180 2932
rect 400140 480 400168 2926
rect 401336 480 401364 3062
rect 402532 480 402560 4150
rect 404280 3466 404308 135526
rect 403624 3460 403676 3466
rect 403624 3402 403676 3408
rect 404268 3460 404320 3466
rect 404268 3402 404320 3408
rect 403636 480 403664 3402
rect 404820 3256 404872 3262
rect 404820 3198 404872 3204
rect 404832 480 404860 3198
rect 405660 2990 405688 138366
rect 406580 135590 406608 138366
rect 407500 136202 407528 138366
rect 407488 136196 407540 136202
rect 407488 136138 407540 136144
rect 407764 136128 407816 136134
rect 407764 136070 407816 136076
rect 406384 135584 406436 135590
rect 406384 135526 406436 135532
rect 406568 135584 406620 135590
rect 406568 135526 406620 135532
rect 407028 135584 407080 135590
rect 407028 135526 407080 135532
rect 406396 11762 406424 135526
rect 406016 11756 406068 11762
rect 406016 11698 406068 11704
rect 406384 11756 406436 11762
rect 406384 11698 406436 11704
rect 405648 2984 405700 2990
rect 405648 2926 405700 2932
rect 406028 480 406056 11698
rect 407040 4894 407068 135526
rect 407776 5370 407804 136070
rect 408420 6914 408448 138366
rect 409156 136202 409184 138366
rect 409144 136196 409196 136202
rect 409144 136138 409196 136144
rect 410076 135318 410104 138366
rect 410064 135312 410116 135318
rect 410064 135254 410116 135260
rect 408328 6886 408448 6914
rect 407764 5364 407816 5370
rect 407764 5306 407816 5312
rect 407028 4888 407080 4894
rect 407028 4830 407080 4836
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 407224 480 407252 3334
rect 408328 2854 408356 6886
rect 409604 4820 409656 4826
rect 409604 4762 409656 4768
rect 408408 3188 408460 3194
rect 408408 3130 408460 3136
rect 408316 2848 408368 2854
rect 408316 2790 408368 2796
rect 408420 480 408448 3130
rect 409616 480 409644 4762
rect 410800 4140 410852 4146
rect 410800 4082 410852 4088
rect 410812 480 410840 4082
rect 411088 3126 411116 138366
rect 411824 135318 411852 138366
rect 412560 138366 412634 138394
rect 413434 138394 413462 138652
rect 414354 138394 414382 138652
rect 415182 138394 415210 138652
rect 416010 138394 416038 138652
rect 416930 138394 416958 138652
rect 417758 138394 417786 138652
rect 418586 138394 418614 138652
rect 419506 138394 419534 138652
rect 413434 138366 413508 138394
rect 414354 138366 414428 138394
rect 415182 138366 415348 138394
rect 416010 138366 416084 138394
rect 416930 138366 417004 138394
rect 417758 138366 418108 138394
rect 418586 138366 418660 138394
rect 411168 135312 411220 135318
rect 411168 135254 411220 135260
rect 411812 135312 411864 135318
rect 411812 135254 411864 135260
rect 412456 135312 412508 135318
rect 412456 135254 412508 135260
rect 411076 3120 411128 3126
rect 411076 3062 411128 3068
rect 411180 2922 411208 135254
rect 412468 4826 412496 135254
rect 412456 4820 412508 4826
rect 412456 4762 412508 4768
rect 411904 3324 411956 3330
rect 411904 3266 411956 3272
rect 411168 2916 411220 2922
rect 411168 2858 411220 2864
rect 411916 480 411944 3266
rect 412560 3194 412588 138366
rect 413480 135318 413508 138366
rect 414400 136066 414428 138366
rect 414388 136060 414440 136066
rect 414388 136002 414440 136008
rect 414664 135992 414716 135998
rect 414664 135934 414716 135940
rect 413468 135312 413520 135318
rect 413468 135254 413520 135260
rect 413928 135312 413980 135318
rect 413928 135254 413980 135260
rect 412640 14476 412692 14482
rect 412640 14418 412692 14424
rect 412548 3188 412600 3194
rect 412548 3130 412600 3136
rect 412652 490 412680 14418
rect 413940 3058 413968 135254
rect 414676 5438 414704 135934
rect 414664 5432 414716 5438
rect 414664 5374 414716 5380
rect 414296 4004 414348 4010
rect 414296 3946 414348 3952
rect 413928 3052 413980 3058
rect 413928 2994 413980 3000
rect 412928 598 413140 626
rect 412928 490 412956 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 462 412956 490
rect 413112 480 413140 598
rect 414308 480 414336 3946
rect 415320 3330 415348 138366
rect 416056 135318 416084 138366
rect 416976 135998 417004 138366
rect 416964 135992 417016 135998
rect 416964 135934 417016 135940
rect 417424 135856 417476 135862
rect 417424 135798 417476 135804
rect 416044 135312 416096 135318
rect 416044 135254 416096 135260
rect 416688 135312 416740 135318
rect 416688 135254 416740 135260
rect 416700 6914 416728 135254
rect 416608 6886 416728 6914
rect 415492 4072 415544 4078
rect 415492 4014 415544 4020
rect 415308 3324 415360 3330
rect 415308 3266 415360 3272
rect 415504 480 415532 4014
rect 416608 3262 416636 6886
rect 417436 5234 417464 135798
rect 416688 5228 416740 5234
rect 416688 5170 416740 5176
rect 417424 5228 417476 5234
rect 417424 5170 417476 5176
rect 416596 3256 416648 3262
rect 416596 3198 416648 3204
rect 416700 480 416728 5170
rect 418080 4010 418108 138366
rect 418632 135590 418660 138366
rect 419368 138366 419534 138394
rect 420334 138394 420362 138652
rect 421162 138394 421190 138652
rect 422082 138394 422110 138652
rect 422910 138394 422938 138652
rect 423830 138394 423858 138652
rect 424658 138394 424686 138652
rect 425486 138394 425514 138652
rect 426406 138394 426434 138652
rect 420334 138366 420408 138394
rect 421162 138366 421236 138394
rect 422082 138366 422156 138394
rect 422910 138366 422984 138394
rect 423830 138366 423904 138394
rect 424658 138366 424732 138394
rect 425486 138366 425560 138394
rect 418620 135584 418672 135590
rect 418620 135526 418672 135532
rect 419368 7614 419396 138366
rect 420380 135590 420408 138366
rect 421208 135590 421236 138366
rect 422128 135998 422156 138366
rect 422116 135992 422168 135998
rect 422116 135934 422168 135940
rect 421564 135924 421616 135930
rect 421564 135866 421616 135872
rect 419448 135584 419500 135590
rect 419448 135526 419500 135532
rect 420368 135584 420420 135590
rect 420368 135526 420420 135532
rect 420828 135584 420880 135590
rect 420828 135526 420880 135532
rect 421196 135584 421248 135590
rect 421196 135526 421248 135532
rect 419356 7608 419408 7614
rect 419356 7550 419408 7556
rect 419460 4146 419488 135526
rect 420184 5364 420236 5370
rect 420184 5306 420236 5312
rect 419448 4140 419500 4146
rect 419448 4082 419500 4088
rect 418068 4004 418120 4010
rect 418068 3946 418120 3952
rect 417884 3936 417936 3942
rect 417884 3878 417936 3884
rect 417896 480 417924 3878
rect 418988 3800 419040 3806
rect 418988 3742 419040 3748
rect 419000 480 419028 3742
rect 420196 480 420224 5306
rect 420840 4078 420868 135526
rect 421576 5370 421604 135866
rect 422956 135590 422984 138366
rect 423876 135590 423904 138366
rect 424704 135862 424732 138366
rect 424692 135856 424744 135862
rect 424692 135798 424744 135804
rect 422208 135584 422260 135590
rect 422208 135526 422260 135532
rect 422944 135584 422996 135590
rect 422944 135526 422996 135532
rect 423588 135584 423640 135590
rect 423588 135526 423640 135532
rect 423864 135584 423916 135590
rect 423864 135526 423916 135532
rect 424968 135584 425020 135590
rect 424968 135526 425020 135532
rect 421564 5364 421616 5370
rect 421564 5306 421616 5312
rect 420828 4072 420880 4078
rect 420828 4014 420880 4020
rect 421380 3732 421432 3738
rect 421380 3674 421432 3680
rect 421392 480 421420 3674
rect 422220 3398 422248 135526
rect 423600 3806 423628 135526
rect 424980 6914 425008 135526
rect 425532 135522 425560 138366
rect 426268 138366 426434 138394
rect 427234 138394 427262 138652
rect 428062 138394 428090 138652
rect 428982 138394 429010 138652
rect 429810 138394 429838 138652
rect 430638 138394 430666 138652
rect 431558 138394 431586 138652
rect 432386 138394 432414 138652
rect 433306 138394 433334 138652
rect 427234 138366 427308 138394
rect 428062 138366 428136 138394
rect 428982 138366 429056 138394
rect 429810 138366 429884 138394
rect 430638 138366 430712 138394
rect 431558 138366 431908 138394
rect 432386 138366 432460 138394
rect 425520 135516 425572 135522
rect 425520 135458 425572 135464
rect 424888 6886 425008 6914
rect 423772 5160 423824 5166
rect 423772 5102 423824 5108
rect 423588 3800 423640 3806
rect 423588 3742 423640 3748
rect 422576 3664 422628 3670
rect 422576 3606 422628 3612
rect 422208 3392 422260 3398
rect 422208 3334 422260 3340
rect 422588 480 422616 3606
rect 423784 480 423812 5102
rect 424888 3942 424916 6886
rect 424876 3936 424928 3942
rect 424876 3878 424928 3884
rect 424968 3868 425020 3874
rect 424968 3810 425020 3816
rect 424980 480 425008 3810
rect 426268 3670 426296 138366
rect 427280 135726 427308 138366
rect 427268 135720 427320 135726
rect 427268 135662 427320 135668
rect 428108 135590 428136 138366
rect 428096 135584 428148 135590
rect 428096 135526 428148 135532
rect 426348 135516 426400 135522
rect 426348 135458 426400 135464
rect 426360 3874 426388 135458
rect 428464 5432 428516 5438
rect 428464 5374 428516 5380
rect 427268 5296 427320 5302
rect 427268 5238 427320 5244
rect 426348 3868 426400 3874
rect 426348 3810 426400 3816
rect 426256 3664 426308 3670
rect 426256 3606 426308 3612
rect 426162 3360 426218 3369
rect 426162 3295 426218 3304
rect 426176 480 426204 3295
rect 427280 480 427308 5238
rect 428476 480 428504 5374
rect 429028 3777 429056 138366
rect 429752 136536 429804 136542
rect 429752 136478 429804 136484
rect 429108 135584 429160 135590
rect 429108 135526 429160 135532
rect 429014 3768 429070 3777
rect 429120 3738 429148 135526
rect 429764 132494 429792 136478
rect 429856 135658 429884 138366
rect 429936 136468 429988 136474
rect 429936 136410 429988 136416
rect 429844 135652 429896 135658
rect 429844 135594 429896 135600
rect 429764 132466 429884 132494
rect 429856 5166 429884 132466
rect 429844 5160 429896 5166
rect 429844 5102 429896 5108
rect 429948 4214 429976 136410
rect 430684 135590 430712 138366
rect 430672 135584 430724 135590
rect 430672 135526 430724 135532
rect 431776 135584 431828 135590
rect 431776 135526 431828 135532
rect 431788 6662 431816 135526
rect 431776 6656 431828 6662
rect 431776 6598 431828 6604
rect 429936 4208 429988 4214
rect 429936 4150 429988 4156
rect 430856 4208 430908 4214
rect 430856 4150 430908 4156
rect 429014 3703 429070 3712
rect 429108 3732 429160 3738
rect 429108 3674 429160 3680
rect 429660 3596 429712 3602
rect 429660 3538 429712 3544
rect 429672 480 429700 3538
rect 430868 480 430896 4150
rect 431880 3602 431908 138366
rect 431960 135856 432012 135862
rect 431960 135798 432012 135804
rect 431972 4214 432000 135798
rect 432432 135794 432460 138366
rect 433260 138366 433334 138394
rect 434134 138394 434162 138652
rect 434962 138394 434990 138652
rect 435882 138394 435910 138652
rect 436710 138394 436738 138652
rect 437538 138394 437566 138652
rect 438458 138394 438486 138652
rect 439286 138394 439314 138652
rect 440114 138394 440142 138652
rect 434134 138366 434208 138394
rect 434962 138366 435036 138394
rect 435882 138366 436048 138394
rect 436710 138366 436784 138394
rect 437538 138366 437612 138394
rect 438458 138366 438532 138394
rect 439286 138366 439360 138394
rect 432420 135788 432472 135794
rect 432420 135730 432472 135736
rect 433260 6594 433288 138366
rect 434180 135590 434208 138366
rect 435008 135862 435036 138366
rect 435364 136604 435416 136610
rect 435364 136546 435416 136552
rect 434996 135856 435048 135862
rect 434996 135798 435048 135804
rect 434168 135584 434220 135590
rect 434168 135526 434220 135532
rect 434628 135584 434680 135590
rect 434628 135526 434680 135532
rect 433248 6588 433300 6594
rect 433248 6530 433300 6536
rect 432052 5092 432104 5098
rect 432052 5034 432104 5040
rect 431960 4208 432012 4214
rect 431960 4150 432012 4156
rect 431868 3596 431920 3602
rect 431868 3538 431920 3544
rect 432064 480 432092 5034
rect 434444 4752 434496 4758
rect 434444 4694 434496 4700
rect 433248 4208 433300 4214
rect 433248 4150 433300 4156
rect 433260 480 433288 4150
rect 434456 480 434484 4694
rect 434640 3641 434668 135526
rect 435376 5030 435404 136546
rect 436020 15910 436048 138366
rect 436652 135720 436704 135726
rect 436652 135662 436704 135668
rect 436664 132494 436692 135662
rect 436756 135590 436784 138366
rect 437584 135590 437612 138366
rect 438504 135726 438532 138366
rect 438492 135720 438544 135726
rect 438492 135662 438544 135668
rect 439332 135590 439360 138366
rect 440068 138366 440142 138394
rect 441034 138394 441062 138652
rect 441862 138394 441890 138652
rect 442782 138394 442810 138652
rect 443610 138394 443638 138652
rect 441034 138366 441108 138394
rect 441862 138366 441936 138394
rect 442782 138366 442856 138394
rect 436744 135584 436796 135590
rect 436744 135526 436796 135532
rect 437388 135584 437440 135590
rect 437388 135526 437440 135532
rect 437572 135584 437624 135590
rect 437572 135526 437624 135532
rect 438768 135584 438820 135590
rect 438768 135526 438820 135532
rect 439320 135584 439372 135590
rect 439320 135526 439372 135532
rect 436664 132466 436784 132494
rect 436008 15904 436060 15910
rect 436008 15846 436060 15852
rect 435548 7676 435600 7682
rect 435548 7618 435600 7624
rect 435364 5024 435416 5030
rect 435364 4966 435416 4972
rect 434626 3632 434682 3641
rect 434626 3567 434682 3576
rect 435560 480 435588 7618
rect 436756 6186 436784 132466
rect 436744 6180 436796 6186
rect 436744 6122 436796 6128
rect 437400 3534 437428 135526
rect 438780 5506 438808 135526
rect 438768 5500 438820 5506
rect 438768 5442 438820 5448
rect 440068 5438 440096 138366
rect 441080 136542 441108 138366
rect 441068 136536 441120 136542
rect 441068 136478 441120 136484
rect 440240 136332 440292 136338
rect 440240 136274 440292 136280
rect 440148 135584 440200 135590
rect 440148 135526 440200 135532
rect 440056 5432 440108 5438
rect 440056 5374 440108 5380
rect 439136 5228 439188 5234
rect 439136 5170 439188 5176
rect 437940 5160 437992 5166
rect 437940 5102 437992 5108
rect 436744 3528 436796 3534
rect 436744 3470 436796 3476
rect 437388 3528 437440 3534
rect 437388 3470 437440 3476
rect 436756 480 436784 3470
rect 437952 480 437980 5102
rect 439148 480 439176 5170
rect 440160 3505 440188 135526
rect 440252 16574 440280 136274
rect 441908 135590 441936 138366
rect 441896 135584 441948 135590
rect 441896 135526 441948 135532
rect 440252 16546 440372 16574
rect 440146 3496 440202 3505
rect 440146 3431 440202 3440
rect 440344 480 440372 16546
rect 442632 5364 442684 5370
rect 442632 5306 442684 5312
rect 441528 4956 441580 4962
rect 441528 4898 441580 4904
rect 441540 480 441568 4898
rect 442644 480 442672 5306
rect 442828 5302 442856 138366
rect 443564 138366 443638 138394
rect 444438 138394 444466 138652
rect 445358 138394 445386 138652
rect 446186 138394 446214 138652
rect 447014 138394 447042 138652
rect 447934 138394 447962 138652
rect 448762 138394 448790 138652
rect 449590 138394 449618 138652
rect 450510 138394 450538 138652
rect 451338 138394 451366 138652
rect 452166 138394 452194 138652
rect 453086 138394 453114 138652
rect 453914 138394 453942 138652
rect 454834 138394 454862 138652
rect 455662 138394 455690 138652
rect 456490 138394 456518 138652
rect 457410 138394 457438 138652
rect 458238 138394 458266 138652
rect 459066 138394 459094 138652
rect 459986 138394 460014 138652
rect 460814 138394 460842 138652
rect 444438 138366 444512 138394
rect 445358 138366 445708 138394
rect 446186 138366 446260 138394
rect 447014 138366 447088 138394
rect 447934 138366 448008 138394
rect 448762 138366 448836 138394
rect 449590 138366 449664 138394
rect 450510 138366 450584 138394
rect 451338 138366 451412 138394
rect 452166 138366 452608 138394
rect 453086 138366 453160 138394
rect 453914 138366 453988 138394
rect 454834 138366 454908 138394
rect 455662 138366 455736 138394
rect 456490 138366 456564 138394
rect 457410 138366 457484 138394
rect 458238 138366 458312 138394
rect 459066 138366 459140 138394
rect 459986 138366 460060 138394
rect 442908 135584 442960 135590
rect 442908 135526 442960 135532
rect 442816 5296 442868 5302
rect 442816 5238 442868 5244
rect 442920 3369 442948 135526
rect 443564 135522 443592 138366
rect 443644 136536 443696 136542
rect 443644 136478 443696 136484
rect 443552 135516 443604 135522
rect 443552 135458 443604 135464
rect 443656 6458 443684 136478
rect 444484 136406 444512 138366
rect 444472 136400 444524 136406
rect 444472 136342 444524 136348
rect 443644 6452 443696 6458
rect 443644 6394 443696 6400
rect 445680 5370 445708 138366
rect 446232 135590 446260 138366
rect 446220 135584 446272 135590
rect 446220 135526 446272 135532
rect 446956 135584 447008 135590
rect 446956 135526 447008 135532
rect 446968 47598 446996 135526
rect 446956 47592 447008 47598
rect 446956 47534 447008 47540
rect 445760 11756 445812 11762
rect 445760 11698 445812 11704
rect 445668 5364 445720 5370
rect 445668 5306 445720 5312
rect 445024 5024 445076 5030
rect 445024 4966 445076 4972
rect 443828 3460 443880 3466
rect 443828 3402 443880 3408
rect 442906 3360 442962 3369
rect 442906 3295 442962 3304
rect 443840 480 443868 3402
rect 445036 480 445064 4966
rect 445772 490 445800 11698
rect 447060 3466 447088 138366
rect 447980 135590 448008 138366
rect 448520 136264 448572 136270
rect 448520 136206 448572 136212
rect 447968 135584 448020 135590
rect 447968 135526 448020 135532
rect 448428 135584 448480 135590
rect 448428 135526 448480 135532
rect 448440 5234 448468 135526
rect 448428 5228 448480 5234
rect 448428 5170 448480 5176
rect 447048 3460 447100 3466
rect 447048 3402 447100 3408
rect 447416 2984 447468 2990
rect 447416 2926 447468 2932
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 2926
rect 448532 2378 448560 136206
rect 448808 135590 448836 138366
rect 449636 136542 449664 138366
rect 449624 136536 449676 136542
rect 449624 136478 449676 136484
rect 450452 136196 450504 136202
rect 450452 136138 450504 136144
rect 448796 135584 448848 135590
rect 448796 135526 448848 135532
rect 449808 135584 449860 135590
rect 449808 135526 449860 135532
rect 449820 11762 449848 135526
rect 450464 132494 450492 136138
rect 450556 135522 450584 138366
rect 451384 136338 451412 138366
rect 451372 136332 451424 136338
rect 451372 136274 451424 136280
rect 450544 135516 450596 135522
rect 450544 135458 450596 135464
rect 451188 135516 451240 135522
rect 451188 135458 451240 135464
rect 450464 132466 450584 132494
rect 449808 11756 449860 11762
rect 449808 11698 449860 11704
rect 448612 4888 448664 4894
rect 448612 4830 448664 4836
rect 448520 2372 448572 2378
rect 448520 2314 448572 2320
rect 448624 480 448652 4830
rect 450556 4418 450584 132466
rect 451200 5166 451228 135458
rect 451188 5160 451240 5166
rect 451188 5102 451240 5108
rect 450544 4412 450596 4418
rect 450544 4354 450596 4360
rect 452108 4412 452160 4418
rect 452108 4354 452160 4360
rect 450912 2848 450964 2854
rect 450912 2790 450964 2796
rect 449808 2372 449860 2378
rect 449808 2314 449860 2320
rect 449820 480 449848 2314
rect 450924 480 450952 2790
rect 452120 480 452148 4354
rect 452580 2854 452608 138366
rect 453132 135658 453160 138366
rect 453960 136474 453988 138366
rect 453948 136468 454000 136474
rect 453948 136410 454000 136416
rect 454880 135658 454908 138366
rect 455708 135658 455736 138366
rect 456536 136202 456564 138366
rect 457456 136270 457484 138366
rect 457444 136264 457496 136270
rect 457444 136206 457496 136212
rect 456524 136196 456576 136202
rect 456524 136138 456576 136144
rect 457536 136060 457588 136066
rect 457536 136002 457588 136008
rect 453120 135652 453172 135658
rect 453120 135594 453172 135600
rect 453948 135652 454000 135658
rect 453948 135594 454000 135600
rect 454868 135652 454920 135658
rect 454868 135594 454920 135600
rect 455328 135652 455380 135658
rect 455328 135594 455380 135600
rect 455696 135652 455748 135658
rect 455696 135594 455748 135600
rect 456708 135652 456760 135658
rect 456708 135594 456760 135600
rect 453960 5098 453988 135594
rect 453948 5092 454000 5098
rect 453948 5034 454000 5040
rect 454500 3120 454552 3126
rect 454500 3062 454552 3068
rect 453304 2916 453356 2922
rect 453304 2858 453356 2864
rect 452568 2848 452620 2854
rect 452568 2790 452620 2796
rect 453316 480 453344 2858
rect 454512 480 454540 3062
rect 455340 2922 455368 135594
rect 456720 5030 456748 135594
rect 457444 135516 457496 135522
rect 457444 135458 457496 135464
rect 456708 5024 456760 5030
rect 456708 4966 456760 4972
rect 455696 4820 455748 4826
rect 455696 4762 455748 4768
rect 455328 2916 455380 2922
rect 455328 2858 455380 2864
rect 455708 480 455736 4762
rect 457456 4690 457484 135458
rect 457444 4684 457496 4690
rect 457444 4626 457496 4632
rect 457548 4214 457576 136002
rect 458284 135318 458312 138366
rect 458272 135312 458324 135318
rect 458272 135254 458324 135260
rect 459112 134978 459140 138366
rect 460032 135318 460060 138366
rect 460768 138366 460842 138394
rect 461642 138394 461670 138652
rect 462562 138394 462590 138652
rect 463390 138394 463418 138652
rect 464310 138394 464338 138652
rect 465138 138394 465166 138652
rect 465966 138394 465994 138652
rect 466886 138394 466914 138652
rect 467714 138394 467742 138652
rect 468542 138394 468570 138652
rect 469462 138394 469490 138652
rect 470290 138394 470318 138652
rect 471118 138394 471146 138652
rect 472038 138394 472066 138652
rect 472866 138394 472894 138652
rect 473786 138394 473814 138652
rect 474614 138394 474642 138652
rect 475442 138394 475470 138652
rect 476362 138394 476390 138652
rect 477190 138394 477218 138652
rect 478018 138394 478046 138652
rect 478938 138394 478966 138652
rect 479766 138394 479794 138652
rect 480594 138394 480622 138652
rect 481514 138394 481542 138652
rect 461642 138366 461716 138394
rect 462562 138366 462636 138394
rect 463390 138366 463648 138394
rect 464310 138366 464384 138394
rect 465138 138366 465212 138394
rect 465966 138366 466040 138394
rect 466886 138366 466960 138394
rect 467714 138366 467788 138394
rect 468542 138366 468616 138394
rect 469462 138366 469536 138394
rect 470290 138366 470548 138394
rect 471118 138366 471192 138394
rect 472038 138366 472112 138394
rect 472866 138366 472940 138394
rect 473786 138366 473860 138394
rect 474614 138366 474688 138394
rect 475442 138366 475516 138394
rect 476362 138366 476436 138394
rect 477190 138366 477264 138394
rect 478018 138366 478092 138394
rect 478938 138366 479012 138394
rect 479766 138366 480116 138394
rect 480594 138366 480668 138394
rect 459376 135312 459428 135318
rect 459376 135254 459428 135260
rect 460020 135312 460072 135318
rect 460020 135254 460072 135260
rect 459100 134972 459152 134978
rect 459100 134914 459152 134920
rect 459388 4962 459416 135254
rect 459376 4956 459428 4962
rect 459376 4898 459428 4904
rect 460768 4826 460796 138366
rect 461584 135992 461636 135998
rect 461584 135934 461636 135940
rect 460848 135312 460900 135318
rect 460848 135254 460900 135260
rect 460756 4820 460808 4826
rect 460756 4762 460808 4768
rect 457536 4208 457588 4214
rect 457536 4150 457588 4156
rect 459192 4208 459244 4214
rect 459192 4150 459244 4156
rect 456892 3188 456944 3194
rect 456892 3130 456944 3136
rect 456904 480 456932 3130
rect 458088 3052 458140 3058
rect 458088 2994 458140 3000
rect 458100 480 458128 2994
rect 459204 480 459232 4150
rect 460388 3324 460440 3330
rect 460388 3266 460440 3272
rect 460400 480 460428 3266
rect 460860 2990 460888 135254
rect 461596 4214 461624 135934
rect 461688 135318 461716 138366
rect 462608 136066 462636 138366
rect 462596 136060 462648 136066
rect 462596 136002 462648 136008
rect 461676 135312 461728 135318
rect 461676 135254 461728 135260
rect 462228 135312 462280 135318
rect 462228 135254 462280 135260
rect 462240 6390 462268 135254
rect 462228 6384 462280 6390
rect 462228 6326 462280 6332
rect 463620 4894 463648 138366
rect 464252 136196 464304 136202
rect 464252 136138 464304 136144
rect 464264 128354 464292 136138
rect 464356 135318 464384 138366
rect 465184 135318 465212 138366
rect 466012 135522 466040 138366
rect 466932 135658 466960 138366
rect 467760 135998 467788 138366
rect 468484 136128 468536 136134
rect 468484 136070 468536 136076
rect 467748 135992 467800 135998
rect 467748 135934 467800 135940
rect 466920 135652 466972 135658
rect 466920 135594 466972 135600
rect 467748 135652 467800 135658
rect 467748 135594 467800 135600
rect 466000 135516 466052 135522
rect 466000 135458 466052 135464
rect 464344 135312 464396 135318
rect 464344 135254 464396 135260
rect 464988 135312 465040 135318
rect 464988 135254 465040 135260
rect 465172 135312 465224 135318
rect 465172 135254 465224 135260
rect 466368 135312 466420 135318
rect 466368 135254 466420 135260
rect 464264 128326 464384 128354
rect 464356 6526 464384 128326
rect 464344 6520 464396 6526
rect 464344 6462 464396 6468
rect 465000 6322 465028 135254
rect 466276 7608 466328 7614
rect 466276 7550 466328 7556
rect 464988 6316 465040 6322
rect 464988 6258 465040 6264
rect 463608 4888 463660 4894
rect 463608 4830 463660 4836
rect 461584 4208 461636 4214
rect 461584 4150 461636 4156
rect 462780 4208 462832 4214
rect 462780 4150 462832 4156
rect 461584 3256 461636 3262
rect 461584 3198 461636 3204
rect 460848 2984 460900 2990
rect 460848 2926 460900 2932
rect 461596 480 461624 3198
rect 462792 480 462820 4150
rect 465172 4140 465224 4146
rect 465172 4082 465224 4088
rect 463976 4004 464028 4010
rect 463976 3946 464028 3952
rect 463988 480 464016 3946
rect 465184 480 465212 4082
rect 466288 480 466316 7550
rect 466380 3058 466408 135254
rect 467760 6254 467788 135594
rect 467748 6248 467800 6254
rect 467748 6190 467800 6196
rect 468496 4214 468524 136070
rect 468588 135658 468616 138366
rect 469508 136202 469536 138366
rect 469496 136196 469548 136202
rect 469496 136138 469548 136144
rect 468576 135652 468628 135658
rect 468576 135594 468628 135600
rect 469128 135652 469180 135658
rect 469128 135594 469180 135600
rect 469140 8974 469168 135594
rect 469128 8968 469180 8974
rect 469128 8910 469180 8916
rect 468484 4208 468536 4214
rect 468484 4150 468536 4156
rect 469864 4208 469916 4214
rect 469864 4150 469916 4156
rect 467472 4072 467524 4078
rect 467472 4014 467524 4020
rect 466368 3052 466420 3058
rect 466368 2994 466420 3000
rect 467484 480 467512 4014
rect 468668 3392 468720 3398
rect 468668 3334 468720 3340
rect 468680 480 468708 3334
rect 469876 480 469904 4150
rect 470520 3126 470548 138366
rect 471164 135590 471192 138366
rect 471244 135924 471296 135930
rect 471244 135866 471296 135872
rect 471152 135584 471204 135590
rect 471152 135526 471204 135532
rect 471256 4214 471284 135866
rect 472084 135590 472112 138366
rect 472912 135930 472940 138366
rect 472900 135924 472952 135930
rect 472900 135866 472952 135872
rect 471888 135584 471940 135590
rect 471888 135526 471940 135532
rect 472072 135584 472124 135590
rect 472072 135526 472124 135532
rect 473268 135584 473320 135590
rect 473268 135526 473320 135532
rect 471900 14482 471928 135526
rect 473280 49026 473308 135526
rect 473832 135522 473860 138366
rect 474660 136134 474688 138366
rect 474648 136128 474700 136134
rect 474648 136070 474700 136076
rect 475488 135590 475516 138366
rect 475476 135584 475528 135590
rect 475476 135526 475528 135532
rect 476028 135584 476080 135590
rect 476028 135526 476080 135532
rect 473820 135516 473872 135522
rect 473820 135458 473872 135464
rect 475384 135448 475436 135454
rect 475384 135390 475436 135396
rect 473268 49020 473320 49026
rect 473268 48962 473320 48968
rect 471888 14476 471940 14482
rect 471888 14418 471940 14424
rect 475396 4758 475424 135390
rect 475384 4752 475436 4758
rect 475384 4694 475436 4700
rect 471244 4208 471296 4214
rect 471244 4150 471296 4156
rect 473452 4208 473504 4214
rect 473452 4150 473504 4156
rect 472256 3936 472308 3942
rect 472256 3878 472308 3884
rect 471060 3800 471112 3806
rect 471060 3742 471112 3748
rect 470508 3120 470560 3126
rect 470508 3062 470560 3068
rect 471072 480 471100 3742
rect 472268 480 472296 3878
rect 473464 480 473492 4150
rect 474556 3868 474608 3874
rect 474556 3810 474608 3816
rect 474568 480 474596 3810
rect 475752 3664 475804 3670
rect 475752 3606 475804 3612
rect 475764 480 475792 3606
rect 476040 3194 476068 135526
rect 476408 135522 476436 138366
rect 476396 135516 476448 135522
rect 476396 135458 476448 135464
rect 477236 134842 477264 138366
rect 478064 135590 478092 138366
rect 478052 135584 478104 135590
rect 478052 135526 478104 135532
rect 478788 135584 478840 135590
rect 478788 135526 478840 135532
rect 477224 134836 477276 134842
rect 477224 134778 477276 134784
rect 476948 6180 477000 6186
rect 476948 6122 477000 6128
rect 476028 3188 476080 3194
rect 476028 3130 476080 3136
rect 476960 480 476988 6122
rect 478144 3732 478196 3738
rect 478144 3674 478196 3680
rect 478156 480 478184 3674
rect 478800 3262 478828 135526
rect 478984 134774 479012 138366
rect 478972 134768 479024 134774
rect 478972 134710 479024 134716
rect 480088 6186 480116 138366
rect 480640 135726 480668 138366
rect 481468 138366 481542 138394
rect 482342 138394 482370 138652
rect 483170 138394 483198 138652
rect 484090 138394 484118 138652
rect 484918 138394 484946 138652
rect 485838 138394 485866 138652
rect 486666 138394 486694 138652
rect 487494 138394 487522 138652
rect 488414 138394 488442 138652
rect 482342 138366 482416 138394
rect 483170 138366 483244 138394
rect 484090 138366 484164 138394
rect 484918 138366 484992 138394
rect 485838 138366 485912 138394
rect 486666 138366 486740 138394
rect 487494 138366 487568 138394
rect 480628 135720 480680 135726
rect 480628 135662 480680 135668
rect 481468 135318 481496 138366
rect 482388 136202 482416 138366
rect 482376 136196 482428 136202
rect 482376 136138 482428 136144
rect 483216 135726 483244 138366
rect 481548 135720 481600 135726
rect 481548 135662 481600 135668
rect 483204 135720 483256 135726
rect 483204 135662 483256 135668
rect 481456 135312 481508 135318
rect 481456 135254 481508 135260
rect 480076 6180 480128 6186
rect 480076 6122 480128 6128
rect 480536 4684 480588 4690
rect 480536 4626 480588 4632
rect 479338 3768 479394 3777
rect 479338 3703 479394 3712
rect 478788 3256 478840 3262
rect 478788 3198 478840 3204
rect 479352 480 479380 3703
rect 480548 480 480576 4626
rect 481560 3330 481588 135662
rect 482284 135380 482336 135386
rect 482284 135322 482336 135328
rect 481732 6656 481784 6662
rect 481732 6598 481784 6604
rect 481548 3324 481600 3330
rect 481548 3266 481600 3272
rect 481744 480 481772 6598
rect 482296 4214 482324 135322
rect 484136 134706 484164 138366
rect 484216 135720 484268 135726
rect 484216 135662 484268 135668
rect 484124 134700 484176 134706
rect 484124 134642 484176 134648
rect 482284 4208 482336 4214
rect 482284 4150 482336 4156
rect 484032 4208 484084 4214
rect 484032 4150 484084 4156
rect 482836 3596 482888 3602
rect 482836 3538 482888 3544
rect 482848 480 482876 3538
rect 484044 480 484072 4150
rect 484228 3398 484256 135662
rect 484964 133210 484992 138366
rect 485884 135726 485912 138366
rect 486424 135856 486476 135862
rect 486424 135798 486476 135804
rect 485872 135720 485924 135726
rect 485872 135662 485924 135668
rect 485044 135448 485096 135454
rect 485044 135390 485096 135396
rect 484952 133204 485004 133210
rect 484952 133146 485004 133152
rect 485056 4214 485084 135390
rect 485228 6588 485280 6594
rect 485228 6530 485280 6536
rect 485044 4208 485096 4214
rect 485044 4150 485096 4156
rect 484216 3392 484268 3398
rect 484216 3334 484268 3340
rect 485240 480 485268 6530
rect 486436 4690 486464 135798
rect 486712 135794 486740 138366
rect 486700 135788 486752 135794
rect 486700 135730 486752 135736
rect 487068 135720 487120 135726
rect 487068 135662 487120 135668
rect 486424 4684 486476 4690
rect 486424 4626 486476 4632
rect 487080 4146 487108 135662
rect 487540 135046 487568 138366
rect 488368 138366 488442 138394
rect 489242 138394 489270 138652
rect 490070 138394 490098 138652
rect 490990 138394 491018 138652
rect 491818 138394 491846 138652
rect 492646 138394 492674 138652
rect 489242 138366 489316 138394
rect 490070 138366 490144 138394
rect 490990 138366 491156 138394
rect 491818 138366 491892 138394
rect 487528 135040 487580 135046
rect 487528 134982 487580 134988
rect 487620 4208 487672 4214
rect 487620 4150 487672 4156
rect 487068 4140 487120 4146
rect 487068 4082 487120 4088
rect 486422 3632 486478 3641
rect 486422 3567 486478 3576
rect 486436 480 486464 3567
rect 487632 480 487660 4150
rect 488368 4010 488396 138366
rect 489288 135726 489316 138366
rect 490116 135726 490144 138366
rect 489276 135720 489328 135726
rect 489276 135662 489328 135668
rect 489828 135720 489880 135726
rect 489828 135662 489880 135668
rect 490104 135720 490156 135726
rect 490104 135662 490156 135668
rect 488632 135312 488684 135318
rect 488632 135254 488684 135260
rect 488644 134910 488672 135254
rect 488632 134904 488684 134910
rect 488632 134846 488684 134852
rect 489840 15910 489868 135662
rect 488816 15904 488868 15910
rect 488816 15846 488868 15852
rect 489828 15904 489880 15910
rect 489828 15846 489880 15852
rect 488356 4004 488408 4010
rect 488356 3946 488408 3952
rect 488828 480 488856 15846
rect 491024 5500 491076 5506
rect 491024 5442 491076 5448
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 489932 480 489960 3470
rect 491036 2802 491064 5442
rect 491128 3806 491156 138366
rect 491864 135726 491892 138366
rect 492600 138366 492674 138394
rect 493566 138394 493594 138652
rect 494394 138394 494422 138652
rect 495314 138394 495342 138652
rect 496142 138394 496170 138652
rect 496970 138394 496998 138652
rect 497890 138394 497918 138652
rect 498718 138394 498746 138652
rect 499546 138394 499574 138652
rect 493566 138366 494008 138394
rect 494394 138366 494468 138394
rect 495314 138366 495388 138394
rect 496142 138366 496216 138394
rect 496970 138366 497044 138394
rect 497890 138366 498056 138394
rect 498718 138366 498792 138394
rect 491208 135720 491260 135726
rect 491208 135662 491260 135668
rect 491852 135720 491904 135726
rect 491852 135662 491904 135668
rect 491220 4078 491248 135662
rect 492312 4684 492364 4690
rect 492312 4626 492364 4632
rect 491208 4072 491260 4078
rect 491208 4014 491260 4020
rect 491116 3800 491168 3806
rect 491116 3742 491168 3748
rect 491036 2774 491156 2802
rect 491128 480 491156 2774
rect 492324 480 492352 4626
rect 492600 3942 492628 138366
rect 493876 135720 493928 135726
rect 493876 135662 493928 135668
rect 493888 134638 493916 135662
rect 493876 134632 493928 134638
rect 493876 134574 493928 134580
rect 492588 3936 492640 3942
rect 492588 3878 492640 3884
rect 493980 3874 494008 138366
rect 494440 135726 494468 138366
rect 494428 135720 494480 135726
rect 494428 135662 494480 135668
rect 494704 5432 494756 5438
rect 494704 5374 494756 5380
rect 493968 3868 494020 3874
rect 493968 3810 494020 3816
rect 493506 3496 493562 3505
rect 493506 3431 493562 3440
rect 493520 480 493548 3431
rect 494716 480 494744 5374
rect 495360 3738 495388 138366
rect 496188 135454 496216 138366
rect 496176 135448 496228 135454
rect 496176 135390 496228 135396
rect 496728 135448 496780 135454
rect 496728 135390 496780 135396
rect 495900 6452 495952 6458
rect 495900 6394 495952 6400
rect 495348 3732 495400 3738
rect 495348 3674 495400 3680
rect 495912 480 495940 6394
rect 496740 3602 496768 135390
rect 497016 134570 497044 138366
rect 497004 134564 497056 134570
rect 497004 134506 497056 134512
rect 496728 3596 496780 3602
rect 496728 3538 496780 3544
rect 498028 3534 498056 138366
rect 498764 135386 498792 138366
rect 499500 138366 499574 138394
rect 500466 138394 500494 138652
rect 501294 138394 501322 138652
rect 502122 138394 502150 138652
rect 503042 138394 503070 138652
rect 503870 138394 503898 138652
rect 500466 138366 500908 138394
rect 501294 138366 501368 138394
rect 502122 138366 502288 138394
rect 503042 138366 503116 138394
rect 503870 138366 503944 138394
rect 499500 135794 499528 138366
rect 499488 135788 499540 135794
rect 499488 135730 499540 135736
rect 499580 135448 499632 135454
rect 499580 135390 499632 135396
rect 498752 135380 498804 135386
rect 498752 135322 498804 135328
rect 499488 135380 499540 135386
rect 499488 135322 499540 135328
rect 498200 5296 498252 5302
rect 498200 5238 498252 5244
rect 498016 3528 498068 3534
rect 498016 3470 498068 3476
rect 497094 3360 497150 3369
rect 497094 3295 497150 3304
rect 497108 480 497136 3295
rect 498212 480 498240 5238
rect 499396 4752 499448 4758
rect 499396 4694 499448 4700
rect 499408 480 499436 4694
rect 499500 3670 499528 135322
rect 499592 16574 499620 135390
rect 499592 16546 500632 16574
rect 499488 3664 499540 3670
rect 499488 3606 499540 3612
rect 500604 480 500632 16546
rect 500880 3777 500908 138366
rect 501340 135454 501368 138366
rect 501328 135448 501380 135454
rect 501328 135390 501380 135396
rect 502156 135448 502208 135454
rect 502156 135390 502208 135396
rect 501788 5364 501840 5370
rect 501788 5306 501840 5312
rect 500866 3768 500922 3777
rect 500866 3703 500922 3712
rect 501800 480 501828 5306
rect 502168 3641 502196 135390
rect 502154 3632 502210 3641
rect 502154 3567 502210 3576
rect 502260 3369 502288 138366
rect 503088 135454 503116 138366
rect 503916 135454 503944 138366
rect 506480 136536 506532 136542
rect 506480 136478 506532 136484
rect 503076 135448 503128 135454
rect 503076 135390 503128 135396
rect 503628 135448 503680 135454
rect 503628 135390 503680 135396
rect 503904 135448 503956 135454
rect 503904 135390 503956 135396
rect 505008 135448 505060 135454
rect 505008 135390 505060 135396
rect 502340 47592 502392 47598
rect 502340 47534 502392 47540
rect 502352 16574 502380 47534
rect 502352 16546 503024 16574
rect 502246 3360 502302 3369
rect 502246 3295 502302 3304
rect 502996 480 503024 16546
rect 503640 3505 503668 135390
rect 503626 3496 503682 3505
rect 505020 3466 505048 135390
rect 505376 5228 505428 5234
rect 505376 5170 505428 5176
rect 503626 3431 503682 3440
rect 504180 3460 504232 3466
rect 504180 3402 504232 3408
rect 505008 3460 505060 3466
rect 505008 3402 505060 3408
rect 504192 480 504220 3402
rect 505388 480 505416 5170
rect 506492 4214 506520 136478
rect 508516 86970 508544 566034
rect 511264 564868 511316 564874
rect 511264 564810 511316 564816
rect 508596 136468 508648 136474
rect 508596 136410 508648 136416
rect 508504 86964 508556 86970
rect 508504 86906 508556 86912
rect 506572 11756 506624 11762
rect 506572 11698 506624 11704
rect 506480 4208 506532 4214
rect 506480 4150 506532 4156
rect 506584 3482 506612 11698
rect 508608 4758 508636 136410
rect 511276 126954 511304 564810
rect 512656 139398 512684 567287
rect 515416 179382 515444 567394
rect 518176 219434 518204 567530
rect 519556 259418 519584 567598
rect 520936 313274 520964 567666
rect 522316 365702 522344 567802
rect 525076 419490 525104 567870
rect 533344 566500 533396 566506
rect 533344 566442 533396 566448
rect 526444 566228 526496 566234
rect 526444 566170 526496 566176
rect 525064 419484 525116 419490
rect 525064 419426 525116 419432
rect 522304 365696 522356 365702
rect 522304 365638 522356 365644
rect 520924 313268 520976 313274
rect 520924 313210 520976 313216
rect 519544 259412 519596 259418
rect 519544 259354 519596 259360
rect 518164 219428 518216 219434
rect 518164 219370 518216 219376
rect 515404 179376 515456 179382
rect 515404 179318 515456 179324
rect 526456 167006 526484 566170
rect 530584 565344 530636 565350
rect 530584 565286 530636 565292
rect 529204 565072 529256 565078
rect 529204 565014 529256 565020
rect 529216 206990 529244 565014
rect 530596 299470 530624 565286
rect 533356 353258 533384 566442
rect 537484 565616 537536 565622
rect 537484 565558 537536 565564
rect 536104 565480 536156 565486
rect 536104 565422 536156 565428
rect 536116 405686 536144 565422
rect 537496 538218 537524 565558
rect 538864 564596 538916 564602
rect 538864 564538 538916 564544
rect 537484 538212 537536 538218
rect 537484 538154 537536 538160
rect 536104 405680 536156 405686
rect 536104 405622 536156 405628
rect 533344 353252 533396 353258
rect 533344 353194 533396 353200
rect 530584 299464 530636 299470
rect 530584 299406 530636 299412
rect 529204 206984 529256 206990
rect 529204 206926 529256 206932
rect 526444 167000 526496 167006
rect 526444 166942 526496 166948
rect 512644 139392 512696 139398
rect 512644 139334 512696 139340
rect 511356 136400 511408 136406
rect 511356 136342 511408 136348
rect 511264 126948 511316 126954
rect 511264 126890 511316 126896
rect 508872 5160 508924 5166
rect 508872 5102 508924 5108
rect 508596 4752 508648 4758
rect 508596 4694 508648 4700
rect 507676 4208 507728 4214
rect 507676 4150 507728 4156
rect 506492 3454 506612 3482
rect 506492 480 506520 3454
rect 507688 480 507716 4150
rect 508884 480 508912 5102
rect 510068 4752 510120 4758
rect 510068 4694 510120 4700
rect 510080 480 510108 4694
rect 511368 4214 511396 136342
rect 529204 136332 529256 136338
rect 529204 136274 529256 136280
rect 517520 136264 517572 136270
rect 517520 136206 517572 136212
rect 512644 135652 512696 135658
rect 512644 135594 512696 135600
rect 512656 11762 512684 135594
rect 515404 135516 515456 135522
rect 515404 135458 515456 135464
rect 512644 11756 512696 11762
rect 512644 11698 512696 11704
rect 512460 5092 512512 5098
rect 512460 5034 512512 5040
rect 511356 4208 511408 4214
rect 511356 4150 511408 4156
rect 511264 2848 511316 2854
rect 511264 2790 511316 2796
rect 511276 480 511304 2790
rect 512472 480 512500 5034
rect 515416 5030 515444 135458
rect 517532 16574 517560 136206
rect 524420 136060 524472 136066
rect 524420 136002 524472 136008
rect 520924 135856 520976 135862
rect 520924 135798 520976 135804
rect 519544 135584 519596 135590
rect 519544 135526 519596 135532
rect 517532 16546 517928 16574
rect 517152 6520 517204 6526
rect 517152 6462 517204 6468
rect 515404 5024 515456 5030
rect 515404 4966 515456 4972
rect 515956 4956 516008 4962
rect 515956 4898 516008 4904
rect 513564 4208 513616 4214
rect 513564 4150 513616 4156
rect 513576 480 513604 4150
rect 514760 2916 514812 2922
rect 514760 2858 514812 2864
rect 514772 480 514800 2858
rect 515968 480 515996 4898
rect 517164 480 517192 6462
rect 517900 490 517928 16546
rect 519556 6458 519584 135526
rect 520280 134972 520332 134978
rect 520280 134914 520332 134920
rect 519544 6452 519596 6458
rect 519544 6394 519596 6400
rect 519544 4752 519596 4758
rect 519544 4694 519596 4700
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 4694
rect 520292 490 520320 134914
rect 520936 7682 520964 135798
rect 522304 135720 522356 135726
rect 522304 135662 522356 135668
rect 520924 7676 520976 7682
rect 520924 7618 520976 7624
rect 522316 7614 522344 135662
rect 524432 16574 524460 136002
rect 526444 135788 526496 135794
rect 526444 135730 526496 135736
rect 524432 16546 525472 16574
rect 522304 7608 522356 7614
rect 522304 7550 522356 7556
rect 524236 6384 524288 6390
rect 524236 6326 524288 6332
rect 523040 4820 523092 4826
rect 523040 4762 523092 4768
rect 521844 2984 521896 2990
rect 521844 2926 521896 2932
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 2926
rect 523052 480 523080 4762
rect 524248 480 524276 6326
rect 525444 480 525472 16546
rect 526456 10334 526484 135730
rect 526444 10328 526496 10334
rect 526444 10270 526496 10276
rect 527824 6316 527876 6322
rect 527824 6258 527876 6264
rect 526628 4888 526680 4894
rect 526628 4830 526680 4836
rect 526640 480 526668 4830
rect 527836 480 527864 6258
rect 529216 4214 529244 136274
rect 536104 136128 536156 136134
rect 536104 136070 536156 136076
rect 531320 135992 531372 135998
rect 531320 135934 531372 135940
rect 531332 16574 531360 135934
rect 531332 16546 532096 16574
rect 530124 11756 530176 11762
rect 530124 11698 530176 11704
rect 529204 4208 529256 4214
rect 529204 4150 529256 4156
rect 529020 3052 529072 3058
rect 529020 2994 529072 3000
rect 529032 480 529060 2994
rect 530136 480 530164 11698
rect 531320 6248 531372 6254
rect 531320 6190 531372 6196
rect 531332 480 531360 6190
rect 532068 490 532096 16546
rect 533712 8968 533764 8974
rect 533712 8910 533764 8916
rect 532344 598 532556 626
rect 532344 490 532372 598
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 462 532372 490
rect 532528 480 532556 598
rect 533724 480 533752 8910
rect 536116 4826 536144 136070
rect 538876 113150 538904 564538
rect 540256 153202 540284 568754
rect 543016 193186 543044 568890
rect 544382 564224 544438 564233
rect 544382 564159 544438 564168
rect 544396 233238 544424 564159
rect 547156 273222 547184 568958
rect 548524 566636 548576 566642
rect 548524 566578 548576 566584
rect 548536 485790 548564 566578
rect 551284 566160 551336 566166
rect 551284 566102 551336 566108
rect 548524 485784 548576 485790
rect 548524 485726 548576 485732
rect 547144 273216 547196 273222
rect 547144 273158 547196 273164
rect 551296 245614 551324 566102
rect 555422 564360 555478 564369
rect 555422 564295 555478 564304
rect 555436 325650 555464 564295
rect 556816 379506 556844 569026
rect 558184 568676 558236 568682
rect 558184 568618 558236 568624
rect 556804 379500 556856 379506
rect 556804 379442 556856 379448
rect 555424 325644 555476 325650
rect 555424 325586 555476 325592
rect 551284 245608 551336 245614
rect 551284 245550 551336 245556
rect 544384 233232 544436 233238
rect 544384 233174 544436 233180
rect 543004 193180 543056 193186
rect 543004 193122 543056 193128
rect 540244 153196 540296 153202
rect 540244 153138 540296 153144
rect 543004 136196 543056 136202
rect 543004 136138 543056 136144
rect 539600 135924 539652 135930
rect 539600 135866 539652 135872
rect 538864 113144 538916 113150
rect 538864 113086 538916 113092
rect 538220 49020 538272 49026
rect 538220 48962 538272 48968
rect 538232 16574 538260 48962
rect 538232 16546 538444 16574
rect 537208 14476 537260 14482
rect 537208 14418 537260 14424
rect 536104 4820 536156 4826
rect 536104 4762 536156 4768
rect 534908 4208 534960 4214
rect 534908 4150 534960 4156
rect 534920 480 534948 4150
rect 536104 3120 536156 3126
rect 536104 3062 536156 3068
rect 536116 480 536144 3062
rect 537220 480 537248 14418
rect 538416 480 538444 16546
rect 539612 480 539640 135866
rect 540796 5024 540848 5030
rect 540796 4966 540848 4972
rect 540808 480 540836 4966
rect 543016 4826 543044 136138
rect 547144 135040 547196 135046
rect 547144 134982 547196 134988
rect 544384 134836 544436 134842
rect 544384 134778 544436 134784
rect 544292 6452 544344 6458
rect 544292 6394 544344 6400
rect 541992 4820 542044 4826
rect 541992 4762 542044 4768
rect 543004 4820 543056 4826
rect 543004 4762 543056 4768
rect 542004 480 542032 4762
rect 544304 3210 544332 6394
rect 544396 3330 544424 134778
rect 544384 3324 544436 3330
rect 544384 3266 544436 3272
rect 545488 3324 545540 3330
rect 545488 3266 545540 3272
rect 544304 3182 544424 3210
rect 543188 3120 543240 3126
rect 543188 3062 543240 3068
rect 543200 480 543228 3062
rect 544396 480 544424 3182
rect 545500 480 545528 3266
rect 547156 3262 547184 134982
rect 550640 134904 550692 134910
rect 550640 134846 550692 134852
rect 547880 134768 547932 134774
rect 547880 134710 547932 134716
rect 547144 3256 547196 3262
rect 547144 3198 547196 3204
rect 546684 3052 546736 3058
rect 546684 2994 546736 3000
rect 546696 480 546724 2994
rect 547892 480 547920 134710
rect 550652 16574 550680 134846
rect 554780 134700 554832 134706
rect 554780 134642 554832 134648
rect 554792 16574 554820 134642
rect 556252 133204 556304 133210
rect 556252 133146 556304 133152
rect 550652 16546 551048 16574
rect 554792 16546 555004 16574
rect 549076 6180 549128 6186
rect 549076 6122 549128 6128
rect 549088 480 549116 6122
rect 550272 3188 550324 3194
rect 550272 3130 550324 3136
rect 550284 480 550312 3130
rect 551020 490 551048 16546
rect 552664 4820 552716 4826
rect 552664 4762 552716 4768
rect 551296 598 551508 626
rect 551296 490 551324 598
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 462 551324 490
rect 551480 480 551508 598
rect 552676 480 552704 4762
rect 553768 3392 553820 3398
rect 553768 3334 553820 3340
rect 553780 480 553808 3334
rect 554976 480 555004 16546
rect 556264 6914 556292 133146
rect 558196 60722 558224 568618
rect 558932 568070 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 560944 568744 560996 568750
rect 560944 568686 560996 568692
rect 558920 568064 558972 568070
rect 558920 568006 558972 568012
rect 560956 100706 560984 568686
rect 580448 565412 580500 565418
rect 580448 565354 580500 565360
rect 580356 565208 580408 565214
rect 580356 565150 580408 565156
rect 580264 564936 580316 564942
rect 580264 564878 580316 564884
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580276 431633 580304 564878
rect 580368 471481 580396 565150
rect 580460 524521 580488 565354
rect 580446 524512 580502 524521
rect 580446 524447 580502 524456
rect 580354 471472 580410 471481
rect 580354 471407 580410 471416
rect 580262 431624 580318 431633
rect 580262 431559 580318 431568
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 564532 134632 564584 134638
rect 564532 134574 564584 134580
rect 560944 100700 560996 100706
rect 560944 100642 560996 100648
rect 558184 60716 558236 60722
rect 558184 60658 558236 60664
rect 564544 16574 564572 134574
rect 572812 134564 572864 134570
rect 572812 134506 572864 134512
rect 564544 16546 565216 16574
rect 562048 15904 562100 15910
rect 562048 15846 562100 15852
rect 558552 7676 558604 7682
rect 558552 7618 558604 7624
rect 556172 6886 556292 6914
rect 556172 480 556200 6886
rect 557356 4140 557408 4146
rect 557356 4082 557408 4088
rect 557368 480 557396 4082
rect 558564 480 558592 7618
rect 560852 4004 560904 4010
rect 560852 3946 560904 3952
rect 559748 3256 559800 3262
rect 559748 3198 559800 3204
rect 559760 480 559788 3198
rect 560864 480 560892 3946
rect 562060 480 562088 15846
rect 563244 4072 563296 4078
rect 563244 4014 563296 4020
rect 563256 480 563284 4014
rect 564440 3800 564492 3806
rect 564440 3742 564492 3748
rect 564452 480 564480 3742
rect 565188 490 565216 16546
rect 569132 7608 569184 7614
rect 569132 7550 569184 7556
rect 566832 3936 566884 3942
rect 566832 3878 566884 3884
rect 565464 598 565676 626
rect 565464 490 565492 598
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 462 565492 490
rect 565648 480 565676 598
rect 566844 480 566872 3878
rect 568028 3868 568080 3874
rect 568028 3810 568080 3816
rect 568040 480 568068 3810
rect 569144 480 569172 7550
rect 572824 6914 572852 134506
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 575848 10328 575900 10334
rect 575848 10270 575900 10276
rect 572732 6886 572852 6914
rect 570328 3732 570380 3738
rect 570328 3674 570380 3680
rect 570340 480 570368 3674
rect 571524 3596 571576 3602
rect 571524 3538 571576 3544
rect 571536 480 571564 3538
rect 572732 480 572760 6886
rect 575112 3664 575164 3670
rect 575112 3606 575164 3612
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 573928 480 573956 3470
rect 575124 480 575152 3606
rect 575860 490 575888 10270
rect 577410 3768 577466 3777
rect 577410 3703 577466 3712
rect 576136 598 576348 626
rect 576136 490 576164 598
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 462 576164 490
rect 576320 480 576348 598
rect 577424 480 577452 3703
rect 578606 3632 578662 3641
rect 578606 3567 578662 3576
rect 578620 480 578648 3567
rect 582194 3496 582250 3505
rect 582194 3431 582250 3440
rect 583392 3460 583444 3466
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582208 480 582236 3431
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3330 553832 3386 553888
rect 3238 527856 3294 527912
rect 3238 501744 3294 501800
rect 3330 475632 3386 475688
rect 3330 449520 3386 449576
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 397432 3386 397488
rect 3330 371320 3386 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3054 293120 3110 293176
rect 2778 254088 2834 254144
rect 3330 214920 3386 214976
rect 2778 201864 2834 201920
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 3790 514800 3846 514856
rect 3698 462576 3754 462632
rect 3606 410488 3662 410544
rect 3514 306176 3570 306232
rect 3514 267144 3570 267200
rect 3514 241032 3570 241088
rect 11702 563760 11758 563816
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3514 71576 3570 71632
rect 3422 58520 3478 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 6458 3304 6514 3360
rect 22742 567432 22798 567488
rect 14738 3576 14794 3632
rect 15934 3440 15990 3496
rect 25502 563896 25558 563952
rect 39302 564032 39358 564088
rect 33782 563624 33838 563680
rect 20626 3712 20682 3768
rect 122746 567296 122802 567352
rect 479798 567432 479854 567488
rect 512642 567296 512698 567352
rect 81990 564576 82046 564632
rect 85026 564576 85082 564632
rect 89350 564576 89406 564632
rect 93122 564576 93178 564632
rect 96342 564576 96398 564632
rect 141514 564576 141570 564632
rect 163778 564576 163834 564632
rect 216034 564576 216090 564632
rect 465078 564576 465134 564632
rect 476118 564576 476174 564632
rect 487342 564576 487398 564632
rect 498566 564576 498622 564632
rect 84382 3304 84438 3360
rect 90454 3576 90510 3632
rect 91282 3440 91338 3496
rect 94778 3712 94834 3768
rect 390374 3304 390430 3360
rect 426162 3304 426218 3360
rect 429014 3712 429070 3768
rect 434626 3576 434682 3632
rect 440146 3440 440202 3496
rect 442906 3304 442962 3360
rect 479338 3712 479394 3768
rect 486422 3576 486478 3632
rect 493506 3440 493562 3496
rect 497094 3304 497150 3360
rect 500866 3712 500922 3768
rect 502154 3576 502210 3632
rect 502246 3304 502302 3360
rect 503626 3440 503682 3496
rect 544382 564168 544438 564224
rect 555422 564304 555478 564360
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 580170 537784 580226 537840
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580446 524456 580502 524512
rect 580354 471416 580410 471472
rect 580262 431568 580318 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 59608 580226 59664
rect 577410 3712 577466 3768
rect 578606 3576 578662 3632
rect 582194 3440 582250 3496
rect 580998 3304 581054 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 22737 567490 22803 567493
rect 479793 567490 479859 567493
rect 22737 567488 479859 567490
rect 22737 567432 22742 567488
rect 22798 567432 479798 567488
rect 479854 567432 479859 567488
rect 22737 567430 479859 567432
rect 22737 567427 22803 567430
rect 479793 567427 479859 567430
rect 122741 567354 122807 567357
rect 512637 567354 512703 567357
rect 122741 567352 512703 567354
rect 122741 567296 122746 567352
rect 122802 567296 512642 567352
rect 512698 567296 512703 567352
rect 122741 567294 512703 567296
rect 122741 567291 122807 567294
rect 512637 567291 512703 567294
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 81985 564634 82051 564637
rect 82670 564634 82676 564636
rect 81985 564632 82676 564634
rect 81985 564576 81990 564632
rect 82046 564576 82676 564632
rect 81985 564574 82676 564576
rect 81985 564571 82051 564574
rect 82670 564572 82676 564574
rect 82740 564572 82746 564636
rect 84694 564572 84700 564636
rect 84764 564634 84770 564636
rect 85021 564634 85087 564637
rect 84764 564632 85087 564634
rect 84764 564576 85026 564632
rect 85082 564576 85087 564632
rect 84764 564574 85087 564576
rect 84764 564572 84770 564574
rect 85021 564571 85087 564574
rect 89345 564634 89411 564637
rect 89478 564634 89484 564636
rect 89345 564632 89484 564634
rect 89345 564576 89350 564632
rect 89406 564576 89484 564632
rect 89345 564574 89484 564576
rect 89345 564571 89411 564574
rect 89478 564572 89484 564574
rect 89548 564572 89554 564636
rect 93117 564634 93183 564637
rect 93710 564634 93716 564636
rect 93117 564632 93716 564634
rect 93117 564576 93122 564632
rect 93178 564576 93716 564632
rect 93117 564574 93716 564576
rect 93117 564571 93183 564574
rect 93710 564572 93716 564574
rect 93780 564572 93786 564636
rect 96337 564634 96403 564637
rect 96470 564634 96476 564636
rect 96337 564632 96476 564634
rect 96337 564576 96342 564632
rect 96398 564576 96476 564632
rect 96337 564574 96476 564576
rect 96337 564571 96403 564574
rect 96470 564572 96476 564574
rect 96540 564572 96546 564636
rect 141509 564634 141575 564637
rect 163773 564634 163839 564637
rect 216029 564636 216095 564637
rect 465073 564636 465139 564637
rect 476113 564636 476179 564637
rect 487337 564636 487403 564637
rect 498561 564636 498627 564637
rect 141509 564632 141618 564634
rect 141509 564576 141514 564632
rect 141570 564576 141618 564632
rect 141509 564571 141618 564576
rect 163773 564632 163882 564634
rect 163773 564576 163778 564632
rect 163834 564576 163882 564632
rect 163773 564571 163882 564576
rect 216029 564632 216076 564636
rect 216140 564634 216146 564636
rect 465022 564634 465028 564636
rect 216029 564576 216034 564632
rect 216029 564572 216076 564576
rect 216140 564574 216186 564634
rect 464982 564574 465028 564634
rect 465092 564632 465139 564636
rect 476062 564634 476068 564636
rect 465134 564576 465139 564632
rect 216140 564572 216146 564574
rect 465022 564572 465028 564574
rect 465092 564572 465139 564576
rect 476022 564574 476068 564634
rect 476132 564632 476179 564636
rect 487286 564634 487292 564636
rect 476174 564576 476179 564632
rect 476062 564572 476068 564574
rect 476132 564572 476179 564576
rect 487246 564574 487292 564634
rect 487356 564632 487403 564636
rect 498510 564634 498516 564636
rect 487398 564576 487403 564632
rect 487286 564572 487292 564574
rect 487356 564572 487403 564576
rect 498470 564574 498516 564634
rect 498580 564632 498627 564636
rect 498622 564576 498627 564632
rect 498510 564572 498516 564574
rect 498580 564572 498627 564576
rect 216029 564571 216095 564572
rect 465073 564571 465139 564572
rect 476113 564571 476179 564572
rect 487337 564571 487403 564572
rect 498561 564571 498627 564572
rect 141558 564226 141618 564571
rect 163822 564362 163882 564571
rect 555417 564362 555483 564365
rect 583520 564362 584960 564452
rect 163822 564360 555483 564362
rect 163822 564304 555422 564360
rect 555478 564304 555483 564360
rect 163822 564302 555483 564304
rect 555417 564299 555483 564302
rect 583342 564302 584960 564362
rect 544377 564226 544443 564229
rect 141558 564224 544443 564226
rect 141558 564168 544382 564224
rect 544438 564168 544443 564224
rect 141558 564166 544443 564168
rect 583342 564226 583402 564302
rect 583520 564226 584960 564302
rect 583342 564212 584960 564226
rect 583342 564166 583586 564212
rect 544377 564163 544443 564166
rect 39297 564090 39363 564093
rect 487286 564090 487292 564092
rect 39297 564088 487292 564090
rect 39297 564032 39302 564088
rect 39358 564032 487292 564088
rect 39297 564030 487292 564032
rect 39297 564027 39363 564030
rect 487286 564028 487292 564030
rect 487356 564028 487362 564092
rect 25497 563954 25563 563957
rect 476062 563954 476068 563956
rect 25497 563952 476068 563954
rect 25497 563896 25502 563952
rect 25558 563896 476068 563952
rect 25497 563894 476068 563896
rect 25497 563891 25563 563894
rect 476062 563892 476068 563894
rect 476132 563892 476138 563956
rect 11697 563818 11763 563821
rect 465022 563818 465028 563820
rect 11697 563816 465028 563818
rect 11697 563760 11702 563816
rect 11758 563760 465028 563816
rect 11697 563758 465028 563760
rect 11697 563755 11763 563758
rect 465022 563756 465028 563758
rect 465092 563756 465098 563820
rect 33777 563682 33843 563685
rect 498510 563682 498516 563684
rect 33777 563680 498516 563682
rect 33777 563624 33782 563680
rect 33838 563624 498516 563680
rect 33777 563622 498516 563624
rect 33777 563619 33843 563622
rect 498510 563620 498516 563622
rect 498580 563620 498586 563684
rect 216070 563076 216076 563140
rect 216140 563138 216146 563140
rect 583526 563138 583586 564166
rect 216140 563078 583586 563138
rect 216140 563076 216146 563078
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3233 527914 3299 527917
rect -960 527912 3299 527914
rect -960 527856 3238 527912
rect 3294 527856 3299 527912
rect -960 527854 3299 527856
rect -960 527764 480 527854
rect 3233 527851 3299 527854
rect 580441 524514 580507 524517
rect 583520 524514 584960 524604
rect 580441 524512 584960 524514
rect 580441 524456 580446 524512
rect 580502 524456 584960 524512
rect 580441 524454 584960 524456
rect 580441 524451 580507 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3785 514858 3851 514861
rect -960 514856 3851 514858
rect -960 514800 3790 514856
rect 3846 514800 3851 514856
rect -960 514798 3851 514800
rect -960 514708 480 514798
rect 3785 514795 3851 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 580349 471474 580415 471477
rect 583520 471474 584960 471564
rect 580349 471472 584960 471474
rect 580349 471416 580354 471472
rect 580410 471416 584960 471472
rect 580349 471414 584960 471416
rect 580349 471411 580415 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3693 462634 3759 462637
rect -960 462632 3759 462634
rect -960 462576 3698 462632
rect 3754 462576 3759 462632
rect -960 462574 3759 462576
rect -960 462484 480 462574
rect 3693 462571 3759 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580257 431626 580323 431629
rect 583520 431626 584960 431716
rect 580257 431624 584960 431626
rect 580257 431568 580262 431624
rect 580318 431568 584960 431624
rect 580257 431566 584960 431568
rect 580257 431563 580323 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3601 410546 3667 410549
rect -960 410544 3667 410546
rect -960 410488 3606 410544
rect 3662 410488 3667 410544
rect -960 410486 3667 410488
rect -960 410396 480 410486
rect 3601 410483 3667 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 96470 71844 96476 71908
rect 96540 71906 96546 71908
rect 583526 71906 583586 72798
rect 96540 71846 583586 71906
rect 96540 71844 96546 71846
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 93710 45596 93716 45660
rect 93780 45658 93786 45660
rect 583526 45658 583586 46142
rect 93780 45598 583586 45658
rect 93780 45596 93786 45598
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 84694 31724 84700 31788
rect 84764 31786 84770 31788
rect 583526 31786 583586 32950
rect 84764 31726 583586 31786
rect 84764 31724 84770 31726
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 89478 19348 89484 19412
rect 89548 19410 89554 19412
rect 583526 19410 583586 19622
rect 89548 19350 583586 19410
rect 89548 19348 89554 19350
rect 583520 6626 584960 6716
rect -960 6490 480 6580
rect 583342 6566 584960 6626
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect 583342 6490 583402 6566
rect 583520 6490 584960 6566
rect 583342 6476 584960 6490
rect 583342 6430 583586 6476
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 82670 5612 82676 5676
rect 82740 5674 82746 5676
rect 583526 5674 583586 6430
rect 82740 5614 583586 5674
rect 82740 5612 82746 5614
rect 20621 3770 20687 3773
rect 94773 3770 94839 3773
rect 20621 3768 94839 3770
rect 20621 3712 20626 3768
rect 20682 3712 94778 3768
rect 94834 3712 94839 3768
rect 20621 3710 94839 3712
rect 20621 3707 20687 3710
rect 94773 3707 94839 3710
rect 429009 3770 429075 3773
rect 479333 3770 479399 3773
rect 429009 3768 479399 3770
rect 429009 3712 429014 3768
rect 429070 3712 479338 3768
rect 479394 3712 479399 3768
rect 429009 3710 479399 3712
rect 429009 3707 429075 3710
rect 479333 3707 479399 3710
rect 500861 3770 500927 3773
rect 577405 3770 577471 3773
rect 500861 3768 577471 3770
rect 500861 3712 500866 3768
rect 500922 3712 577410 3768
rect 577466 3712 577471 3768
rect 500861 3710 577471 3712
rect 500861 3707 500927 3710
rect 577405 3707 577471 3710
rect 14733 3634 14799 3637
rect 90449 3634 90515 3637
rect 14733 3632 90515 3634
rect 14733 3576 14738 3632
rect 14794 3576 90454 3632
rect 90510 3576 90515 3632
rect 14733 3574 90515 3576
rect 14733 3571 14799 3574
rect 90449 3571 90515 3574
rect 434621 3634 434687 3637
rect 486417 3634 486483 3637
rect 434621 3632 486483 3634
rect 434621 3576 434626 3632
rect 434682 3576 486422 3632
rect 486478 3576 486483 3632
rect 434621 3574 486483 3576
rect 434621 3571 434687 3574
rect 486417 3571 486483 3574
rect 502149 3634 502215 3637
rect 578601 3634 578667 3637
rect 502149 3632 578667 3634
rect 502149 3576 502154 3632
rect 502210 3576 578606 3632
rect 578662 3576 578667 3632
rect 502149 3574 578667 3576
rect 502149 3571 502215 3574
rect 578601 3571 578667 3574
rect 15929 3498 15995 3501
rect 91277 3498 91343 3501
rect 15929 3496 91343 3498
rect 15929 3440 15934 3496
rect 15990 3440 91282 3496
rect 91338 3440 91343 3496
rect 15929 3438 91343 3440
rect 15929 3435 15995 3438
rect 91277 3435 91343 3438
rect 440141 3498 440207 3501
rect 493501 3498 493567 3501
rect 440141 3496 493567 3498
rect 440141 3440 440146 3496
rect 440202 3440 493506 3496
rect 493562 3440 493567 3496
rect 440141 3438 493567 3440
rect 440141 3435 440207 3438
rect 493501 3435 493567 3438
rect 503621 3498 503687 3501
rect 582189 3498 582255 3501
rect 503621 3496 582255 3498
rect 503621 3440 503626 3496
rect 503682 3440 582194 3496
rect 582250 3440 582255 3496
rect 503621 3438 582255 3440
rect 503621 3435 503687 3438
rect 582189 3435 582255 3438
rect 6453 3362 6519 3365
rect 84377 3362 84443 3365
rect 6453 3360 84443 3362
rect 6453 3304 6458 3360
rect 6514 3304 84382 3360
rect 84438 3304 84443 3360
rect 6453 3302 84443 3304
rect 6453 3299 6519 3302
rect 84377 3299 84443 3302
rect 390369 3362 390435 3365
rect 426157 3362 426223 3365
rect 390369 3360 426223 3362
rect 390369 3304 390374 3360
rect 390430 3304 426162 3360
rect 426218 3304 426223 3360
rect 390369 3302 426223 3304
rect 390369 3299 390435 3302
rect 426157 3299 426223 3302
rect 442901 3362 442967 3365
rect 497089 3362 497155 3365
rect 442901 3360 497155 3362
rect 442901 3304 442906 3360
rect 442962 3304 497094 3360
rect 497150 3304 497155 3360
rect 442901 3302 497155 3304
rect 442901 3299 442967 3302
rect 497089 3299 497155 3302
rect 502241 3362 502307 3365
rect 580993 3362 581059 3365
rect 502241 3360 581059 3362
rect 502241 3304 502246 3360
rect 502302 3304 580998 3360
rect 581054 3304 581059 3360
rect 502241 3302 581059 3304
rect 502241 3299 502307 3302
rect 580993 3299 581059 3302
<< via3 >>
rect 82676 564572 82740 564636
rect 84700 564572 84764 564636
rect 89484 564572 89548 564636
rect 93716 564572 93780 564636
rect 96476 564572 96540 564636
rect 216076 564632 216140 564636
rect 216076 564576 216090 564632
rect 216090 564576 216140 564632
rect 216076 564572 216140 564576
rect 465028 564632 465092 564636
rect 465028 564576 465078 564632
rect 465078 564576 465092 564632
rect 465028 564572 465092 564576
rect 476068 564632 476132 564636
rect 476068 564576 476118 564632
rect 476118 564576 476132 564632
rect 476068 564572 476132 564576
rect 487292 564632 487356 564636
rect 487292 564576 487342 564632
rect 487342 564576 487356 564632
rect 487292 564572 487356 564576
rect 498516 564632 498580 564636
rect 498516 564576 498566 564632
rect 498566 564576 498580 564632
rect 498516 564572 498580 564576
rect 487292 564028 487356 564092
rect 476068 563892 476132 563956
rect 465028 563756 465092 563820
rect 498516 563620 498580 563684
rect 216076 563076 216140 563140
rect 96476 71844 96540 71908
rect 93716 45596 93780 45660
rect 84700 31724 84764 31788
rect 89484 19348 89548 19412
rect 82676 5612 82740 5676
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 567304 78134 582618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 567304 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 567304 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 567304 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 567304 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 567304 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 567304 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 567304 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 567304 114134 582618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 567304 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 567304 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 567304 128414 596898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 567304 132134 600618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 567304 135854 568338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 567304 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 567304 146414 578898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 567304 150134 582618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 567304 153854 586338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 567304 157574 590058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 567304 164414 596898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 567304 168134 600618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 567304 171854 568338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 567304 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 567304 182414 578898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 567304 186134 582618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 567304 189854 586338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 567304 193574 590058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 567304 200414 596898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 567304 204134 600618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 567304 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 567304 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 567304 218414 578898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 567304 222134 582618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 567304 225854 586338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 567304 229574 590058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 567304 236414 596898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 567304 240134 600618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 567304 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 567304 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 567304 254414 578898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 567304 258134 582618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 567304 261854 586338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 567304 265574 590058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 567304 272414 596898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 567304 276134 600618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 567304 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 567304 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 567304 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 567304 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 567304 297854 586338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 567304 301574 590058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 567304 308414 596898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 567304 312134 600618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 567304 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 567304 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 567304 326414 578898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 567304 330134 582618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 567304 333854 586338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 567304 337574 590058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 567304 344414 596898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 567304 348134 600618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 567304 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 567304 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 567304 362414 578898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 567304 366134 582618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 567304 369854 586338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 567304 373574 590058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 567304 380414 596898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 567304 384134 600618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 567304 387854 568338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 567304 391574 572058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 567304 398414 578898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 567304 402134 582618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 567304 405854 586338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 567304 409574 590058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 567304 416414 596898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 567304 420134 600618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 567304 423854 568338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 567304 427574 572058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 567304 434414 578898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 567304 438134 582618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 567304 441854 586338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 567304 445574 590058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 567304 452414 596898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 567304 456134 600618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 567304 459854 568338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 567304 463574 572058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 567304 470414 578898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 567304 474134 582618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 567304 477854 586338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 567304 481574 590058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 567304 488414 596898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 567304 492134 600618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 567304 495854 568338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 567304 499574 572058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 567304 506414 578898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 82675 564636 82741 564637
rect 82675 564572 82676 564636
rect 82740 564572 82741 564636
rect 82675 564571 82741 564572
rect 84699 564636 84765 564637
rect 84699 564572 84700 564636
rect 84764 564572 84765 564636
rect 84699 564571 84765 564572
rect 89483 564636 89549 564637
rect 89483 564572 89484 564636
rect 89548 564572 89549 564636
rect 89483 564571 89549 564572
rect 93715 564636 93781 564637
rect 93715 564572 93716 564636
rect 93780 564572 93781 564636
rect 93715 564571 93781 564572
rect 96475 564636 96541 564637
rect 96475 564572 96476 564636
rect 96540 564572 96541 564636
rect 96475 564571 96541 564572
rect 216075 564636 216141 564637
rect 216075 564572 216076 564636
rect 216140 564572 216141 564636
rect 216075 564571 216141 564572
rect 465027 564636 465093 564637
rect 465027 564572 465028 564636
rect 465092 564572 465093 564636
rect 465027 564571 465093 564572
rect 476067 564636 476133 564637
rect 476067 564572 476068 564636
rect 476132 564572 476133 564636
rect 476067 564571 476133 564572
rect 487291 564636 487357 564637
rect 487291 564572 487292 564636
rect 487356 564572 487357 564636
rect 487291 564571 487357 564572
rect 498515 564636 498581 564637
rect 498515 564572 498516 564636
rect 498580 564572 498581 564636
rect 498515 564571 498581 564572
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 115174 78134 136600
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 118894 81854 136600
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 82678 5677 82738 564571
rect 84008 543454 84328 543486
rect 84008 543218 84050 543454
rect 84286 543218 84328 543454
rect 84008 543134 84328 543218
rect 84008 542898 84050 543134
rect 84286 542898 84328 543134
rect 84008 542866 84328 542898
rect 84008 507454 84328 507486
rect 84008 507218 84050 507454
rect 84286 507218 84328 507454
rect 84008 507134 84328 507218
rect 84008 506898 84050 507134
rect 84286 506898 84328 507134
rect 84008 506866 84328 506898
rect 84008 471454 84328 471486
rect 84008 471218 84050 471454
rect 84286 471218 84328 471454
rect 84008 471134 84328 471218
rect 84008 470898 84050 471134
rect 84286 470898 84328 471134
rect 84008 470866 84328 470898
rect 84008 435454 84328 435486
rect 84008 435218 84050 435454
rect 84286 435218 84328 435454
rect 84008 435134 84328 435218
rect 84008 434898 84050 435134
rect 84286 434898 84328 435134
rect 84008 434866 84328 434898
rect 84008 399454 84328 399486
rect 84008 399218 84050 399454
rect 84286 399218 84328 399454
rect 84008 399134 84328 399218
rect 84008 398898 84050 399134
rect 84286 398898 84328 399134
rect 84008 398866 84328 398898
rect 84008 363454 84328 363486
rect 84008 363218 84050 363454
rect 84286 363218 84328 363454
rect 84008 363134 84328 363218
rect 84008 362898 84050 363134
rect 84286 362898 84328 363134
rect 84008 362866 84328 362898
rect 84008 327454 84328 327486
rect 84008 327218 84050 327454
rect 84286 327218 84328 327454
rect 84008 327134 84328 327218
rect 84008 326898 84050 327134
rect 84286 326898 84328 327134
rect 84008 326866 84328 326898
rect 84008 291454 84328 291486
rect 84008 291218 84050 291454
rect 84286 291218 84328 291454
rect 84008 291134 84328 291218
rect 84008 290898 84050 291134
rect 84286 290898 84328 291134
rect 84008 290866 84328 290898
rect 84008 255454 84328 255486
rect 84008 255218 84050 255454
rect 84286 255218 84328 255454
rect 84008 255134 84328 255218
rect 84008 254898 84050 255134
rect 84286 254898 84328 255134
rect 84008 254866 84328 254898
rect 84008 219454 84328 219486
rect 84008 219218 84050 219454
rect 84286 219218 84328 219454
rect 84008 219134 84328 219218
rect 84008 218898 84050 219134
rect 84286 218898 84328 219134
rect 84008 218866 84328 218898
rect 84008 183454 84328 183486
rect 84008 183218 84050 183454
rect 84286 183218 84328 183454
rect 84008 183134 84328 183218
rect 84008 182898 84050 183134
rect 84286 182898 84328 183134
rect 84008 182866 84328 182898
rect 84008 147454 84328 147486
rect 84008 147218 84050 147454
rect 84286 147218 84328 147454
rect 84008 147134 84328 147218
rect 84008 146898 84050 147134
rect 84286 146898 84328 147134
rect 84008 146866 84328 146898
rect 84702 31789 84762 564571
rect 84954 122614 85574 136600
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84699 31788 84765 31789
rect 84699 31724 84700 31788
rect 84764 31724 84765 31788
rect 84699 31723 84765 31724
rect 84954 14614 85574 50058
rect 89486 19413 89546 564571
rect 91794 129454 92414 136600
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 93718 45661 93778 564571
rect 95514 133174 96134 136600
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 96478 71909 96538 564571
rect 216078 563141 216138 564571
rect 465030 563821 465090 564571
rect 476070 563957 476130 564571
rect 487294 564093 487354 564571
rect 487291 564092 487357 564093
rect 487291 564028 487292 564092
rect 487356 564028 487357 564092
rect 487291 564027 487357 564028
rect 476067 563956 476133 563957
rect 476067 563892 476068 563956
rect 476132 563892 476133 563956
rect 476067 563891 476133 563892
rect 465027 563820 465093 563821
rect 465027 563756 465028 563820
rect 465092 563756 465093 563820
rect 465027 563755 465093 563756
rect 498518 563685 498578 564571
rect 498515 563684 498581 563685
rect 498515 563620 498516 563684
rect 498580 563620 498581 563684
rect 498515 563619 498581 563620
rect 216075 563140 216141 563141
rect 216075 563076 216076 563140
rect 216140 563076 216141 563140
rect 216075 563075 216141 563076
rect 99368 561454 99688 561486
rect 99368 561218 99410 561454
rect 99646 561218 99688 561454
rect 99368 561134 99688 561218
rect 99368 560898 99410 561134
rect 99646 560898 99688 561134
rect 99368 560866 99688 560898
rect 130088 561454 130408 561486
rect 130088 561218 130130 561454
rect 130366 561218 130408 561454
rect 130088 561134 130408 561218
rect 130088 560898 130130 561134
rect 130366 560898 130408 561134
rect 130088 560866 130408 560898
rect 160808 561454 161128 561486
rect 160808 561218 160850 561454
rect 161086 561218 161128 561454
rect 160808 561134 161128 561218
rect 160808 560898 160850 561134
rect 161086 560898 161128 561134
rect 160808 560866 161128 560898
rect 191528 561454 191848 561486
rect 191528 561218 191570 561454
rect 191806 561218 191848 561454
rect 191528 561134 191848 561218
rect 191528 560898 191570 561134
rect 191806 560898 191848 561134
rect 191528 560866 191848 560898
rect 222248 561454 222568 561486
rect 222248 561218 222290 561454
rect 222526 561218 222568 561454
rect 222248 561134 222568 561218
rect 222248 560898 222290 561134
rect 222526 560898 222568 561134
rect 222248 560866 222568 560898
rect 252968 561454 253288 561486
rect 252968 561218 253010 561454
rect 253246 561218 253288 561454
rect 252968 561134 253288 561218
rect 252968 560898 253010 561134
rect 253246 560898 253288 561134
rect 252968 560866 253288 560898
rect 283688 561454 284008 561486
rect 283688 561218 283730 561454
rect 283966 561218 284008 561454
rect 283688 561134 284008 561218
rect 283688 560898 283730 561134
rect 283966 560898 284008 561134
rect 283688 560866 284008 560898
rect 314408 561454 314728 561486
rect 314408 561218 314450 561454
rect 314686 561218 314728 561454
rect 314408 561134 314728 561218
rect 314408 560898 314450 561134
rect 314686 560898 314728 561134
rect 314408 560866 314728 560898
rect 345128 561454 345448 561486
rect 345128 561218 345170 561454
rect 345406 561218 345448 561454
rect 345128 561134 345448 561218
rect 345128 560898 345170 561134
rect 345406 560898 345448 561134
rect 345128 560866 345448 560898
rect 375848 561454 376168 561486
rect 375848 561218 375890 561454
rect 376126 561218 376168 561454
rect 375848 561134 376168 561218
rect 375848 560898 375890 561134
rect 376126 560898 376168 561134
rect 375848 560866 376168 560898
rect 406568 561454 406888 561486
rect 406568 561218 406610 561454
rect 406846 561218 406888 561454
rect 406568 561134 406888 561218
rect 406568 560898 406610 561134
rect 406846 560898 406888 561134
rect 406568 560866 406888 560898
rect 437288 561454 437608 561486
rect 437288 561218 437330 561454
rect 437566 561218 437608 561454
rect 437288 561134 437608 561218
rect 437288 560898 437330 561134
rect 437566 560898 437608 561134
rect 437288 560866 437608 560898
rect 468008 561454 468328 561486
rect 468008 561218 468050 561454
rect 468286 561218 468328 561454
rect 468008 561134 468328 561218
rect 468008 560898 468050 561134
rect 468286 560898 468328 561134
rect 468008 560866 468328 560898
rect 498728 561454 499048 561486
rect 498728 561218 498770 561454
rect 499006 561218 499048 561454
rect 498728 561134 499048 561218
rect 498728 560898 498770 561134
rect 499006 560898 499048 561134
rect 498728 560866 499048 560898
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 114728 543454 115048 543486
rect 114728 543218 114770 543454
rect 115006 543218 115048 543454
rect 114728 543134 115048 543218
rect 114728 542898 114770 543134
rect 115006 542898 115048 543134
rect 114728 542866 115048 542898
rect 145448 543454 145768 543486
rect 145448 543218 145490 543454
rect 145726 543218 145768 543454
rect 145448 543134 145768 543218
rect 145448 542898 145490 543134
rect 145726 542898 145768 543134
rect 145448 542866 145768 542898
rect 176168 543454 176488 543486
rect 176168 543218 176210 543454
rect 176446 543218 176488 543454
rect 176168 543134 176488 543218
rect 176168 542898 176210 543134
rect 176446 542898 176488 543134
rect 176168 542866 176488 542898
rect 206888 543454 207208 543486
rect 206888 543218 206930 543454
rect 207166 543218 207208 543454
rect 206888 543134 207208 543218
rect 206888 542898 206930 543134
rect 207166 542898 207208 543134
rect 206888 542866 207208 542898
rect 237608 543454 237928 543486
rect 237608 543218 237650 543454
rect 237886 543218 237928 543454
rect 237608 543134 237928 543218
rect 237608 542898 237650 543134
rect 237886 542898 237928 543134
rect 237608 542866 237928 542898
rect 268328 543454 268648 543486
rect 268328 543218 268370 543454
rect 268606 543218 268648 543454
rect 268328 543134 268648 543218
rect 268328 542898 268370 543134
rect 268606 542898 268648 543134
rect 268328 542866 268648 542898
rect 299048 543454 299368 543486
rect 299048 543218 299090 543454
rect 299326 543218 299368 543454
rect 299048 543134 299368 543218
rect 299048 542898 299090 543134
rect 299326 542898 299368 543134
rect 299048 542866 299368 542898
rect 329768 543454 330088 543486
rect 329768 543218 329810 543454
rect 330046 543218 330088 543454
rect 329768 543134 330088 543218
rect 329768 542898 329810 543134
rect 330046 542898 330088 543134
rect 329768 542866 330088 542898
rect 360488 543454 360808 543486
rect 360488 543218 360530 543454
rect 360766 543218 360808 543454
rect 360488 543134 360808 543218
rect 360488 542898 360530 543134
rect 360766 542898 360808 543134
rect 360488 542866 360808 542898
rect 391208 543454 391528 543486
rect 391208 543218 391250 543454
rect 391486 543218 391528 543454
rect 391208 543134 391528 543218
rect 391208 542898 391250 543134
rect 391486 542898 391528 543134
rect 391208 542866 391528 542898
rect 421928 543454 422248 543486
rect 421928 543218 421970 543454
rect 422206 543218 422248 543454
rect 421928 543134 422248 543218
rect 421928 542898 421970 543134
rect 422206 542898 422248 543134
rect 421928 542866 422248 542898
rect 452648 543454 452968 543486
rect 452648 543218 452690 543454
rect 452926 543218 452968 543454
rect 452648 543134 452968 543218
rect 452648 542898 452690 543134
rect 452926 542898 452968 543134
rect 452648 542866 452968 542898
rect 483368 543454 483688 543486
rect 483368 543218 483410 543454
rect 483646 543218 483688 543454
rect 483368 543134 483688 543218
rect 483368 542898 483410 543134
rect 483646 542898 483688 543134
rect 483368 542866 483688 542898
rect 99368 525454 99688 525486
rect 99368 525218 99410 525454
rect 99646 525218 99688 525454
rect 99368 525134 99688 525218
rect 99368 524898 99410 525134
rect 99646 524898 99688 525134
rect 99368 524866 99688 524898
rect 130088 525454 130408 525486
rect 130088 525218 130130 525454
rect 130366 525218 130408 525454
rect 130088 525134 130408 525218
rect 130088 524898 130130 525134
rect 130366 524898 130408 525134
rect 130088 524866 130408 524898
rect 160808 525454 161128 525486
rect 160808 525218 160850 525454
rect 161086 525218 161128 525454
rect 160808 525134 161128 525218
rect 160808 524898 160850 525134
rect 161086 524898 161128 525134
rect 160808 524866 161128 524898
rect 191528 525454 191848 525486
rect 191528 525218 191570 525454
rect 191806 525218 191848 525454
rect 191528 525134 191848 525218
rect 191528 524898 191570 525134
rect 191806 524898 191848 525134
rect 191528 524866 191848 524898
rect 222248 525454 222568 525486
rect 222248 525218 222290 525454
rect 222526 525218 222568 525454
rect 222248 525134 222568 525218
rect 222248 524898 222290 525134
rect 222526 524898 222568 525134
rect 222248 524866 222568 524898
rect 252968 525454 253288 525486
rect 252968 525218 253010 525454
rect 253246 525218 253288 525454
rect 252968 525134 253288 525218
rect 252968 524898 253010 525134
rect 253246 524898 253288 525134
rect 252968 524866 253288 524898
rect 283688 525454 284008 525486
rect 283688 525218 283730 525454
rect 283966 525218 284008 525454
rect 283688 525134 284008 525218
rect 283688 524898 283730 525134
rect 283966 524898 284008 525134
rect 283688 524866 284008 524898
rect 314408 525454 314728 525486
rect 314408 525218 314450 525454
rect 314686 525218 314728 525454
rect 314408 525134 314728 525218
rect 314408 524898 314450 525134
rect 314686 524898 314728 525134
rect 314408 524866 314728 524898
rect 345128 525454 345448 525486
rect 345128 525218 345170 525454
rect 345406 525218 345448 525454
rect 345128 525134 345448 525218
rect 345128 524898 345170 525134
rect 345406 524898 345448 525134
rect 345128 524866 345448 524898
rect 375848 525454 376168 525486
rect 375848 525218 375890 525454
rect 376126 525218 376168 525454
rect 375848 525134 376168 525218
rect 375848 524898 375890 525134
rect 376126 524898 376168 525134
rect 375848 524866 376168 524898
rect 406568 525454 406888 525486
rect 406568 525218 406610 525454
rect 406846 525218 406888 525454
rect 406568 525134 406888 525218
rect 406568 524898 406610 525134
rect 406846 524898 406888 525134
rect 406568 524866 406888 524898
rect 437288 525454 437608 525486
rect 437288 525218 437330 525454
rect 437566 525218 437608 525454
rect 437288 525134 437608 525218
rect 437288 524898 437330 525134
rect 437566 524898 437608 525134
rect 437288 524866 437608 524898
rect 468008 525454 468328 525486
rect 468008 525218 468050 525454
rect 468286 525218 468328 525454
rect 468008 525134 468328 525218
rect 468008 524898 468050 525134
rect 468286 524898 468328 525134
rect 468008 524866 468328 524898
rect 498728 525454 499048 525486
rect 498728 525218 498770 525454
rect 499006 525218 499048 525454
rect 498728 525134 499048 525218
rect 498728 524898 498770 525134
rect 499006 524898 499048 525134
rect 498728 524866 499048 524898
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 114728 507454 115048 507486
rect 114728 507218 114770 507454
rect 115006 507218 115048 507454
rect 114728 507134 115048 507218
rect 114728 506898 114770 507134
rect 115006 506898 115048 507134
rect 114728 506866 115048 506898
rect 145448 507454 145768 507486
rect 145448 507218 145490 507454
rect 145726 507218 145768 507454
rect 145448 507134 145768 507218
rect 145448 506898 145490 507134
rect 145726 506898 145768 507134
rect 145448 506866 145768 506898
rect 176168 507454 176488 507486
rect 176168 507218 176210 507454
rect 176446 507218 176488 507454
rect 176168 507134 176488 507218
rect 176168 506898 176210 507134
rect 176446 506898 176488 507134
rect 176168 506866 176488 506898
rect 206888 507454 207208 507486
rect 206888 507218 206930 507454
rect 207166 507218 207208 507454
rect 206888 507134 207208 507218
rect 206888 506898 206930 507134
rect 207166 506898 207208 507134
rect 206888 506866 207208 506898
rect 237608 507454 237928 507486
rect 237608 507218 237650 507454
rect 237886 507218 237928 507454
rect 237608 507134 237928 507218
rect 237608 506898 237650 507134
rect 237886 506898 237928 507134
rect 237608 506866 237928 506898
rect 268328 507454 268648 507486
rect 268328 507218 268370 507454
rect 268606 507218 268648 507454
rect 268328 507134 268648 507218
rect 268328 506898 268370 507134
rect 268606 506898 268648 507134
rect 268328 506866 268648 506898
rect 299048 507454 299368 507486
rect 299048 507218 299090 507454
rect 299326 507218 299368 507454
rect 299048 507134 299368 507218
rect 299048 506898 299090 507134
rect 299326 506898 299368 507134
rect 299048 506866 299368 506898
rect 329768 507454 330088 507486
rect 329768 507218 329810 507454
rect 330046 507218 330088 507454
rect 329768 507134 330088 507218
rect 329768 506898 329810 507134
rect 330046 506898 330088 507134
rect 329768 506866 330088 506898
rect 360488 507454 360808 507486
rect 360488 507218 360530 507454
rect 360766 507218 360808 507454
rect 360488 507134 360808 507218
rect 360488 506898 360530 507134
rect 360766 506898 360808 507134
rect 360488 506866 360808 506898
rect 391208 507454 391528 507486
rect 391208 507218 391250 507454
rect 391486 507218 391528 507454
rect 391208 507134 391528 507218
rect 391208 506898 391250 507134
rect 391486 506898 391528 507134
rect 391208 506866 391528 506898
rect 421928 507454 422248 507486
rect 421928 507218 421970 507454
rect 422206 507218 422248 507454
rect 421928 507134 422248 507218
rect 421928 506898 421970 507134
rect 422206 506898 422248 507134
rect 421928 506866 422248 506898
rect 452648 507454 452968 507486
rect 452648 507218 452690 507454
rect 452926 507218 452968 507454
rect 452648 507134 452968 507218
rect 452648 506898 452690 507134
rect 452926 506898 452968 507134
rect 452648 506866 452968 506898
rect 483368 507454 483688 507486
rect 483368 507218 483410 507454
rect 483646 507218 483688 507454
rect 483368 507134 483688 507218
rect 483368 506898 483410 507134
rect 483646 506898 483688 507134
rect 483368 506866 483688 506898
rect 99368 489454 99688 489486
rect 99368 489218 99410 489454
rect 99646 489218 99688 489454
rect 99368 489134 99688 489218
rect 99368 488898 99410 489134
rect 99646 488898 99688 489134
rect 99368 488866 99688 488898
rect 130088 489454 130408 489486
rect 130088 489218 130130 489454
rect 130366 489218 130408 489454
rect 130088 489134 130408 489218
rect 130088 488898 130130 489134
rect 130366 488898 130408 489134
rect 130088 488866 130408 488898
rect 160808 489454 161128 489486
rect 160808 489218 160850 489454
rect 161086 489218 161128 489454
rect 160808 489134 161128 489218
rect 160808 488898 160850 489134
rect 161086 488898 161128 489134
rect 160808 488866 161128 488898
rect 191528 489454 191848 489486
rect 191528 489218 191570 489454
rect 191806 489218 191848 489454
rect 191528 489134 191848 489218
rect 191528 488898 191570 489134
rect 191806 488898 191848 489134
rect 191528 488866 191848 488898
rect 222248 489454 222568 489486
rect 222248 489218 222290 489454
rect 222526 489218 222568 489454
rect 222248 489134 222568 489218
rect 222248 488898 222290 489134
rect 222526 488898 222568 489134
rect 222248 488866 222568 488898
rect 252968 489454 253288 489486
rect 252968 489218 253010 489454
rect 253246 489218 253288 489454
rect 252968 489134 253288 489218
rect 252968 488898 253010 489134
rect 253246 488898 253288 489134
rect 252968 488866 253288 488898
rect 283688 489454 284008 489486
rect 283688 489218 283730 489454
rect 283966 489218 284008 489454
rect 283688 489134 284008 489218
rect 283688 488898 283730 489134
rect 283966 488898 284008 489134
rect 283688 488866 284008 488898
rect 314408 489454 314728 489486
rect 314408 489218 314450 489454
rect 314686 489218 314728 489454
rect 314408 489134 314728 489218
rect 314408 488898 314450 489134
rect 314686 488898 314728 489134
rect 314408 488866 314728 488898
rect 345128 489454 345448 489486
rect 345128 489218 345170 489454
rect 345406 489218 345448 489454
rect 345128 489134 345448 489218
rect 345128 488898 345170 489134
rect 345406 488898 345448 489134
rect 345128 488866 345448 488898
rect 375848 489454 376168 489486
rect 375848 489218 375890 489454
rect 376126 489218 376168 489454
rect 375848 489134 376168 489218
rect 375848 488898 375890 489134
rect 376126 488898 376168 489134
rect 375848 488866 376168 488898
rect 406568 489454 406888 489486
rect 406568 489218 406610 489454
rect 406846 489218 406888 489454
rect 406568 489134 406888 489218
rect 406568 488898 406610 489134
rect 406846 488898 406888 489134
rect 406568 488866 406888 488898
rect 437288 489454 437608 489486
rect 437288 489218 437330 489454
rect 437566 489218 437608 489454
rect 437288 489134 437608 489218
rect 437288 488898 437330 489134
rect 437566 488898 437608 489134
rect 437288 488866 437608 488898
rect 468008 489454 468328 489486
rect 468008 489218 468050 489454
rect 468286 489218 468328 489454
rect 468008 489134 468328 489218
rect 468008 488898 468050 489134
rect 468286 488898 468328 489134
rect 468008 488866 468328 488898
rect 498728 489454 499048 489486
rect 498728 489218 498770 489454
rect 499006 489218 499048 489454
rect 498728 489134 499048 489218
rect 498728 488898 498770 489134
rect 499006 488898 499048 489134
rect 498728 488866 499048 488898
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 114728 471454 115048 471486
rect 114728 471218 114770 471454
rect 115006 471218 115048 471454
rect 114728 471134 115048 471218
rect 114728 470898 114770 471134
rect 115006 470898 115048 471134
rect 114728 470866 115048 470898
rect 145448 471454 145768 471486
rect 145448 471218 145490 471454
rect 145726 471218 145768 471454
rect 145448 471134 145768 471218
rect 145448 470898 145490 471134
rect 145726 470898 145768 471134
rect 145448 470866 145768 470898
rect 176168 471454 176488 471486
rect 176168 471218 176210 471454
rect 176446 471218 176488 471454
rect 176168 471134 176488 471218
rect 176168 470898 176210 471134
rect 176446 470898 176488 471134
rect 176168 470866 176488 470898
rect 206888 471454 207208 471486
rect 206888 471218 206930 471454
rect 207166 471218 207208 471454
rect 206888 471134 207208 471218
rect 206888 470898 206930 471134
rect 207166 470898 207208 471134
rect 206888 470866 207208 470898
rect 237608 471454 237928 471486
rect 237608 471218 237650 471454
rect 237886 471218 237928 471454
rect 237608 471134 237928 471218
rect 237608 470898 237650 471134
rect 237886 470898 237928 471134
rect 237608 470866 237928 470898
rect 268328 471454 268648 471486
rect 268328 471218 268370 471454
rect 268606 471218 268648 471454
rect 268328 471134 268648 471218
rect 268328 470898 268370 471134
rect 268606 470898 268648 471134
rect 268328 470866 268648 470898
rect 299048 471454 299368 471486
rect 299048 471218 299090 471454
rect 299326 471218 299368 471454
rect 299048 471134 299368 471218
rect 299048 470898 299090 471134
rect 299326 470898 299368 471134
rect 299048 470866 299368 470898
rect 329768 471454 330088 471486
rect 329768 471218 329810 471454
rect 330046 471218 330088 471454
rect 329768 471134 330088 471218
rect 329768 470898 329810 471134
rect 330046 470898 330088 471134
rect 329768 470866 330088 470898
rect 360488 471454 360808 471486
rect 360488 471218 360530 471454
rect 360766 471218 360808 471454
rect 360488 471134 360808 471218
rect 360488 470898 360530 471134
rect 360766 470898 360808 471134
rect 360488 470866 360808 470898
rect 391208 471454 391528 471486
rect 391208 471218 391250 471454
rect 391486 471218 391528 471454
rect 391208 471134 391528 471218
rect 391208 470898 391250 471134
rect 391486 470898 391528 471134
rect 391208 470866 391528 470898
rect 421928 471454 422248 471486
rect 421928 471218 421970 471454
rect 422206 471218 422248 471454
rect 421928 471134 422248 471218
rect 421928 470898 421970 471134
rect 422206 470898 422248 471134
rect 421928 470866 422248 470898
rect 452648 471454 452968 471486
rect 452648 471218 452690 471454
rect 452926 471218 452968 471454
rect 452648 471134 452968 471218
rect 452648 470898 452690 471134
rect 452926 470898 452968 471134
rect 452648 470866 452968 470898
rect 483368 471454 483688 471486
rect 483368 471218 483410 471454
rect 483646 471218 483688 471454
rect 483368 471134 483688 471218
rect 483368 470898 483410 471134
rect 483646 470898 483688 471134
rect 483368 470866 483688 470898
rect 99368 453454 99688 453486
rect 99368 453218 99410 453454
rect 99646 453218 99688 453454
rect 99368 453134 99688 453218
rect 99368 452898 99410 453134
rect 99646 452898 99688 453134
rect 99368 452866 99688 452898
rect 130088 453454 130408 453486
rect 130088 453218 130130 453454
rect 130366 453218 130408 453454
rect 130088 453134 130408 453218
rect 130088 452898 130130 453134
rect 130366 452898 130408 453134
rect 130088 452866 130408 452898
rect 160808 453454 161128 453486
rect 160808 453218 160850 453454
rect 161086 453218 161128 453454
rect 160808 453134 161128 453218
rect 160808 452898 160850 453134
rect 161086 452898 161128 453134
rect 160808 452866 161128 452898
rect 191528 453454 191848 453486
rect 191528 453218 191570 453454
rect 191806 453218 191848 453454
rect 191528 453134 191848 453218
rect 191528 452898 191570 453134
rect 191806 452898 191848 453134
rect 191528 452866 191848 452898
rect 222248 453454 222568 453486
rect 222248 453218 222290 453454
rect 222526 453218 222568 453454
rect 222248 453134 222568 453218
rect 222248 452898 222290 453134
rect 222526 452898 222568 453134
rect 222248 452866 222568 452898
rect 252968 453454 253288 453486
rect 252968 453218 253010 453454
rect 253246 453218 253288 453454
rect 252968 453134 253288 453218
rect 252968 452898 253010 453134
rect 253246 452898 253288 453134
rect 252968 452866 253288 452898
rect 283688 453454 284008 453486
rect 283688 453218 283730 453454
rect 283966 453218 284008 453454
rect 283688 453134 284008 453218
rect 283688 452898 283730 453134
rect 283966 452898 284008 453134
rect 283688 452866 284008 452898
rect 314408 453454 314728 453486
rect 314408 453218 314450 453454
rect 314686 453218 314728 453454
rect 314408 453134 314728 453218
rect 314408 452898 314450 453134
rect 314686 452898 314728 453134
rect 314408 452866 314728 452898
rect 345128 453454 345448 453486
rect 345128 453218 345170 453454
rect 345406 453218 345448 453454
rect 345128 453134 345448 453218
rect 345128 452898 345170 453134
rect 345406 452898 345448 453134
rect 345128 452866 345448 452898
rect 375848 453454 376168 453486
rect 375848 453218 375890 453454
rect 376126 453218 376168 453454
rect 375848 453134 376168 453218
rect 375848 452898 375890 453134
rect 376126 452898 376168 453134
rect 375848 452866 376168 452898
rect 406568 453454 406888 453486
rect 406568 453218 406610 453454
rect 406846 453218 406888 453454
rect 406568 453134 406888 453218
rect 406568 452898 406610 453134
rect 406846 452898 406888 453134
rect 406568 452866 406888 452898
rect 437288 453454 437608 453486
rect 437288 453218 437330 453454
rect 437566 453218 437608 453454
rect 437288 453134 437608 453218
rect 437288 452898 437330 453134
rect 437566 452898 437608 453134
rect 437288 452866 437608 452898
rect 468008 453454 468328 453486
rect 468008 453218 468050 453454
rect 468286 453218 468328 453454
rect 468008 453134 468328 453218
rect 468008 452898 468050 453134
rect 468286 452898 468328 453134
rect 468008 452866 468328 452898
rect 498728 453454 499048 453486
rect 498728 453218 498770 453454
rect 499006 453218 499048 453454
rect 498728 453134 499048 453218
rect 498728 452898 498770 453134
rect 499006 452898 499048 453134
rect 498728 452866 499048 452898
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 114728 435454 115048 435486
rect 114728 435218 114770 435454
rect 115006 435218 115048 435454
rect 114728 435134 115048 435218
rect 114728 434898 114770 435134
rect 115006 434898 115048 435134
rect 114728 434866 115048 434898
rect 145448 435454 145768 435486
rect 145448 435218 145490 435454
rect 145726 435218 145768 435454
rect 145448 435134 145768 435218
rect 145448 434898 145490 435134
rect 145726 434898 145768 435134
rect 145448 434866 145768 434898
rect 176168 435454 176488 435486
rect 176168 435218 176210 435454
rect 176446 435218 176488 435454
rect 176168 435134 176488 435218
rect 176168 434898 176210 435134
rect 176446 434898 176488 435134
rect 176168 434866 176488 434898
rect 206888 435454 207208 435486
rect 206888 435218 206930 435454
rect 207166 435218 207208 435454
rect 206888 435134 207208 435218
rect 206888 434898 206930 435134
rect 207166 434898 207208 435134
rect 206888 434866 207208 434898
rect 237608 435454 237928 435486
rect 237608 435218 237650 435454
rect 237886 435218 237928 435454
rect 237608 435134 237928 435218
rect 237608 434898 237650 435134
rect 237886 434898 237928 435134
rect 237608 434866 237928 434898
rect 268328 435454 268648 435486
rect 268328 435218 268370 435454
rect 268606 435218 268648 435454
rect 268328 435134 268648 435218
rect 268328 434898 268370 435134
rect 268606 434898 268648 435134
rect 268328 434866 268648 434898
rect 299048 435454 299368 435486
rect 299048 435218 299090 435454
rect 299326 435218 299368 435454
rect 299048 435134 299368 435218
rect 299048 434898 299090 435134
rect 299326 434898 299368 435134
rect 299048 434866 299368 434898
rect 329768 435454 330088 435486
rect 329768 435218 329810 435454
rect 330046 435218 330088 435454
rect 329768 435134 330088 435218
rect 329768 434898 329810 435134
rect 330046 434898 330088 435134
rect 329768 434866 330088 434898
rect 360488 435454 360808 435486
rect 360488 435218 360530 435454
rect 360766 435218 360808 435454
rect 360488 435134 360808 435218
rect 360488 434898 360530 435134
rect 360766 434898 360808 435134
rect 360488 434866 360808 434898
rect 391208 435454 391528 435486
rect 391208 435218 391250 435454
rect 391486 435218 391528 435454
rect 391208 435134 391528 435218
rect 391208 434898 391250 435134
rect 391486 434898 391528 435134
rect 391208 434866 391528 434898
rect 421928 435454 422248 435486
rect 421928 435218 421970 435454
rect 422206 435218 422248 435454
rect 421928 435134 422248 435218
rect 421928 434898 421970 435134
rect 422206 434898 422248 435134
rect 421928 434866 422248 434898
rect 452648 435454 452968 435486
rect 452648 435218 452690 435454
rect 452926 435218 452968 435454
rect 452648 435134 452968 435218
rect 452648 434898 452690 435134
rect 452926 434898 452968 435134
rect 452648 434866 452968 434898
rect 483368 435454 483688 435486
rect 483368 435218 483410 435454
rect 483646 435218 483688 435454
rect 483368 435134 483688 435218
rect 483368 434898 483410 435134
rect 483646 434898 483688 435134
rect 483368 434866 483688 434898
rect 99368 417454 99688 417486
rect 99368 417218 99410 417454
rect 99646 417218 99688 417454
rect 99368 417134 99688 417218
rect 99368 416898 99410 417134
rect 99646 416898 99688 417134
rect 99368 416866 99688 416898
rect 130088 417454 130408 417486
rect 130088 417218 130130 417454
rect 130366 417218 130408 417454
rect 130088 417134 130408 417218
rect 130088 416898 130130 417134
rect 130366 416898 130408 417134
rect 130088 416866 130408 416898
rect 160808 417454 161128 417486
rect 160808 417218 160850 417454
rect 161086 417218 161128 417454
rect 160808 417134 161128 417218
rect 160808 416898 160850 417134
rect 161086 416898 161128 417134
rect 160808 416866 161128 416898
rect 191528 417454 191848 417486
rect 191528 417218 191570 417454
rect 191806 417218 191848 417454
rect 191528 417134 191848 417218
rect 191528 416898 191570 417134
rect 191806 416898 191848 417134
rect 191528 416866 191848 416898
rect 222248 417454 222568 417486
rect 222248 417218 222290 417454
rect 222526 417218 222568 417454
rect 222248 417134 222568 417218
rect 222248 416898 222290 417134
rect 222526 416898 222568 417134
rect 222248 416866 222568 416898
rect 252968 417454 253288 417486
rect 252968 417218 253010 417454
rect 253246 417218 253288 417454
rect 252968 417134 253288 417218
rect 252968 416898 253010 417134
rect 253246 416898 253288 417134
rect 252968 416866 253288 416898
rect 283688 417454 284008 417486
rect 283688 417218 283730 417454
rect 283966 417218 284008 417454
rect 283688 417134 284008 417218
rect 283688 416898 283730 417134
rect 283966 416898 284008 417134
rect 283688 416866 284008 416898
rect 314408 417454 314728 417486
rect 314408 417218 314450 417454
rect 314686 417218 314728 417454
rect 314408 417134 314728 417218
rect 314408 416898 314450 417134
rect 314686 416898 314728 417134
rect 314408 416866 314728 416898
rect 345128 417454 345448 417486
rect 345128 417218 345170 417454
rect 345406 417218 345448 417454
rect 345128 417134 345448 417218
rect 345128 416898 345170 417134
rect 345406 416898 345448 417134
rect 345128 416866 345448 416898
rect 375848 417454 376168 417486
rect 375848 417218 375890 417454
rect 376126 417218 376168 417454
rect 375848 417134 376168 417218
rect 375848 416898 375890 417134
rect 376126 416898 376168 417134
rect 375848 416866 376168 416898
rect 406568 417454 406888 417486
rect 406568 417218 406610 417454
rect 406846 417218 406888 417454
rect 406568 417134 406888 417218
rect 406568 416898 406610 417134
rect 406846 416898 406888 417134
rect 406568 416866 406888 416898
rect 437288 417454 437608 417486
rect 437288 417218 437330 417454
rect 437566 417218 437608 417454
rect 437288 417134 437608 417218
rect 437288 416898 437330 417134
rect 437566 416898 437608 417134
rect 437288 416866 437608 416898
rect 468008 417454 468328 417486
rect 468008 417218 468050 417454
rect 468286 417218 468328 417454
rect 468008 417134 468328 417218
rect 468008 416898 468050 417134
rect 468286 416898 468328 417134
rect 468008 416866 468328 416898
rect 498728 417454 499048 417486
rect 498728 417218 498770 417454
rect 499006 417218 499048 417454
rect 498728 417134 499048 417218
rect 498728 416898 498770 417134
rect 499006 416898 499048 417134
rect 498728 416866 499048 416898
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 114728 399454 115048 399486
rect 114728 399218 114770 399454
rect 115006 399218 115048 399454
rect 114728 399134 115048 399218
rect 114728 398898 114770 399134
rect 115006 398898 115048 399134
rect 114728 398866 115048 398898
rect 145448 399454 145768 399486
rect 145448 399218 145490 399454
rect 145726 399218 145768 399454
rect 145448 399134 145768 399218
rect 145448 398898 145490 399134
rect 145726 398898 145768 399134
rect 145448 398866 145768 398898
rect 176168 399454 176488 399486
rect 176168 399218 176210 399454
rect 176446 399218 176488 399454
rect 176168 399134 176488 399218
rect 176168 398898 176210 399134
rect 176446 398898 176488 399134
rect 176168 398866 176488 398898
rect 206888 399454 207208 399486
rect 206888 399218 206930 399454
rect 207166 399218 207208 399454
rect 206888 399134 207208 399218
rect 206888 398898 206930 399134
rect 207166 398898 207208 399134
rect 206888 398866 207208 398898
rect 237608 399454 237928 399486
rect 237608 399218 237650 399454
rect 237886 399218 237928 399454
rect 237608 399134 237928 399218
rect 237608 398898 237650 399134
rect 237886 398898 237928 399134
rect 237608 398866 237928 398898
rect 268328 399454 268648 399486
rect 268328 399218 268370 399454
rect 268606 399218 268648 399454
rect 268328 399134 268648 399218
rect 268328 398898 268370 399134
rect 268606 398898 268648 399134
rect 268328 398866 268648 398898
rect 299048 399454 299368 399486
rect 299048 399218 299090 399454
rect 299326 399218 299368 399454
rect 299048 399134 299368 399218
rect 299048 398898 299090 399134
rect 299326 398898 299368 399134
rect 299048 398866 299368 398898
rect 329768 399454 330088 399486
rect 329768 399218 329810 399454
rect 330046 399218 330088 399454
rect 329768 399134 330088 399218
rect 329768 398898 329810 399134
rect 330046 398898 330088 399134
rect 329768 398866 330088 398898
rect 360488 399454 360808 399486
rect 360488 399218 360530 399454
rect 360766 399218 360808 399454
rect 360488 399134 360808 399218
rect 360488 398898 360530 399134
rect 360766 398898 360808 399134
rect 360488 398866 360808 398898
rect 391208 399454 391528 399486
rect 391208 399218 391250 399454
rect 391486 399218 391528 399454
rect 391208 399134 391528 399218
rect 391208 398898 391250 399134
rect 391486 398898 391528 399134
rect 391208 398866 391528 398898
rect 421928 399454 422248 399486
rect 421928 399218 421970 399454
rect 422206 399218 422248 399454
rect 421928 399134 422248 399218
rect 421928 398898 421970 399134
rect 422206 398898 422248 399134
rect 421928 398866 422248 398898
rect 452648 399454 452968 399486
rect 452648 399218 452690 399454
rect 452926 399218 452968 399454
rect 452648 399134 452968 399218
rect 452648 398898 452690 399134
rect 452926 398898 452968 399134
rect 452648 398866 452968 398898
rect 483368 399454 483688 399486
rect 483368 399218 483410 399454
rect 483646 399218 483688 399454
rect 483368 399134 483688 399218
rect 483368 398898 483410 399134
rect 483646 398898 483688 399134
rect 483368 398866 483688 398898
rect 99368 381454 99688 381486
rect 99368 381218 99410 381454
rect 99646 381218 99688 381454
rect 99368 381134 99688 381218
rect 99368 380898 99410 381134
rect 99646 380898 99688 381134
rect 99368 380866 99688 380898
rect 130088 381454 130408 381486
rect 130088 381218 130130 381454
rect 130366 381218 130408 381454
rect 130088 381134 130408 381218
rect 130088 380898 130130 381134
rect 130366 380898 130408 381134
rect 130088 380866 130408 380898
rect 160808 381454 161128 381486
rect 160808 381218 160850 381454
rect 161086 381218 161128 381454
rect 160808 381134 161128 381218
rect 160808 380898 160850 381134
rect 161086 380898 161128 381134
rect 160808 380866 161128 380898
rect 191528 381454 191848 381486
rect 191528 381218 191570 381454
rect 191806 381218 191848 381454
rect 191528 381134 191848 381218
rect 191528 380898 191570 381134
rect 191806 380898 191848 381134
rect 191528 380866 191848 380898
rect 222248 381454 222568 381486
rect 222248 381218 222290 381454
rect 222526 381218 222568 381454
rect 222248 381134 222568 381218
rect 222248 380898 222290 381134
rect 222526 380898 222568 381134
rect 222248 380866 222568 380898
rect 252968 381454 253288 381486
rect 252968 381218 253010 381454
rect 253246 381218 253288 381454
rect 252968 381134 253288 381218
rect 252968 380898 253010 381134
rect 253246 380898 253288 381134
rect 252968 380866 253288 380898
rect 283688 381454 284008 381486
rect 283688 381218 283730 381454
rect 283966 381218 284008 381454
rect 283688 381134 284008 381218
rect 283688 380898 283730 381134
rect 283966 380898 284008 381134
rect 283688 380866 284008 380898
rect 314408 381454 314728 381486
rect 314408 381218 314450 381454
rect 314686 381218 314728 381454
rect 314408 381134 314728 381218
rect 314408 380898 314450 381134
rect 314686 380898 314728 381134
rect 314408 380866 314728 380898
rect 345128 381454 345448 381486
rect 345128 381218 345170 381454
rect 345406 381218 345448 381454
rect 345128 381134 345448 381218
rect 345128 380898 345170 381134
rect 345406 380898 345448 381134
rect 345128 380866 345448 380898
rect 375848 381454 376168 381486
rect 375848 381218 375890 381454
rect 376126 381218 376168 381454
rect 375848 381134 376168 381218
rect 375848 380898 375890 381134
rect 376126 380898 376168 381134
rect 375848 380866 376168 380898
rect 406568 381454 406888 381486
rect 406568 381218 406610 381454
rect 406846 381218 406888 381454
rect 406568 381134 406888 381218
rect 406568 380898 406610 381134
rect 406846 380898 406888 381134
rect 406568 380866 406888 380898
rect 437288 381454 437608 381486
rect 437288 381218 437330 381454
rect 437566 381218 437608 381454
rect 437288 381134 437608 381218
rect 437288 380898 437330 381134
rect 437566 380898 437608 381134
rect 437288 380866 437608 380898
rect 468008 381454 468328 381486
rect 468008 381218 468050 381454
rect 468286 381218 468328 381454
rect 468008 381134 468328 381218
rect 468008 380898 468050 381134
rect 468286 380898 468328 381134
rect 468008 380866 468328 380898
rect 498728 381454 499048 381486
rect 498728 381218 498770 381454
rect 499006 381218 499048 381454
rect 498728 381134 499048 381218
rect 498728 380898 498770 381134
rect 499006 380898 499048 381134
rect 498728 380866 499048 380898
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 114728 363454 115048 363486
rect 114728 363218 114770 363454
rect 115006 363218 115048 363454
rect 114728 363134 115048 363218
rect 114728 362898 114770 363134
rect 115006 362898 115048 363134
rect 114728 362866 115048 362898
rect 145448 363454 145768 363486
rect 145448 363218 145490 363454
rect 145726 363218 145768 363454
rect 145448 363134 145768 363218
rect 145448 362898 145490 363134
rect 145726 362898 145768 363134
rect 145448 362866 145768 362898
rect 176168 363454 176488 363486
rect 176168 363218 176210 363454
rect 176446 363218 176488 363454
rect 176168 363134 176488 363218
rect 176168 362898 176210 363134
rect 176446 362898 176488 363134
rect 176168 362866 176488 362898
rect 206888 363454 207208 363486
rect 206888 363218 206930 363454
rect 207166 363218 207208 363454
rect 206888 363134 207208 363218
rect 206888 362898 206930 363134
rect 207166 362898 207208 363134
rect 206888 362866 207208 362898
rect 237608 363454 237928 363486
rect 237608 363218 237650 363454
rect 237886 363218 237928 363454
rect 237608 363134 237928 363218
rect 237608 362898 237650 363134
rect 237886 362898 237928 363134
rect 237608 362866 237928 362898
rect 268328 363454 268648 363486
rect 268328 363218 268370 363454
rect 268606 363218 268648 363454
rect 268328 363134 268648 363218
rect 268328 362898 268370 363134
rect 268606 362898 268648 363134
rect 268328 362866 268648 362898
rect 299048 363454 299368 363486
rect 299048 363218 299090 363454
rect 299326 363218 299368 363454
rect 299048 363134 299368 363218
rect 299048 362898 299090 363134
rect 299326 362898 299368 363134
rect 299048 362866 299368 362898
rect 329768 363454 330088 363486
rect 329768 363218 329810 363454
rect 330046 363218 330088 363454
rect 329768 363134 330088 363218
rect 329768 362898 329810 363134
rect 330046 362898 330088 363134
rect 329768 362866 330088 362898
rect 360488 363454 360808 363486
rect 360488 363218 360530 363454
rect 360766 363218 360808 363454
rect 360488 363134 360808 363218
rect 360488 362898 360530 363134
rect 360766 362898 360808 363134
rect 360488 362866 360808 362898
rect 391208 363454 391528 363486
rect 391208 363218 391250 363454
rect 391486 363218 391528 363454
rect 391208 363134 391528 363218
rect 391208 362898 391250 363134
rect 391486 362898 391528 363134
rect 391208 362866 391528 362898
rect 421928 363454 422248 363486
rect 421928 363218 421970 363454
rect 422206 363218 422248 363454
rect 421928 363134 422248 363218
rect 421928 362898 421970 363134
rect 422206 362898 422248 363134
rect 421928 362866 422248 362898
rect 452648 363454 452968 363486
rect 452648 363218 452690 363454
rect 452926 363218 452968 363454
rect 452648 363134 452968 363218
rect 452648 362898 452690 363134
rect 452926 362898 452968 363134
rect 452648 362866 452968 362898
rect 483368 363454 483688 363486
rect 483368 363218 483410 363454
rect 483646 363218 483688 363454
rect 483368 363134 483688 363218
rect 483368 362898 483410 363134
rect 483646 362898 483688 363134
rect 483368 362866 483688 362898
rect 99368 345454 99688 345486
rect 99368 345218 99410 345454
rect 99646 345218 99688 345454
rect 99368 345134 99688 345218
rect 99368 344898 99410 345134
rect 99646 344898 99688 345134
rect 99368 344866 99688 344898
rect 130088 345454 130408 345486
rect 130088 345218 130130 345454
rect 130366 345218 130408 345454
rect 130088 345134 130408 345218
rect 130088 344898 130130 345134
rect 130366 344898 130408 345134
rect 130088 344866 130408 344898
rect 160808 345454 161128 345486
rect 160808 345218 160850 345454
rect 161086 345218 161128 345454
rect 160808 345134 161128 345218
rect 160808 344898 160850 345134
rect 161086 344898 161128 345134
rect 160808 344866 161128 344898
rect 191528 345454 191848 345486
rect 191528 345218 191570 345454
rect 191806 345218 191848 345454
rect 191528 345134 191848 345218
rect 191528 344898 191570 345134
rect 191806 344898 191848 345134
rect 191528 344866 191848 344898
rect 222248 345454 222568 345486
rect 222248 345218 222290 345454
rect 222526 345218 222568 345454
rect 222248 345134 222568 345218
rect 222248 344898 222290 345134
rect 222526 344898 222568 345134
rect 222248 344866 222568 344898
rect 252968 345454 253288 345486
rect 252968 345218 253010 345454
rect 253246 345218 253288 345454
rect 252968 345134 253288 345218
rect 252968 344898 253010 345134
rect 253246 344898 253288 345134
rect 252968 344866 253288 344898
rect 283688 345454 284008 345486
rect 283688 345218 283730 345454
rect 283966 345218 284008 345454
rect 283688 345134 284008 345218
rect 283688 344898 283730 345134
rect 283966 344898 284008 345134
rect 283688 344866 284008 344898
rect 314408 345454 314728 345486
rect 314408 345218 314450 345454
rect 314686 345218 314728 345454
rect 314408 345134 314728 345218
rect 314408 344898 314450 345134
rect 314686 344898 314728 345134
rect 314408 344866 314728 344898
rect 345128 345454 345448 345486
rect 345128 345218 345170 345454
rect 345406 345218 345448 345454
rect 345128 345134 345448 345218
rect 345128 344898 345170 345134
rect 345406 344898 345448 345134
rect 345128 344866 345448 344898
rect 375848 345454 376168 345486
rect 375848 345218 375890 345454
rect 376126 345218 376168 345454
rect 375848 345134 376168 345218
rect 375848 344898 375890 345134
rect 376126 344898 376168 345134
rect 375848 344866 376168 344898
rect 406568 345454 406888 345486
rect 406568 345218 406610 345454
rect 406846 345218 406888 345454
rect 406568 345134 406888 345218
rect 406568 344898 406610 345134
rect 406846 344898 406888 345134
rect 406568 344866 406888 344898
rect 437288 345454 437608 345486
rect 437288 345218 437330 345454
rect 437566 345218 437608 345454
rect 437288 345134 437608 345218
rect 437288 344898 437330 345134
rect 437566 344898 437608 345134
rect 437288 344866 437608 344898
rect 468008 345454 468328 345486
rect 468008 345218 468050 345454
rect 468286 345218 468328 345454
rect 468008 345134 468328 345218
rect 468008 344898 468050 345134
rect 468286 344898 468328 345134
rect 468008 344866 468328 344898
rect 498728 345454 499048 345486
rect 498728 345218 498770 345454
rect 499006 345218 499048 345454
rect 498728 345134 499048 345218
rect 498728 344898 498770 345134
rect 499006 344898 499048 345134
rect 498728 344866 499048 344898
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 114728 327454 115048 327486
rect 114728 327218 114770 327454
rect 115006 327218 115048 327454
rect 114728 327134 115048 327218
rect 114728 326898 114770 327134
rect 115006 326898 115048 327134
rect 114728 326866 115048 326898
rect 145448 327454 145768 327486
rect 145448 327218 145490 327454
rect 145726 327218 145768 327454
rect 145448 327134 145768 327218
rect 145448 326898 145490 327134
rect 145726 326898 145768 327134
rect 145448 326866 145768 326898
rect 176168 327454 176488 327486
rect 176168 327218 176210 327454
rect 176446 327218 176488 327454
rect 176168 327134 176488 327218
rect 176168 326898 176210 327134
rect 176446 326898 176488 327134
rect 176168 326866 176488 326898
rect 206888 327454 207208 327486
rect 206888 327218 206930 327454
rect 207166 327218 207208 327454
rect 206888 327134 207208 327218
rect 206888 326898 206930 327134
rect 207166 326898 207208 327134
rect 206888 326866 207208 326898
rect 237608 327454 237928 327486
rect 237608 327218 237650 327454
rect 237886 327218 237928 327454
rect 237608 327134 237928 327218
rect 237608 326898 237650 327134
rect 237886 326898 237928 327134
rect 237608 326866 237928 326898
rect 268328 327454 268648 327486
rect 268328 327218 268370 327454
rect 268606 327218 268648 327454
rect 268328 327134 268648 327218
rect 268328 326898 268370 327134
rect 268606 326898 268648 327134
rect 268328 326866 268648 326898
rect 299048 327454 299368 327486
rect 299048 327218 299090 327454
rect 299326 327218 299368 327454
rect 299048 327134 299368 327218
rect 299048 326898 299090 327134
rect 299326 326898 299368 327134
rect 299048 326866 299368 326898
rect 329768 327454 330088 327486
rect 329768 327218 329810 327454
rect 330046 327218 330088 327454
rect 329768 327134 330088 327218
rect 329768 326898 329810 327134
rect 330046 326898 330088 327134
rect 329768 326866 330088 326898
rect 360488 327454 360808 327486
rect 360488 327218 360530 327454
rect 360766 327218 360808 327454
rect 360488 327134 360808 327218
rect 360488 326898 360530 327134
rect 360766 326898 360808 327134
rect 360488 326866 360808 326898
rect 391208 327454 391528 327486
rect 391208 327218 391250 327454
rect 391486 327218 391528 327454
rect 391208 327134 391528 327218
rect 391208 326898 391250 327134
rect 391486 326898 391528 327134
rect 391208 326866 391528 326898
rect 421928 327454 422248 327486
rect 421928 327218 421970 327454
rect 422206 327218 422248 327454
rect 421928 327134 422248 327218
rect 421928 326898 421970 327134
rect 422206 326898 422248 327134
rect 421928 326866 422248 326898
rect 452648 327454 452968 327486
rect 452648 327218 452690 327454
rect 452926 327218 452968 327454
rect 452648 327134 452968 327218
rect 452648 326898 452690 327134
rect 452926 326898 452968 327134
rect 452648 326866 452968 326898
rect 483368 327454 483688 327486
rect 483368 327218 483410 327454
rect 483646 327218 483688 327454
rect 483368 327134 483688 327218
rect 483368 326898 483410 327134
rect 483646 326898 483688 327134
rect 483368 326866 483688 326898
rect 99368 309454 99688 309486
rect 99368 309218 99410 309454
rect 99646 309218 99688 309454
rect 99368 309134 99688 309218
rect 99368 308898 99410 309134
rect 99646 308898 99688 309134
rect 99368 308866 99688 308898
rect 130088 309454 130408 309486
rect 130088 309218 130130 309454
rect 130366 309218 130408 309454
rect 130088 309134 130408 309218
rect 130088 308898 130130 309134
rect 130366 308898 130408 309134
rect 130088 308866 130408 308898
rect 160808 309454 161128 309486
rect 160808 309218 160850 309454
rect 161086 309218 161128 309454
rect 160808 309134 161128 309218
rect 160808 308898 160850 309134
rect 161086 308898 161128 309134
rect 160808 308866 161128 308898
rect 191528 309454 191848 309486
rect 191528 309218 191570 309454
rect 191806 309218 191848 309454
rect 191528 309134 191848 309218
rect 191528 308898 191570 309134
rect 191806 308898 191848 309134
rect 191528 308866 191848 308898
rect 222248 309454 222568 309486
rect 222248 309218 222290 309454
rect 222526 309218 222568 309454
rect 222248 309134 222568 309218
rect 222248 308898 222290 309134
rect 222526 308898 222568 309134
rect 222248 308866 222568 308898
rect 252968 309454 253288 309486
rect 252968 309218 253010 309454
rect 253246 309218 253288 309454
rect 252968 309134 253288 309218
rect 252968 308898 253010 309134
rect 253246 308898 253288 309134
rect 252968 308866 253288 308898
rect 283688 309454 284008 309486
rect 283688 309218 283730 309454
rect 283966 309218 284008 309454
rect 283688 309134 284008 309218
rect 283688 308898 283730 309134
rect 283966 308898 284008 309134
rect 283688 308866 284008 308898
rect 314408 309454 314728 309486
rect 314408 309218 314450 309454
rect 314686 309218 314728 309454
rect 314408 309134 314728 309218
rect 314408 308898 314450 309134
rect 314686 308898 314728 309134
rect 314408 308866 314728 308898
rect 345128 309454 345448 309486
rect 345128 309218 345170 309454
rect 345406 309218 345448 309454
rect 345128 309134 345448 309218
rect 345128 308898 345170 309134
rect 345406 308898 345448 309134
rect 345128 308866 345448 308898
rect 375848 309454 376168 309486
rect 375848 309218 375890 309454
rect 376126 309218 376168 309454
rect 375848 309134 376168 309218
rect 375848 308898 375890 309134
rect 376126 308898 376168 309134
rect 375848 308866 376168 308898
rect 406568 309454 406888 309486
rect 406568 309218 406610 309454
rect 406846 309218 406888 309454
rect 406568 309134 406888 309218
rect 406568 308898 406610 309134
rect 406846 308898 406888 309134
rect 406568 308866 406888 308898
rect 437288 309454 437608 309486
rect 437288 309218 437330 309454
rect 437566 309218 437608 309454
rect 437288 309134 437608 309218
rect 437288 308898 437330 309134
rect 437566 308898 437608 309134
rect 437288 308866 437608 308898
rect 468008 309454 468328 309486
rect 468008 309218 468050 309454
rect 468286 309218 468328 309454
rect 468008 309134 468328 309218
rect 468008 308898 468050 309134
rect 468286 308898 468328 309134
rect 468008 308866 468328 308898
rect 498728 309454 499048 309486
rect 498728 309218 498770 309454
rect 499006 309218 499048 309454
rect 498728 309134 499048 309218
rect 498728 308898 498770 309134
rect 499006 308898 499048 309134
rect 498728 308866 499048 308898
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 114728 291454 115048 291486
rect 114728 291218 114770 291454
rect 115006 291218 115048 291454
rect 114728 291134 115048 291218
rect 114728 290898 114770 291134
rect 115006 290898 115048 291134
rect 114728 290866 115048 290898
rect 145448 291454 145768 291486
rect 145448 291218 145490 291454
rect 145726 291218 145768 291454
rect 145448 291134 145768 291218
rect 145448 290898 145490 291134
rect 145726 290898 145768 291134
rect 145448 290866 145768 290898
rect 176168 291454 176488 291486
rect 176168 291218 176210 291454
rect 176446 291218 176488 291454
rect 176168 291134 176488 291218
rect 176168 290898 176210 291134
rect 176446 290898 176488 291134
rect 176168 290866 176488 290898
rect 206888 291454 207208 291486
rect 206888 291218 206930 291454
rect 207166 291218 207208 291454
rect 206888 291134 207208 291218
rect 206888 290898 206930 291134
rect 207166 290898 207208 291134
rect 206888 290866 207208 290898
rect 237608 291454 237928 291486
rect 237608 291218 237650 291454
rect 237886 291218 237928 291454
rect 237608 291134 237928 291218
rect 237608 290898 237650 291134
rect 237886 290898 237928 291134
rect 237608 290866 237928 290898
rect 268328 291454 268648 291486
rect 268328 291218 268370 291454
rect 268606 291218 268648 291454
rect 268328 291134 268648 291218
rect 268328 290898 268370 291134
rect 268606 290898 268648 291134
rect 268328 290866 268648 290898
rect 299048 291454 299368 291486
rect 299048 291218 299090 291454
rect 299326 291218 299368 291454
rect 299048 291134 299368 291218
rect 299048 290898 299090 291134
rect 299326 290898 299368 291134
rect 299048 290866 299368 290898
rect 329768 291454 330088 291486
rect 329768 291218 329810 291454
rect 330046 291218 330088 291454
rect 329768 291134 330088 291218
rect 329768 290898 329810 291134
rect 330046 290898 330088 291134
rect 329768 290866 330088 290898
rect 360488 291454 360808 291486
rect 360488 291218 360530 291454
rect 360766 291218 360808 291454
rect 360488 291134 360808 291218
rect 360488 290898 360530 291134
rect 360766 290898 360808 291134
rect 360488 290866 360808 290898
rect 391208 291454 391528 291486
rect 391208 291218 391250 291454
rect 391486 291218 391528 291454
rect 391208 291134 391528 291218
rect 391208 290898 391250 291134
rect 391486 290898 391528 291134
rect 391208 290866 391528 290898
rect 421928 291454 422248 291486
rect 421928 291218 421970 291454
rect 422206 291218 422248 291454
rect 421928 291134 422248 291218
rect 421928 290898 421970 291134
rect 422206 290898 422248 291134
rect 421928 290866 422248 290898
rect 452648 291454 452968 291486
rect 452648 291218 452690 291454
rect 452926 291218 452968 291454
rect 452648 291134 452968 291218
rect 452648 290898 452690 291134
rect 452926 290898 452968 291134
rect 452648 290866 452968 290898
rect 483368 291454 483688 291486
rect 483368 291218 483410 291454
rect 483646 291218 483688 291454
rect 483368 291134 483688 291218
rect 483368 290898 483410 291134
rect 483646 290898 483688 291134
rect 483368 290866 483688 290898
rect 99368 273454 99688 273486
rect 99368 273218 99410 273454
rect 99646 273218 99688 273454
rect 99368 273134 99688 273218
rect 99368 272898 99410 273134
rect 99646 272898 99688 273134
rect 99368 272866 99688 272898
rect 130088 273454 130408 273486
rect 130088 273218 130130 273454
rect 130366 273218 130408 273454
rect 130088 273134 130408 273218
rect 130088 272898 130130 273134
rect 130366 272898 130408 273134
rect 130088 272866 130408 272898
rect 160808 273454 161128 273486
rect 160808 273218 160850 273454
rect 161086 273218 161128 273454
rect 160808 273134 161128 273218
rect 160808 272898 160850 273134
rect 161086 272898 161128 273134
rect 160808 272866 161128 272898
rect 191528 273454 191848 273486
rect 191528 273218 191570 273454
rect 191806 273218 191848 273454
rect 191528 273134 191848 273218
rect 191528 272898 191570 273134
rect 191806 272898 191848 273134
rect 191528 272866 191848 272898
rect 222248 273454 222568 273486
rect 222248 273218 222290 273454
rect 222526 273218 222568 273454
rect 222248 273134 222568 273218
rect 222248 272898 222290 273134
rect 222526 272898 222568 273134
rect 222248 272866 222568 272898
rect 252968 273454 253288 273486
rect 252968 273218 253010 273454
rect 253246 273218 253288 273454
rect 252968 273134 253288 273218
rect 252968 272898 253010 273134
rect 253246 272898 253288 273134
rect 252968 272866 253288 272898
rect 283688 273454 284008 273486
rect 283688 273218 283730 273454
rect 283966 273218 284008 273454
rect 283688 273134 284008 273218
rect 283688 272898 283730 273134
rect 283966 272898 284008 273134
rect 283688 272866 284008 272898
rect 314408 273454 314728 273486
rect 314408 273218 314450 273454
rect 314686 273218 314728 273454
rect 314408 273134 314728 273218
rect 314408 272898 314450 273134
rect 314686 272898 314728 273134
rect 314408 272866 314728 272898
rect 345128 273454 345448 273486
rect 345128 273218 345170 273454
rect 345406 273218 345448 273454
rect 345128 273134 345448 273218
rect 345128 272898 345170 273134
rect 345406 272898 345448 273134
rect 345128 272866 345448 272898
rect 375848 273454 376168 273486
rect 375848 273218 375890 273454
rect 376126 273218 376168 273454
rect 375848 273134 376168 273218
rect 375848 272898 375890 273134
rect 376126 272898 376168 273134
rect 375848 272866 376168 272898
rect 406568 273454 406888 273486
rect 406568 273218 406610 273454
rect 406846 273218 406888 273454
rect 406568 273134 406888 273218
rect 406568 272898 406610 273134
rect 406846 272898 406888 273134
rect 406568 272866 406888 272898
rect 437288 273454 437608 273486
rect 437288 273218 437330 273454
rect 437566 273218 437608 273454
rect 437288 273134 437608 273218
rect 437288 272898 437330 273134
rect 437566 272898 437608 273134
rect 437288 272866 437608 272898
rect 468008 273454 468328 273486
rect 468008 273218 468050 273454
rect 468286 273218 468328 273454
rect 468008 273134 468328 273218
rect 468008 272898 468050 273134
rect 468286 272898 468328 273134
rect 468008 272866 468328 272898
rect 498728 273454 499048 273486
rect 498728 273218 498770 273454
rect 499006 273218 499048 273454
rect 498728 273134 499048 273218
rect 498728 272898 498770 273134
rect 499006 272898 499048 273134
rect 498728 272866 499048 272898
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 114728 255454 115048 255486
rect 114728 255218 114770 255454
rect 115006 255218 115048 255454
rect 114728 255134 115048 255218
rect 114728 254898 114770 255134
rect 115006 254898 115048 255134
rect 114728 254866 115048 254898
rect 145448 255454 145768 255486
rect 145448 255218 145490 255454
rect 145726 255218 145768 255454
rect 145448 255134 145768 255218
rect 145448 254898 145490 255134
rect 145726 254898 145768 255134
rect 145448 254866 145768 254898
rect 176168 255454 176488 255486
rect 176168 255218 176210 255454
rect 176446 255218 176488 255454
rect 176168 255134 176488 255218
rect 176168 254898 176210 255134
rect 176446 254898 176488 255134
rect 176168 254866 176488 254898
rect 206888 255454 207208 255486
rect 206888 255218 206930 255454
rect 207166 255218 207208 255454
rect 206888 255134 207208 255218
rect 206888 254898 206930 255134
rect 207166 254898 207208 255134
rect 206888 254866 207208 254898
rect 237608 255454 237928 255486
rect 237608 255218 237650 255454
rect 237886 255218 237928 255454
rect 237608 255134 237928 255218
rect 237608 254898 237650 255134
rect 237886 254898 237928 255134
rect 237608 254866 237928 254898
rect 268328 255454 268648 255486
rect 268328 255218 268370 255454
rect 268606 255218 268648 255454
rect 268328 255134 268648 255218
rect 268328 254898 268370 255134
rect 268606 254898 268648 255134
rect 268328 254866 268648 254898
rect 299048 255454 299368 255486
rect 299048 255218 299090 255454
rect 299326 255218 299368 255454
rect 299048 255134 299368 255218
rect 299048 254898 299090 255134
rect 299326 254898 299368 255134
rect 299048 254866 299368 254898
rect 329768 255454 330088 255486
rect 329768 255218 329810 255454
rect 330046 255218 330088 255454
rect 329768 255134 330088 255218
rect 329768 254898 329810 255134
rect 330046 254898 330088 255134
rect 329768 254866 330088 254898
rect 360488 255454 360808 255486
rect 360488 255218 360530 255454
rect 360766 255218 360808 255454
rect 360488 255134 360808 255218
rect 360488 254898 360530 255134
rect 360766 254898 360808 255134
rect 360488 254866 360808 254898
rect 391208 255454 391528 255486
rect 391208 255218 391250 255454
rect 391486 255218 391528 255454
rect 391208 255134 391528 255218
rect 391208 254898 391250 255134
rect 391486 254898 391528 255134
rect 391208 254866 391528 254898
rect 421928 255454 422248 255486
rect 421928 255218 421970 255454
rect 422206 255218 422248 255454
rect 421928 255134 422248 255218
rect 421928 254898 421970 255134
rect 422206 254898 422248 255134
rect 421928 254866 422248 254898
rect 452648 255454 452968 255486
rect 452648 255218 452690 255454
rect 452926 255218 452968 255454
rect 452648 255134 452968 255218
rect 452648 254898 452690 255134
rect 452926 254898 452968 255134
rect 452648 254866 452968 254898
rect 483368 255454 483688 255486
rect 483368 255218 483410 255454
rect 483646 255218 483688 255454
rect 483368 255134 483688 255218
rect 483368 254898 483410 255134
rect 483646 254898 483688 255134
rect 483368 254866 483688 254898
rect 99368 237454 99688 237486
rect 99368 237218 99410 237454
rect 99646 237218 99688 237454
rect 99368 237134 99688 237218
rect 99368 236898 99410 237134
rect 99646 236898 99688 237134
rect 99368 236866 99688 236898
rect 130088 237454 130408 237486
rect 130088 237218 130130 237454
rect 130366 237218 130408 237454
rect 130088 237134 130408 237218
rect 130088 236898 130130 237134
rect 130366 236898 130408 237134
rect 130088 236866 130408 236898
rect 160808 237454 161128 237486
rect 160808 237218 160850 237454
rect 161086 237218 161128 237454
rect 160808 237134 161128 237218
rect 160808 236898 160850 237134
rect 161086 236898 161128 237134
rect 160808 236866 161128 236898
rect 191528 237454 191848 237486
rect 191528 237218 191570 237454
rect 191806 237218 191848 237454
rect 191528 237134 191848 237218
rect 191528 236898 191570 237134
rect 191806 236898 191848 237134
rect 191528 236866 191848 236898
rect 222248 237454 222568 237486
rect 222248 237218 222290 237454
rect 222526 237218 222568 237454
rect 222248 237134 222568 237218
rect 222248 236898 222290 237134
rect 222526 236898 222568 237134
rect 222248 236866 222568 236898
rect 252968 237454 253288 237486
rect 252968 237218 253010 237454
rect 253246 237218 253288 237454
rect 252968 237134 253288 237218
rect 252968 236898 253010 237134
rect 253246 236898 253288 237134
rect 252968 236866 253288 236898
rect 283688 237454 284008 237486
rect 283688 237218 283730 237454
rect 283966 237218 284008 237454
rect 283688 237134 284008 237218
rect 283688 236898 283730 237134
rect 283966 236898 284008 237134
rect 283688 236866 284008 236898
rect 314408 237454 314728 237486
rect 314408 237218 314450 237454
rect 314686 237218 314728 237454
rect 314408 237134 314728 237218
rect 314408 236898 314450 237134
rect 314686 236898 314728 237134
rect 314408 236866 314728 236898
rect 345128 237454 345448 237486
rect 345128 237218 345170 237454
rect 345406 237218 345448 237454
rect 345128 237134 345448 237218
rect 345128 236898 345170 237134
rect 345406 236898 345448 237134
rect 345128 236866 345448 236898
rect 375848 237454 376168 237486
rect 375848 237218 375890 237454
rect 376126 237218 376168 237454
rect 375848 237134 376168 237218
rect 375848 236898 375890 237134
rect 376126 236898 376168 237134
rect 375848 236866 376168 236898
rect 406568 237454 406888 237486
rect 406568 237218 406610 237454
rect 406846 237218 406888 237454
rect 406568 237134 406888 237218
rect 406568 236898 406610 237134
rect 406846 236898 406888 237134
rect 406568 236866 406888 236898
rect 437288 237454 437608 237486
rect 437288 237218 437330 237454
rect 437566 237218 437608 237454
rect 437288 237134 437608 237218
rect 437288 236898 437330 237134
rect 437566 236898 437608 237134
rect 437288 236866 437608 236898
rect 468008 237454 468328 237486
rect 468008 237218 468050 237454
rect 468286 237218 468328 237454
rect 468008 237134 468328 237218
rect 468008 236898 468050 237134
rect 468286 236898 468328 237134
rect 468008 236866 468328 236898
rect 498728 237454 499048 237486
rect 498728 237218 498770 237454
rect 499006 237218 499048 237454
rect 498728 237134 499048 237218
rect 498728 236898 498770 237134
rect 499006 236898 499048 237134
rect 498728 236866 499048 236898
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 114728 219454 115048 219486
rect 114728 219218 114770 219454
rect 115006 219218 115048 219454
rect 114728 219134 115048 219218
rect 114728 218898 114770 219134
rect 115006 218898 115048 219134
rect 114728 218866 115048 218898
rect 145448 219454 145768 219486
rect 145448 219218 145490 219454
rect 145726 219218 145768 219454
rect 145448 219134 145768 219218
rect 145448 218898 145490 219134
rect 145726 218898 145768 219134
rect 145448 218866 145768 218898
rect 176168 219454 176488 219486
rect 176168 219218 176210 219454
rect 176446 219218 176488 219454
rect 176168 219134 176488 219218
rect 176168 218898 176210 219134
rect 176446 218898 176488 219134
rect 176168 218866 176488 218898
rect 206888 219454 207208 219486
rect 206888 219218 206930 219454
rect 207166 219218 207208 219454
rect 206888 219134 207208 219218
rect 206888 218898 206930 219134
rect 207166 218898 207208 219134
rect 206888 218866 207208 218898
rect 237608 219454 237928 219486
rect 237608 219218 237650 219454
rect 237886 219218 237928 219454
rect 237608 219134 237928 219218
rect 237608 218898 237650 219134
rect 237886 218898 237928 219134
rect 237608 218866 237928 218898
rect 268328 219454 268648 219486
rect 268328 219218 268370 219454
rect 268606 219218 268648 219454
rect 268328 219134 268648 219218
rect 268328 218898 268370 219134
rect 268606 218898 268648 219134
rect 268328 218866 268648 218898
rect 299048 219454 299368 219486
rect 299048 219218 299090 219454
rect 299326 219218 299368 219454
rect 299048 219134 299368 219218
rect 299048 218898 299090 219134
rect 299326 218898 299368 219134
rect 299048 218866 299368 218898
rect 329768 219454 330088 219486
rect 329768 219218 329810 219454
rect 330046 219218 330088 219454
rect 329768 219134 330088 219218
rect 329768 218898 329810 219134
rect 330046 218898 330088 219134
rect 329768 218866 330088 218898
rect 360488 219454 360808 219486
rect 360488 219218 360530 219454
rect 360766 219218 360808 219454
rect 360488 219134 360808 219218
rect 360488 218898 360530 219134
rect 360766 218898 360808 219134
rect 360488 218866 360808 218898
rect 391208 219454 391528 219486
rect 391208 219218 391250 219454
rect 391486 219218 391528 219454
rect 391208 219134 391528 219218
rect 391208 218898 391250 219134
rect 391486 218898 391528 219134
rect 391208 218866 391528 218898
rect 421928 219454 422248 219486
rect 421928 219218 421970 219454
rect 422206 219218 422248 219454
rect 421928 219134 422248 219218
rect 421928 218898 421970 219134
rect 422206 218898 422248 219134
rect 421928 218866 422248 218898
rect 452648 219454 452968 219486
rect 452648 219218 452690 219454
rect 452926 219218 452968 219454
rect 452648 219134 452968 219218
rect 452648 218898 452690 219134
rect 452926 218898 452968 219134
rect 452648 218866 452968 218898
rect 483368 219454 483688 219486
rect 483368 219218 483410 219454
rect 483646 219218 483688 219454
rect 483368 219134 483688 219218
rect 483368 218898 483410 219134
rect 483646 218898 483688 219134
rect 483368 218866 483688 218898
rect 99368 201454 99688 201486
rect 99368 201218 99410 201454
rect 99646 201218 99688 201454
rect 99368 201134 99688 201218
rect 99368 200898 99410 201134
rect 99646 200898 99688 201134
rect 99368 200866 99688 200898
rect 130088 201454 130408 201486
rect 130088 201218 130130 201454
rect 130366 201218 130408 201454
rect 130088 201134 130408 201218
rect 130088 200898 130130 201134
rect 130366 200898 130408 201134
rect 130088 200866 130408 200898
rect 160808 201454 161128 201486
rect 160808 201218 160850 201454
rect 161086 201218 161128 201454
rect 160808 201134 161128 201218
rect 160808 200898 160850 201134
rect 161086 200898 161128 201134
rect 160808 200866 161128 200898
rect 191528 201454 191848 201486
rect 191528 201218 191570 201454
rect 191806 201218 191848 201454
rect 191528 201134 191848 201218
rect 191528 200898 191570 201134
rect 191806 200898 191848 201134
rect 191528 200866 191848 200898
rect 222248 201454 222568 201486
rect 222248 201218 222290 201454
rect 222526 201218 222568 201454
rect 222248 201134 222568 201218
rect 222248 200898 222290 201134
rect 222526 200898 222568 201134
rect 222248 200866 222568 200898
rect 252968 201454 253288 201486
rect 252968 201218 253010 201454
rect 253246 201218 253288 201454
rect 252968 201134 253288 201218
rect 252968 200898 253010 201134
rect 253246 200898 253288 201134
rect 252968 200866 253288 200898
rect 283688 201454 284008 201486
rect 283688 201218 283730 201454
rect 283966 201218 284008 201454
rect 283688 201134 284008 201218
rect 283688 200898 283730 201134
rect 283966 200898 284008 201134
rect 283688 200866 284008 200898
rect 314408 201454 314728 201486
rect 314408 201218 314450 201454
rect 314686 201218 314728 201454
rect 314408 201134 314728 201218
rect 314408 200898 314450 201134
rect 314686 200898 314728 201134
rect 314408 200866 314728 200898
rect 345128 201454 345448 201486
rect 345128 201218 345170 201454
rect 345406 201218 345448 201454
rect 345128 201134 345448 201218
rect 345128 200898 345170 201134
rect 345406 200898 345448 201134
rect 345128 200866 345448 200898
rect 375848 201454 376168 201486
rect 375848 201218 375890 201454
rect 376126 201218 376168 201454
rect 375848 201134 376168 201218
rect 375848 200898 375890 201134
rect 376126 200898 376168 201134
rect 375848 200866 376168 200898
rect 406568 201454 406888 201486
rect 406568 201218 406610 201454
rect 406846 201218 406888 201454
rect 406568 201134 406888 201218
rect 406568 200898 406610 201134
rect 406846 200898 406888 201134
rect 406568 200866 406888 200898
rect 437288 201454 437608 201486
rect 437288 201218 437330 201454
rect 437566 201218 437608 201454
rect 437288 201134 437608 201218
rect 437288 200898 437330 201134
rect 437566 200898 437608 201134
rect 437288 200866 437608 200898
rect 468008 201454 468328 201486
rect 468008 201218 468050 201454
rect 468286 201218 468328 201454
rect 468008 201134 468328 201218
rect 468008 200898 468050 201134
rect 468286 200898 468328 201134
rect 468008 200866 468328 200898
rect 498728 201454 499048 201486
rect 498728 201218 498770 201454
rect 499006 201218 499048 201454
rect 498728 201134 499048 201218
rect 498728 200898 498770 201134
rect 499006 200898 499048 201134
rect 498728 200866 499048 200898
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 114728 183454 115048 183486
rect 114728 183218 114770 183454
rect 115006 183218 115048 183454
rect 114728 183134 115048 183218
rect 114728 182898 114770 183134
rect 115006 182898 115048 183134
rect 114728 182866 115048 182898
rect 145448 183454 145768 183486
rect 145448 183218 145490 183454
rect 145726 183218 145768 183454
rect 145448 183134 145768 183218
rect 145448 182898 145490 183134
rect 145726 182898 145768 183134
rect 145448 182866 145768 182898
rect 176168 183454 176488 183486
rect 176168 183218 176210 183454
rect 176446 183218 176488 183454
rect 176168 183134 176488 183218
rect 176168 182898 176210 183134
rect 176446 182898 176488 183134
rect 176168 182866 176488 182898
rect 206888 183454 207208 183486
rect 206888 183218 206930 183454
rect 207166 183218 207208 183454
rect 206888 183134 207208 183218
rect 206888 182898 206930 183134
rect 207166 182898 207208 183134
rect 206888 182866 207208 182898
rect 237608 183454 237928 183486
rect 237608 183218 237650 183454
rect 237886 183218 237928 183454
rect 237608 183134 237928 183218
rect 237608 182898 237650 183134
rect 237886 182898 237928 183134
rect 237608 182866 237928 182898
rect 268328 183454 268648 183486
rect 268328 183218 268370 183454
rect 268606 183218 268648 183454
rect 268328 183134 268648 183218
rect 268328 182898 268370 183134
rect 268606 182898 268648 183134
rect 268328 182866 268648 182898
rect 299048 183454 299368 183486
rect 299048 183218 299090 183454
rect 299326 183218 299368 183454
rect 299048 183134 299368 183218
rect 299048 182898 299090 183134
rect 299326 182898 299368 183134
rect 299048 182866 299368 182898
rect 329768 183454 330088 183486
rect 329768 183218 329810 183454
rect 330046 183218 330088 183454
rect 329768 183134 330088 183218
rect 329768 182898 329810 183134
rect 330046 182898 330088 183134
rect 329768 182866 330088 182898
rect 360488 183454 360808 183486
rect 360488 183218 360530 183454
rect 360766 183218 360808 183454
rect 360488 183134 360808 183218
rect 360488 182898 360530 183134
rect 360766 182898 360808 183134
rect 360488 182866 360808 182898
rect 391208 183454 391528 183486
rect 391208 183218 391250 183454
rect 391486 183218 391528 183454
rect 391208 183134 391528 183218
rect 391208 182898 391250 183134
rect 391486 182898 391528 183134
rect 391208 182866 391528 182898
rect 421928 183454 422248 183486
rect 421928 183218 421970 183454
rect 422206 183218 422248 183454
rect 421928 183134 422248 183218
rect 421928 182898 421970 183134
rect 422206 182898 422248 183134
rect 421928 182866 422248 182898
rect 452648 183454 452968 183486
rect 452648 183218 452690 183454
rect 452926 183218 452968 183454
rect 452648 183134 452968 183218
rect 452648 182898 452690 183134
rect 452926 182898 452968 183134
rect 452648 182866 452968 182898
rect 483368 183454 483688 183486
rect 483368 183218 483410 183454
rect 483646 183218 483688 183454
rect 483368 183134 483688 183218
rect 483368 182898 483410 183134
rect 483646 182898 483688 183134
rect 483368 182866 483688 182898
rect 99368 165454 99688 165486
rect 99368 165218 99410 165454
rect 99646 165218 99688 165454
rect 99368 165134 99688 165218
rect 99368 164898 99410 165134
rect 99646 164898 99688 165134
rect 99368 164866 99688 164898
rect 130088 165454 130408 165486
rect 130088 165218 130130 165454
rect 130366 165218 130408 165454
rect 130088 165134 130408 165218
rect 130088 164898 130130 165134
rect 130366 164898 130408 165134
rect 130088 164866 130408 164898
rect 160808 165454 161128 165486
rect 160808 165218 160850 165454
rect 161086 165218 161128 165454
rect 160808 165134 161128 165218
rect 160808 164898 160850 165134
rect 161086 164898 161128 165134
rect 160808 164866 161128 164898
rect 191528 165454 191848 165486
rect 191528 165218 191570 165454
rect 191806 165218 191848 165454
rect 191528 165134 191848 165218
rect 191528 164898 191570 165134
rect 191806 164898 191848 165134
rect 191528 164866 191848 164898
rect 222248 165454 222568 165486
rect 222248 165218 222290 165454
rect 222526 165218 222568 165454
rect 222248 165134 222568 165218
rect 222248 164898 222290 165134
rect 222526 164898 222568 165134
rect 222248 164866 222568 164898
rect 252968 165454 253288 165486
rect 252968 165218 253010 165454
rect 253246 165218 253288 165454
rect 252968 165134 253288 165218
rect 252968 164898 253010 165134
rect 253246 164898 253288 165134
rect 252968 164866 253288 164898
rect 283688 165454 284008 165486
rect 283688 165218 283730 165454
rect 283966 165218 284008 165454
rect 283688 165134 284008 165218
rect 283688 164898 283730 165134
rect 283966 164898 284008 165134
rect 283688 164866 284008 164898
rect 314408 165454 314728 165486
rect 314408 165218 314450 165454
rect 314686 165218 314728 165454
rect 314408 165134 314728 165218
rect 314408 164898 314450 165134
rect 314686 164898 314728 165134
rect 314408 164866 314728 164898
rect 345128 165454 345448 165486
rect 345128 165218 345170 165454
rect 345406 165218 345448 165454
rect 345128 165134 345448 165218
rect 345128 164898 345170 165134
rect 345406 164898 345448 165134
rect 345128 164866 345448 164898
rect 375848 165454 376168 165486
rect 375848 165218 375890 165454
rect 376126 165218 376168 165454
rect 375848 165134 376168 165218
rect 375848 164898 375890 165134
rect 376126 164898 376168 165134
rect 375848 164866 376168 164898
rect 406568 165454 406888 165486
rect 406568 165218 406610 165454
rect 406846 165218 406888 165454
rect 406568 165134 406888 165218
rect 406568 164898 406610 165134
rect 406846 164898 406888 165134
rect 406568 164866 406888 164898
rect 437288 165454 437608 165486
rect 437288 165218 437330 165454
rect 437566 165218 437608 165454
rect 437288 165134 437608 165218
rect 437288 164898 437330 165134
rect 437566 164898 437608 165134
rect 437288 164866 437608 164898
rect 468008 165454 468328 165486
rect 468008 165218 468050 165454
rect 468286 165218 468328 165454
rect 468008 165134 468328 165218
rect 468008 164898 468050 165134
rect 468286 164898 468328 165134
rect 468008 164866 468328 164898
rect 498728 165454 499048 165486
rect 498728 165218 498770 165454
rect 499006 165218 499048 165454
rect 498728 165134 499048 165218
rect 498728 164898 498770 165134
rect 499006 164898 499048 165134
rect 498728 164866 499048 164898
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 114728 147454 115048 147486
rect 114728 147218 114770 147454
rect 115006 147218 115048 147454
rect 114728 147134 115048 147218
rect 114728 146898 114770 147134
rect 115006 146898 115048 147134
rect 114728 146866 115048 146898
rect 145448 147454 145768 147486
rect 145448 147218 145490 147454
rect 145726 147218 145768 147454
rect 145448 147134 145768 147218
rect 145448 146898 145490 147134
rect 145726 146898 145768 147134
rect 145448 146866 145768 146898
rect 176168 147454 176488 147486
rect 176168 147218 176210 147454
rect 176446 147218 176488 147454
rect 176168 147134 176488 147218
rect 176168 146898 176210 147134
rect 176446 146898 176488 147134
rect 176168 146866 176488 146898
rect 206888 147454 207208 147486
rect 206888 147218 206930 147454
rect 207166 147218 207208 147454
rect 206888 147134 207208 147218
rect 206888 146898 206930 147134
rect 207166 146898 207208 147134
rect 206888 146866 207208 146898
rect 237608 147454 237928 147486
rect 237608 147218 237650 147454
rect 237886 147218 237928 147454
rect 237608 147134 237928 147218
rect 237608 146898 237650 147134
rect 237886 146898 237928 147134
rect 237608 146866 237928 146898
rect 268328 147454 268648 147486
rect 268328 147218 268370 147454
rect 268606 147218 268648 147454
rect 268328 147134 268648 147218
rect 268328 146898 268370 147134
rect 268606 146898 268648 147134
rect 268328 146866 268648 146898
rect 299048 147454 299368 147486
rect 299048 147218 299090 147454
rect 299326 147218 299368 147454
rect 299048 147134 299368 147218
rect 299048 146898 299090 147134
rect 299326 146898 299368 147134
rect 299048 146866 299368 146898
rect 329768 147454 330088 147486
rect 329768 147218 329810 147454
rect 330046 147218 330088 147454
rect 329768 147134 330088 147218
rect 329768 146898 329810 147134
rect 330046 146898 330088 147134
rect 329768 146866 330088 146898
rect 360488 147454 360808 147486
rect 360488 147218 360530 147454
rect 360766 147218 360808 147454
rect 360488 147134 360808 147218
rect 360488 146898 360530 147134
rect 360766 146898 360808 147134
rect 360488 146866 360808 146898
rect 391208 147454 391528 147486
rect 391208 147218 391250 147454
rect 391486 147218 391528 147454
rect 391208 147134 391528 147218
rect 391208 146898 391250 147134
rect 391486 146898 391528 147134
rect 391208 146866 391528 146898
rect 421928 147454 422248 147486
rect 421928 147218 421970 147454
rect 422206 147218 422248 147454
rect 421928 147134 422248 147218
rect 421928 146898 421970 147134
rect 422206 146898 422248 147134
rect 421928 146866 422248 146898
rect 452648 147454 452968 147486
rect 452648 147218 452690 147454
rect 452926 147218 452968 147454
rect 452648 147134 452968 147218
rect 452648 146898 452690 147134
rect 452926 146898 452968 147134
rect 452648 146866 452968 146898
rect 483368 147454 483688 147486
rect 483368 147218 483410 147454
rect 483646 147218 483688 147454
rect 483368 147134 483688 147218
rect 483368 146898 483410 147134
rect 483646 146898 483688 147134
rect 483368 146866 483688 146898
rect 99234 100894 99854 136600
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 96475 71908 96541 71909
rect 96475 71844 96476 71908
rect 96540 71844 96541 71908
rect 96475 71843 96541 71844
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 93715 45660 93781 45661
rect 93715 45596 93716 45660
rect 93780 45596 93781 45660
rect 93715 45595 93781 45596
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 89483 19412 89549 19413
rect 89483 19348 89484 19412
rect 89548 19348 89549 19412
rect 89483 19347 89549 19348
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 82675 5676 82741 5677
rect 82675 5612 82676 5676
rect 82740 5612 82741 5676
rect 82675 5611 82741 5612
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 104614 103574 136600
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 111454 110414 136600
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 115174 114134 136600
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 118894 117854 136600
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 122614 121574 136600
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 129454 128414 136600
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 133174 132134 136600
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 100894 135854 136600
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 104614 139574 136600
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 111454 146414 136600
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 115174 150134 136600
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 118894 153854 136600
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 122614 157574 136600
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 129454 164414 136600
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 133174 168134 136600
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 100894 171854 136600
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 104614 175574 136600
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 111454 182414 136600
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 115174 186134 136600
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 118894 189854 136600
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 122614 193574 136600
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 129454 200414 136600
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 133174 204134 136600
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 100894 207854 136600
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 104614 211574 136600
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 111454 218414 136600
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 115174 222134 136600
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 118894 225854 136600
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 122614 229574 136600
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 129454 236414 136600
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 133174 240134 136600
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 100894 243854 136600
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 104614 247574 136600
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 111454 254414 136600
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 115174 258134 136600
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 118894 261854 136600
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 122614 265574 136600
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 129454 272414 136600
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 133174 276134 136600
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 100894 279854 136600
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 104614 283574 136600
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 111454 290414 136600
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 115174 294134 136600
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 118894 297854 136600
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 122614 301574 136600
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 129454 308414 136600
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 133174 312134 136600
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 100894 315854 136600
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 104614 319574 136600
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 111454 326414 136600
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 115174 330134 136600
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 118894 333854 136600
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 122614 337574 136600
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 129454 344414 136600
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 133174 348134 136600
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 100894 351854 136600
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 104614 355574 136600
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 111454 362414 136600
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 115174 366134 136600
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 118894 369854 136600
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 122614 373574 136600
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 129454 380414 136600
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 133174 384134 136600
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 100894 387854 136600
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 104614 391574 136600
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 111454 398414 136600
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 115174 402134 136600
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 118894 405854 136600
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 122614 409574 136600
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 129454 416414 136600
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 133174 420134 136600
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 100894 423854 136600
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 104614 427574 136600
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 111454 434414 136600
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 115174 438134 136600
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 118894 441854 136600
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 122614 445574 136600
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 129454 452414 136600
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 133174 456134 136600
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 100894 459854 136600
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 104614 463574 136600
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 111454 470414 136600
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 115174 474134 136600
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 118894 477854 136600
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 122614 481574 136600
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 129454 488414 136600
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 133174 492134 136600
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 100894 495854 136600
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 104614 499574 136600
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 111454 506414 136600
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 84050 543218 84286 543454
rect 84050 542898 84286 543134
rect 84050 507218 84286 507454
rect 84050 506898 84286 507134
rect 84050 471218 84286 471454
rect 84050 470898 84286 471134
rect 84050 435218 84286 435454
rect 84050 434898 84286 435134
rect 84050 399218 84286 399454
rect 84050 398898 84286 399134
rect 84050 363218 84286 363454
rect 84050 362898 84286 363134
rect 84050 327218 84286 327454
rect 84050 326898 84286 327134
rect 84050 291218 84286 291454
rect 84050 290898 84286 291134
rect 84050 255218 84286 255454
rect 84050 254898 84286 255134
rect 84050 219218 84286 219454
rect 84050 218898 84286 219134
rect 84050 183218 84286 183454
rect 84050 182898 84286 183134
rect 84050 147218 84286 147454
rect 84050 146898 84286 147134
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 99410 561218 99646 561454
rect 99410 560898 99646 561134
rect 130130 561218 130366 561454
rect 130130 560898 130366 561134
rect 160850 561218 161086 561454
rect 160850 560898 161086 561134
rect 191570 561218 191806 561454
rect 191570 560898 191806 561134
rect 222290 561218 222526 561454
rect 222290 560898 222526 561134
rect 253010 561218 253246 561454
rect 253010 560898 253246 561134
rect 283730 561218 283966 561454
rect 283730 560898 283966 561134
rect 314450 561218 314686 561454
rect 314450 560898 314686 561134
rect 345170 561218 345406 561454
rect 345170 560898 345406 561134
rect 375890 561218 376126 561454
rect 375890 560898 376126 561134
rect 406610 561218 406846 561454
rect 406610 560898 406846 561134
rect 437330 561218 437566 561454
rect 437330 560898 437566 561134
rect 468050 561218 468286 561454
rect 468050 560898 468286 561134
rect 498770 561218 499006 561454
rect 498770 560898 499006 561134
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 114770 543218 115006 543454
rect 114770 542898 115006 543134
rect 145490 543218 145726 543454
rect 145490 542898 145726 543134
rect 176210 543218 176446 543454
rect 176210 542898 176446 543134
rect 206930 543218 207166 543454
rect 206930 542898 207166 543134
rect 237650 543218 237886 543454
rect 237650 542898 237886 543134
rect 268370 543218 268606 543454
rect 268370 542898 268606 543134
rect 299090 543218 299326 543454
rect 299090 542898 299326 543134
rect 329810 543218 330046 543454
rect 329810 542898 330046 543134
rect 360530 543218 360766 543454
rect 360530 542898 360766 543134
rect 391250 543218 391486 543454
rect 391250 542898 391486 543134
rect 421970 543218 422206 543454
rect 421970 542898 422206 543134
rect 452690 543218 452926 543454
rect 452690 542898 452926 543134
rect 483410 543218 483646 543454
rect 483410 542898 483646 543134
rect 99410 525218 99646 525454
rect 99410 524898 99646 525134
rect 130130 525218 130366 525454
rect 130130 524898 130366 525134
rect 160850 525218 161086 525454
rect 160850 524898 161086 525134
rect 191570 525218 191806 525454
rect 191570 524898 191806 525134
rect 222290 525218 222526 525454
rect 222290 524898 222526 525134
rect 253010 525218 253246 525454
rect 253010 524898 253246 525134
rect 283730 525218 283966 525454
rect 283730 524898 283966 525134
rect 314450 525218 314686 525454
rect 314450 524898 314686 525134
rect 345170 525218 345406 525454
rect 345170 524898 345406 525134
rect 375890 525218 376126 525454
rect 375890 524898 376126 525134
rect 406610 525218 406846 525454
rect 406610 524898 406846 525134
rect 437330 525218 437566 525454
rect 437330 524898 437566 525134
rect 468050 525218 468286 525454
rect 468050 524898 468286 525134
rect 498770 525218 499006 525454
rect 498770 524898 499006 525134
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 114770 507218 115006 507454
rect 114770 506898 115006 507134
rect 145490 507218 145726 507454
rect 145490 506898 145726 507134
rect 176210 507218 176446 507454
rect 176210 506898 176446 507134
rect 206930 507218 207166 507454
rect 206930 506898 207166 507134
rect 237650 507218 237886 507454
rect 237650 506898 237886 507134
rect 268370 507218 268606 507454
rect 268370 506898 268606 507134
rect 299090 507218 299326 507454
rect 299090 506898 299326 507134
rect 329810 507218 330046 507454
rect 329810 506898 330046 507134
rect 360530 507218 360766 507454
rect 360530 506898 360766 507134
rect 391250 507218 391486 507454
rect 391250 506898 391486 507134
rect 421970 507218 422206 507454
rect 421970 506898 422206 507134
rect 452690 507218 452926 507454
rect 452690 506898 452926 507134
rect 483410 507218 483646 507454
rect 483410 506898 483646 507134
rect 99410 489218 99646 489454
rect 99410 488898 99646 489134
rect 130130 489218 130366 489454
rect 130130 488898 130366 489134
rect 160850 489218 161086 489454
rect 160850 488898 161086 489134
rect 191570 489218 191806 489454
rect 191570 488898 191806 489134
rect 222290 489218 222526 489454
rect 222290 488898 222526 489134
rect 253010 489218 253246 489454
rect 253010 488898 253246 489134
rect 283730 489218 283966 489454
rect 283730 488898 283966 489134
rect 314450 489218 314686 489454
rect 314450 488898 314686 489134
rect 345170 489218 345406 489454
rect 345170 488898 345406 489134
rect 375890 489218 376126 489454
rect 375890 488898 376126 489134
rect 406610 489218 406846 489454
rect 406610 488898 406846 489134
rect 437330 489218 437566 489454
rect 437330 488898 437566 489134
rect 468050 489218 468286 489454
rect 468050 488898 468286 489134
rect 498770 489218 499006 489454
rect 498770 488898 499006 489134
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 114770 471218 115006 471454
rect 114770 470898 115006 471134
rect 145490 471218 145726 471454
rect 145490 470898 145726 471134
rect 176210 471218 176446 471454
rect 176210 470898 176446 471134
rect 206930 471218 207166 471454
rect 206930 470898 207166 471134
rect 237650 471218 237886 471454
rect 237650 470898 237886 471134
rect 268370 471218 268606 471454
rect 268370 470898 268606 471134
rect 299090 471218 299326 471454
rect 299090 470898 299326 471134
rect 329810 471218 330046 471454
rect 329810 470898 330046 471134
rect 360530 471218 360766 471454
rect 360530 470898 360766 471134
rect 391250 471218 391486 471454
rect 391250 470898 391486 471134
rect 421970 471218 422206 471454
rect 421970 470898 422206 471134
rect 452690 471218 452926 471454
rect 452690 470898 452926 471134
rect 483410 471218 483646 471454
rect 483410 470898 483646 471134
rect 99410 453218 99646 453454
rect 99410 452898 99646 453134
rect 130130 453218 130366 453454
rect 130130 452898 130366 453134
rect 160850 453218 161086 453454
rect 160850 452898 161086 453134
rect 191570 453218 191806 453454
rect 191570 452898 191806 453134
rect 222290 453218 222526 453454
rect 222290 452898 222526 453134
rect 253010 453218 253246 453454
rect 253010 452898 253246 453134
rect 283730 453218 283966 453454
rect 283730 452898 283966 453134
rect 314450 453218 314686 453454
rect 314450 452898 314686 453134
rect 345170 453218 345406 453454
rect 345170 452898 345406 453134
rect 375890 453218 376126 453454
rect 375890 452898 376126 453134
rect 406610 453218 406846 453454
rect 406610 452898 406846 453134
rect 437330 453218 437566 453454
rect 437330 452898 437566 453134
rect 468050 453218 468286 453454
rect 468050 452898 468286 453134
rect 498770 453218 499006 453454
rect 498770 452898 499006 453134
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 114770 435218 115006 435454
rect 114770 434898 115006 435134
rect 145490 435218 145726 435454
rect 145490 434898 145726 435134
rect 176210 435218 176446 435454
rect 176210 434898 176446 435134
rect 206930 435218 207166 435454
rect 206930 434898 207166 435134
rect 237650 435218 237886 435454
rect 237650 434898 237886 435134
rect 268370 435218 268606 435454
rect 268370 434898 268606 435134
rect 299090 435218 299326 435454
rect 299090 434898 299326 435134
rect 329810 435218 330046 435454
rect 329810 434898 330046 435134
rect 360530 435218 360766 435454
rect 360530 434898 360766 435134
rect 391250 435218 391486 435454
rect 391250 434898 391486 435134
rect 421970 435218 422206 435454
rect 421970 434898 422206 435134
rect 452690 435218 452926 435454
rect 452690 434898 452926 435134
rect 483410 435218 483646 435454
rect 483410 434898 483646 435134
rect 99410 417218 99646 417454
rect 99410 416898 99646 417134
rect 130130 417218 130366 417454
rect 130130 416898 130366 417134
rect 160850 417218 161086 417454
rect 160850 416898 161086 417134
rect 191570 417218 191806 417454
rect 191570 416898 191806 417134
rect 222290 417218 222526 417454
rect 222290 416898 222526 417134
rect 253010 417218 253246 417454
rect 253010 416898 253246 417134
rect 283730 417218 283966 417454
rect 283730 416898 283966 417134
rect 314450 417218 314686 417454
rect 314450 416898 314686 417134
rect 345170 417218 345406 417454
rect 345170 416898 345406 417134
rect 375890 417218 376126 417454
rect 375890 416898 376126 417134
rect 406610 417218 406846 417454
rect 406610 416898 406846 417134
rect 437330 417218 437566 417454
rect 437330 416898 437566 417134
rect 468050 417218 468286 417454
rect 468050 416898 468286 417134
rect 498770 417218 499006 417454
rect 498770 416898 499006 417134
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 114770 399218 115006 399454
rect 114770 398898 115006 399134
rect 145490 399218 145726 399454
rect 145490 398898 145726 399134
rect 176210 399218 176446 399454
rect 176210 398898 176446 399134
rect 206930 399218 207166 399454
rect 206930 398898 207166 399134
rect 237650 399218 237886 399454
rect 237650 398898 237886 399134
rect 268370 399218 268606 399454
rect 268370 398898 268606 399134
rect 299090 399218 299326 399454
rect 299090 398898 299326 399134
rect 329810 399218 330046 399454
rect 329810 398898 330046 399134
rect 360530 399218 360766 399454
rect 360530 398898 360766 399134
rect 391250 399218 391486 399454
rect 391250 398898 391486 399134
rect 421970 399218 422206 399454
rect 421970 398898 422206 399134
rect 452690 399218 452926 399454
rect 452690 398898 452926 399134
rect 483410 399218 483646 399454
rect 483410 398898 483646 399134
rect 99410 381218 99646 381454
rect 99410 380898 99646 381134
rect 130130 381218 130366 381454
rect 130130 380898 130366 381134
rect 160850 381218 161086 381454
rect 160850 380898 161086 381134
rect 191570 381218 191806 381454
rect 191570 380898 191806 381134
rect 222290 381218 222526 381454
rect 222290 380898 222526 381134
rect 253010 381218 253246 381454
rect 253010 380898 253246 381134
rect 283730 381218 283966 381454
rect 283730 380898 283966 381134
rect 314450 381218 314686 381454
rect 314450 380898 314686 381134
rect 345170 381218 345406 381454
rect 345170 380898 345406 381134
rect 375890 381218 376126 381454
rect 375890 380898 376126 381134
rect 406610 381218 406846 381454
rect 406610 380898 406846 381134
rect 437330 381218 437566 381454
rect 437330 380898 437566 381134
rect 468050 381218 468286 381454
rect 468050 380898 468286 381134
rect 498770 381218 499006 381454
rect 498770 380898 499006 381134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 114770 363218 115006 363454
rect 114770 362898 115006 363134
rect 145490 363218 145726 363454
rect 145490 362898 145726 363134
rect 176210 363218 176446 363454
rect 176210 362898 176446 363134
rect 206930 363218 207166 363454
rect 206930 362898 207166 363134
rect 237650 363218 237886 363454
rect 237650 362898 237886 363134
rect 268370 363218 268606 363454
rect 268370 362898 268606 363134
rect 299090 363218 299326 363454
rect 299090 362898 299326 363134
rect 329810 363218 330046 363454
rect 329810 362898 330046 363134
rect 360530 363218 360766 363454
rect 360530 362898 360766 363134
rect 391250 363218 391486 363454
rect 391250 362898 391486 363134
rect 421970 363218 422206 363454
rect 421970 362898 422206 363134
rect 452690 363218 452926 363454
rect 452690 362898 452926 363134
rect 483410 363218 483646 363454
rect 483410 362898 483646 363134
rect 99410 345218 99646 345454
rect 99410 344898 99646 345134
rect 130130 345218 130366 345454
rect 130130 344898 130366 345134
rect 160850 345218 161086 345454
rect 160850 344898 161086 345134
rect 191570 345218 191806 345454
rect 191570 344898 191806 345134
rect 222290 345218 222526 345454
rect 222290 344898 222526 345134
rect 253010 345218 253246 345454
rect 253010 344898 253246 345134
rect 283730 345218 283966 345454
rect 283730 344898 283966 345134
rect 314450 345218 314686 345454
rect 314450 344898 314686 345134
rect 345170 345218 345406 345454
rect 345170 344898 345406 345134
rect 375890 345218 376126 345454
rect 375890 344898 376126 345134
rect 406610 345218 406846 345454
rect 406610 344898 406846 345134
rect 437330 345218 437566 345454
rect 437330 344898 437566 345134
rect 468050 345218 468286 345454
rect 468050 344898 468286 345134
rect 498770 345218 499006 345454
rect 498770 344898 499006 345134
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 114770 327218 115006 327454
rect 114770 326898 115006 327134
rect 145490 327218 145726 327454
rect 145490 326898 145726 327134
rect 176210 327218 176446 327454
rect 176210 326898 176446 327134
rect 206930 327218 207166 327454
rect 206930 326898 207166 327134
rect 237650 327218 237886 327454
rect 237650 326898 237886 327134
rect 268370 327218 268606 327454
rect 268370 326898 268606 327134
rect 299090 327218 299326 327454
rect 299090 326898 299326 327134
rect 329810 327218 330046 327454
rect 329810 326898 330046 327134
rect 360530 327218 360766 327454
rect 360530 326898 360766 327134
rect 391250 327218 391486 327454
rect 391250 326898 391486 327134
rect 421970 327218 422206 327454
rect 421970 326898 422206 327134
rect 452690 327218 452926 327454
rect 452690 326898 452926 327134
rect 483410 327218 483646 327454
rect 483410 326898 483646 327134
rect 99410 309218 99646 309454
rect 99410 308898 99646 309134
rect 130130 309218 130366 309454
rect 130130 308898 130366 309134
rect 160850 309218 161086 309454
rect 160850 308898 161086 309134
rect 191570 309218 191806 309454
rect 191570 308898 191806 309134
rect 222290 309218 222526 309454
rect 222290 308898 222526 309134
rect 253010 309218 253246 309454
rect 253010 308898 253246 309134
rect 283730 309218 283966 309454
rect 283730 308898 283966 309134
rect 314450 309218 314686 309454
rect 314450 308898 314686 309134
rect 345170 309218 345406 309454
rect 345170 308898 345406 309134
rect 375890 309218 376126 309454
rect 375890 308898 376126 309134
rect 406610 309218 406846 309454
rect 406610 308898 406846 309134
rect 437330 309218 437566 309454
rect 437330 308898 437566 309134
rect 468050 309218 468286 309454
rect 468050 308898 468286 309134
rect 498770 309218 499006 309454
rect 498770 308898 499006 309134
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 114770 291218 115006 291454
rect 114770 290898 115006 291134
rect 145490 291218 145726 291454
rect 145490 290898 145726 291134
rect 176210 291218 176446 291454
rect 176210 290898 176446 291134
rect 206930 291218 207166 291454
rect 206930 290898 207166 291134
rect 237650 291218 237886 291454
rect 237650 290898 237886 291134
rect 268370 291218 268606 291454
rect 268370 290898 268606 291134
rect 299090 291218 299326 291454
rect 299090 290898 299326 291134
rect 329810 291218 330046 291454
rect 329810 290898 330046 291134
rect 360530 291218 360766 291454
rect 360530 290898 360766 291134
rect 391250 291218 391486 291454
rect 391250 290898 391486 291134
rect 421970 291218 422206 291454
rect 421970 290898 422206 291134
rect 452690 291218 452926 291454
rect 452690 290898 452926 291134
rect 483410 291218 483646 291454
rect 483410 290898 483646 291134
rect 99410 273218 99646 273454
rect 99410 272898 99646 273134
rect 130130 273218 130366 273454
rect 130130 272898 130366 273134
rect 160850 273218 161086 273454
rect 160850 272898 161086 273134
rect 191570 273218 191806 273454
rect 191570 272898 191806 273134
rect 222290 273218 222526 273454
rect 222290 272898 222526 273134
rect 253010 273218 253246 273454
rect 253010 272898 253246 273134
rect 283730 273218 283966 273454
rect 283730 272898 283966 273134
rect 314450 273218 314686 273454
rect 314450 272898 314686 273134
rect 345170 273218 345406 273454
rect 345170 272898 345406 273134
rect 375890 273218 376126 273454
rect 375890 272898 376126 273134
rect 406610 273218 406846 273454
rect 406610 272898 406846 273134
rect 437330 273218 437566 273454
rect 437330 272898 437566 273134
rect 468050 273218 468286 273454
rect 468050 272898 468286 273134
rect 498770 273218 499006 273454
rect 498770 272898 499006 273134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 114770 255218 115006 255454
rect 114770 254898 115006 255134
rect 145490 255218 145726 255454
rect 145490 254898 145726 255134
rect 176210 255218 176446 255454
rect 176210 254898 176446 255134
rect 206930 255218 207166 255454
rect 206930 254898 207166 255134
rect 237650 255218 237886 255454
rect 237650 254898 237886 255134
rect 268370 255218 268606 255454
rect 268370 254898 268606 255134
rect 299090 255218 299326 255454
rect 299090 254898 299326 255134
rect 329810 255218 330046 255454
rect 329810 254898 330046 255134
rect 360530 255218 360766 255454
rect 360530 254898 360766 255134
rect 391250 255218 391486 255454
rect 391250 254898 391486 255134
rect 421970 255218 422206 255454
rect 421970 254898 422206 255134
rect 452690 255218 452926 255454
rect 452690 254898 452926 255134
rect 483410 255218 483646 255454
rect 483410 254898 483646 255134
rect 99410 237218 99646 237454
rect 99410 236898 99646 237134
rect 130130 237218 130366 237454
rect 130130 236898 130366 237134
rect 160850 237218 161086 237454
rect 160850 236898 161086 237134
rect 191570 237218 191806 237454
rect 191570 236898 191806 237134
rect 222290 237218 222526 237454
rect 222290 236898 222526 237134
rect 253010 237218 253246 237454
rect 253010 236898 253246 237134
rect 283730 237218 283966 237454
rect 283730 236898 283966 237134
rect 314450 237218 314686 237454
rect 314450 236898 314686 237134
rect 345170 237218 345406 237454
rect 345170 236898 345406 237134
rect 375890 237218 376126 237454
rect 375890 236898 376126 237134
rect 406610 237218 406846 237454
rect 406610 236898 406846 237134
rect 437330 237218 437566 237454
rect 437330 236898 437566 237134
rect 468050 237218 468286 237454
rect 468050 236898 468286 237134
rect 498770 237218 499006 237454
rect 498770 236898 499006 237134
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 114770 219218 115006 219454
rect 114770 218898 115006 219134
rect 145490 219218 145726 219454
rect 145490 218898 145726 219134
rect 176210 219218 176446 219454
rect 176210 218898 176446 219134
rect 206930 219218 207166 219454
rect 206930 218898 207166 219134
rect 237650 219218 237886 219454
rect 237650 218898 237886 219134
rect 268370 219218 268606 219454
rect 268370 218898 268606 219134
rect 299090 219218 299326 219454
rect 299090 218898 299326 219134
rect 329810 219218 330046 219454
rect 329810 218898 330046 219134
rect 360530 219218 360766 219454
rect 360530 218898 360766 219134
rect 391250 219218 391486 219454
rect 391250 218898 391486 219134
rect 421970 219218 422206 219454
rect 421970 218898 422206 219134
rect 452690 219218 452926 219454
rect 452690 218898 452926 219134
rect 483410 219218 483646 219454
rect 483410 218898 483646 219134
rect 99410 201218 99646 201454
rect 99410 200898 99646 201134
rect 130130 201218 130366 201454
rect 130130 200898 130366 201134
rect 160850 201218 161086 201454
rect 160850 200898 161086 201134
rect 191570 201218 191806 201454
rect 191570 200898 191806 201134
rect 222290 201218 222526 201454
rect 222290 200898 222526 201134
rect 253010 201218 253246 201454
rect 253010 200898 253246 201134
rect 283730 201218 283966 201454
rect 283730 200898 283966 201134
rect 314450 201218 314686 201454
rect 314450 200898 314686 201134
rect 345170 201218 345406 201454
rect 345170 200898 345406 201134
rect 375890 201218 376126 201454
rect 375890 200898 376126 201134
rect 406610 201218 406846 201454
rect 406610 200898 406846 201134
rect 437330 201218 437566 201454
rect 437330 200898 437566 201134
rect 468050 201218 468286 201454
rect 468050 200898 468286 201134
rect 498770 201218 499006 201454
rect 498770 200898 499006 201134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 114770 183218 115006 183454
rect 114770 182898 115006 183134
rect 145490 183218 145726 183454
rect 145490 182898 145726 183134
rect 176210 183218 176446 183454
rect 176210 182898 176446 183134
rect 206930 183218 207166 183454
rect 206930 182898 207166 183134
rect 237650 183218 237886 183454
rect 237650 182898 237886 183134
rect 268370 183218 268606 183454
rect 268370 182898 268606 183134
rect 299090 183218 299326 183454
rect 299090 182898 299326 183134
rect 329810 183218 330046 183454
rect 329810 182898 330046 183134
rect 360530 183218 360766 183454
rect 360530 182898 360766 183134
rect 391250 183218 391486 183454
rect 391250 182898 391486 183134
rect 421970 183218 422206 183454
rect 421970 182898 422206 183134
rect 452690 183218 452926 183454
rect 452690 182898 452926 183134
rect 483410 183218 483646 183454
rect 483410 182898 483646 183134
rect 99410 165218 99646 165454
rect 99410 164898 99646 165134
rect 130130 165218 130366 165454
rect 130130 164898 130366 165134
rect 160850 165218 161086 165454
rect 160850 164898 161086 165134
rect 191570 165218 191806 165454
rect 191570 164898 191806 165134
rect 222290 165218 222526 165454
rect 222290 164898 222526 165134
rect 253010 165218 253246 165454
rect 253010 164898 253246 165134
rect 283730 165218 283966 165454
rect 283730 164898 283966 165134
rect 314450 165218 314686 165454
rect 314450 164898 314686 165134
rect 345170 165218 345406 165454
rect 345170 164898 345406 165134
rect 375890 165218 376126 165454
rect 375890 164898 376126 165134
rect 406610 165218 406846 165454
rect 406610 164898 406846 165134
rect 437330 165218 437566 165454
rect 437330 164898 437566 165134
rect 468050 165218 468286 165454
rect 468050 164898 468286 165134
rect 498770 165218 499006 165454
rect 498770 164898 499006 165134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 114770 147218 115006 147454
rect 114770 146898 115006 147134
rect 145490 147218 145726 147454
rect 145490 146898 145726 147134
rect 176210 147218 176446 147454
rect 176210 146898 176446 147134
rect 206930 147218 207166 147454
rect 206930 146898 207166 147134
rect 237650 147218 237886 147454
rect 237650 146898 237886 147134
rect 268370 147218 268606 147454
rect 268370 146898 268606 147134
rect 299090 147218 299326 147454
rect 299090 146898 299326 147134
rect 329810 147218 330046 147454
rect 329810 146898 330046 147134
rect 360530 147218 360766 147454
rect 360530 146898 360766 147134
rect 391250 147218 391486 147454
rect 391250 146898 391486 147134
rect 421970 147218 422206 147454
rect 421970 146898 422206 147134
rect 452690 147218 452926 147454
rect 452690 146898 452926 147134
rect 483410 147218 483646 147454
rect 483410 146898 483646 147134
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 99410 561454
rect 99646 561218 130130 561454
rect 130366 561218 160850 561454
rect 161086 561218 191570 561454
rect 191806 561218 222290 561454
rect 222526 561218 253010 561454
rect 253246 561218 283730 561454
rect 283966 561218 314450 561454
rect 314686 561218 345170 561454
rect 345406 561218 375890 561454
rect 376126 561218 406610 561454
rect 406846 561218 437330 561454
rect 437566 561218 468050 561454
rect 468286 561218 498770 561454
rect 499006 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 99410 561134
rect 99646 560898 130130 561134
rect 130366 560898 160850 561134
rect 161086 560898 191570 561134
rect 191806 560898 222290 561134
rect 222526 560898 253010 561134
rect 253246 560898 283730 561134
rect 283966 560898 314450 561134
rect 314686 560898 345170 561134
rect 345406 560898 375890 561134
rect 376126 560898 406610 561134
rect 406846 560898 437330 561134
rect 437566 560898 468050 561134
rect 468286 560898 498770 561134
rect 499006 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 84050 543454
rect 84286 543218 114770 543454
rect 115006 543218 145490 543454
rect 145726 543218 176210 543454
rect 176446 543218 206930 543454
rect 207166 543218 237650 543454
rect 237886 543218 268370 543454
rect 268606 543218 299090 543454
rect 299326 543218 329810 543454
rect 330046 543218 360530 543454
rect 360766 543218 391250 543454
rect 391486 543218 421970 543454
rect 422206 543218 452690 543454
rect 452926 543218 483410 543454
rect 483646 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 84050 543134
rect 84286 542898 114770 543134
rect 115006 542898 145490 543134
rect 145726 542898 176210 543134
rect 176446 542898 206930 543134
rect 207166 542898 237650 543134
rect 237886 542898 268370 543134
rect 268606 542898 299090 543134
rect 299326 542898 329810 543134
rect 330046 542898 360530 543134
rect 360766 542898 391250 543134
rect 391486 542898 421970 543134
rect 422206 542898 452690 543134
rect 452926 542898 483410 543134
rect 483646 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 99410 525454
rect 99646 525218 130130 525454
rect 130366 525218 160850 525454
rect 161086 525218 191570 525454
rect 191806 525218 222290 525454
rect 222526 525218 253010 525454
rect 253246 525218 283730 525454
rect 283966 525218 314450 525454
rect 314686 525218 345170 525454
rect 345406 525218 375890 525454
rect 376126 525218 406610 525454
rect 406846 525218 437330 525454
rect 437566 525218 468050 525454
rect 468286 525218 498770 525454
rect 499006 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 99410 525134
rect 99646 524898 130130 525134
rect 130366 524898 160850 525134
rect 161086 524898 191570 525134
rect 191806 524898 222290 525134
rect 222526 524898 253010 525134
rect 253246 524898 283730 525134
rect 283966 524898 314450 525134
rect 314686 524898 345170 525134
rect 345406 524898 375890 525134
rect 376126 524898 406610 525134
rect 406846 524898 437330 525134
rect 437566 524898 468050 525134
rect 468286 524898 498770 525134
rect 499006 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 84050 507454
rect 84286 507218 114770 507454
rect 115006 507218 145490 507454
rect 145726 507218 176210 507454
rect 176446 507218 206930 507454
rect 207166 507218 237650 507454
rect 237886 507218 268370 507454
rect 268606 507218 299090 507454
rect 299326 507218 329810 507454
rect 330046 507218 360530 507454
rect 360766 507218 391250 507454
rect 391486 507218 421970 507454
rect 422206 507218 452690 507454
rect 452926 507218 483410 507454
rect 483646 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 84050 507134
rect 84286 506898 114770 507134
rect 115006 506898 145490 507134
rect 145726 506898 176210 507134
rect 176446 506898 206930 507134
rect 207166 506898 237650 507134
rect 237886 506898 268370 507134
rect 268606 506898 299090 507134
rect 299326 506898 329810 507134
rect 330046 506898 360530 507134
rect 360766 506898 391250 507134
rect 391486 506898 421970 507134
rect 422206 506898 452690 507134
rect 452926 506898 483410 507134
rect 483646 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 99410 489454
rect 99646 489218 130130 489454
rect 130366 489218 160850 489454
rect 161086 489218 191570 489454
rect 191806 489218 222290 489454
rect 222526 489218 253010 489454
rect 253246 489218 283730 489454
rect 283966 489218 314450 489454
rect 314686 489218 345170 489454
rect 345406 489218 375890 489454
rect 376126 489218 406610 489454
rect 406846 489218 437330 489454
rect 437566 489218 468050 489454
rect 468286 489218 498770 489454
rect 499006 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 99410 489134
rect 99646 488898 130130 489134
rect 130366 488898 160850 489134
rect 161086 488898 191570 489134
rect 191806 488898 222290 489134
rect 222526 488898 253010 489134
rect 253246 488898 283730 489134
rect 283966 488898 314450 489134
rect 314686 488898 345170 489134
rect 345406 488898 375890 489134
rect 376126 488898 406610 489134
rect 406846 488898 437330 489134
rect 437566 488898 468050 489134
rect 468286 488898 498770 489134
rect 499006 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 84050 471454
rect 84286 471218 114770 471454
rect 115006 471218 145490 471454
rect 145726 471218 176210 471454
rect 176446 471218 206930 471454
rect 207166 471218 237650 471454
rect 237886 471218 268370 471454
rect 268606 471218 299090 471454
rect 299326 471218 329810 471454
rect 330046 471218 360530 471454
rect 360766 471218 391250 471454
rect 391486 471218 421970 471454
rect 422206 471218 452690 471454
rect 452926 471218 483410 471454
rect 483646 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 84050 471134
rect 84286 470898 114770 471134
rect 115006 470898 145490 471134
rect 145726 470898 176210 471134
rect 176446 470898 206930 471134
rect 207166 470898 237650 471134
rect 237886 470898 268370 471134
rect 268606 470898 299090 471134
rect 299326 470898 329810 471134
rect 330046 470898 360530 471134
rect 360766 470898 391250 471134
rect 391486 470898 421970 471134
rect 422206 470898 452690 471134
rect 452926 470898 483410 471134
rect 483646 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 99410 453454
rect 99646 453218 130130 453454
rect 130366 453218 160850 453454
rect 161086 453218 191570 453454
rect 191806 453218 222290 453454
rect 222526 453218 253010 453454
rect 253246 453218 283730 453454
rect 283966 453218 314450 453454
rect 314686 453218 345170 453454
rect 345406 453218 375890 453454
rect 376126 453218 406610 453454
rect 406846 453218 437330 453454
rect 437566 453218 468050 453454
rect 468286 453218 498770 453454
rect 499006 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 99410 453134
rect 99646 452898 130130 453134
rect 130366 452898 160850 453134
rect 161086 452898 191570 453134
rect 191806 452898 222290 453134
rect 222526 452898 253010 453134
rect 253246 452898 283730 453134
rect 283966 452898 314450 453134
rect 314686 452898 345170 453134
rect 345406 452898 375890 453134
rect 376126 452898 406610 453134
rect 406846 452898 437330 453134
rect 437566 452898 468050 453134
rect 468286 452898 498770 453134
rect 499006 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 84050 435454
rect 84286 435218 114770 435454
rect 115006 435218 145490 435454
rect 145726 435218 176210 435454
rect 176446 435218 206930 435454
rect 207166 435218 237650 435454
rect 237886 435218 268370 435454
rect 268606 435218 299090 435454
rect 299326 435218 329810 435454
rect 330046 435218 360530 435454
rect 360766 435218 391250 435454
rect 391486 435218 421970 435454
rect 422206 435218 452690 435454
rect 452926 435218 483410 435454
rect 483646 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 84050 435134
rect 84286 434898 114770 435134
rect 115006 434898 145490 435134
rect 145726 434898 176210 435134
rect 176446 434898 206930 435134
rect 207166 434898 237650 435134
rect 237886 434898 268370 435134
rect 268606 434898 299090 435134
rect 299326 434898 329810 435134
rect 330046 434898 360530 435134
rect 360766 434898 391250 435134
rect 391486 434898 421970 435134
rect 422206 434898 452690 435134
rect 452926 434898 483410 435134
rect 483646 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 99410 417454
rect 99646 417218 130130 417454
rect 130366 417218 160850 417454
rect 161086 417218 191570 417454
rect 191806 417218 222290 417454
rect 222526 417218 253010 417454
rect 253246 417218 283730 417454
rect 283966 417218 314450 417454
rect 314686 417218 345170 417454
rect 345406 417218 375890 417454
rect 376126 417218 406610 417454
rect 406846 417218 437330 417454
rect 437566 417218 468050 417454
rect 468286 417218 498770 417454
rect 499006 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 99410 417134
rect 99646 416898 130130 417134
rect 130366 416898 160850 417134
rect 161086 416898 191570 417134
rect 191806 416898 222290 417134
rect 222526 416898 253010 417134
rect 253246 416898 283730 417134
rect 283966 416898 314450 417134
rect 314686 416898 345170 417134
rect 345406 416898 375890 417134
rect 376126 416898 406610 417134
rect 406846 416898 437330 417134
rect 437566 416898 468050 417134
rect 468286 416898 498770 417134
rect 499006 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 84050 399454
rect 84286 399218 114770 399454
rect 115006 399218 145490 399454
rect 145726 399218 176210 399454
rect 176446 399218 206930 399454
rect 207166 399218 237650 399454
rect 237886 399218 268370 399454
rect 268606 399218 299090 399454
rect 299326 399218 329810 399454
rect 330046 399218 360530 399454
rect 360766 399218 391250 399454
rect 391486 399218 421970 399454
rect 422206 399218 452690 399454
rect 452926 399218 483410 399454
rect 483646 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 84050 399134
rect 84286 398898 114770 399134
rect 115006 398898 145490 399134
rect 145726 398898 176210 399134
rect 176446 398898 206930 399134
rect 207166 398898 237650 399134
rect 237886 398898 268370 399134
rect 268606 398898 299090 399134
rect 299326 398898 329810 399134
rect 330046 398898 360530 399134
rect 360766 398898 391250 399134
rect 391486 398898 421970 399134
rect 422206 398898 452690 399134
rect 452926 398898 483410 399134
rect 483646 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 99410 381454
rect 99646 381218 130130 381454
rect 130366 381218 160850 381454
rect 161086 381218 191570 381454
rect 191806 381218 222290 381454
rect 222526 381218 253010 381454
rect 253246 381218 283730 381454
rect 283966 381218 314450 381454
rect 314686 381218 345170 381454
rect 345406 381218 375890 381454
rect 376126 381218 406610 381454
rect 406846 381218 437330 381454
rect 437566 381218 468050 381454
rect 468286 381218 498770 381454
rect 499006 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 99410 381134
rect 99646 380898 130130 381134
rect 130366 380898 160850 381134
rect 161086 380898 191570 381134
rect 191806 380898 222290 381134
rect 222526 380898 253010 381134
rect 253246 380898 283730 381134
rect 283966 380898 314450 381134
rect 314686 380898 345170 381134
rect 345406 380898 375890 381134
rect 376126 380898 406610 381134
rect 406846 380898 437330 381134
rect 437566 380898 468050 381134
rect 468286 380898 498770 381134
rect 499006 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 84050 363454
rect 84286 363218 114770 363454
rect 115006 363218 145490 363454
rect 145726 363218 176210 363454
rect 176446 363218 206930 363454
rect 207166 363218 237650 363454
rect 237886 363218 268370 363454
rect 268606 363218 299090 363454
rect 299326 363218 329810 363454
rect 330046 363218 360530 363454
rect 360766 363218 391250 363454
rect 391486 363218 421970 363454
rect 422206 363218 452690 363454
rect 452926 363218 483410 363454
rect 483646 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 84050 363134
rect 84286 362898 114770 363134
rect 115006 362898 145490 363134
rect 145726 362898 176210 363134
rect 176446 362898 206930 363134
rect 207166 362898 237650 363134
rect 237886 362898 268370 363134
rect 268606 362898 299090 363134
rect 299326 362898 329810 363134
rect 330046 362898 360530 363134
rect 360766 362898 391250 363134
rect 391486 362898 421970 363134
rect 422206 362898 452690 363134
rect 452926 362898 483410 363134
rect 483646 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 99410 345454
rect 99646 345218 130130 345454
rect 130366 345218 160850 345454
rect 161086 345218 191570 345454
rect 191806 345218 222290 345454
rect 222526 345218 253010 345454
rect 253246 345218 283730 345454
rect 283966 345218 314450 345454
rect 314686 345218 345170 345454
rect 345406 345218 375890 345454
rect 376126 345218 406610 345454
rect 406846 345218 437330 345454
rect 437566 345218 468050 345454
rect 468286 345218 498770 345454
rect 499006 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 99410 345134
rect 99646 344898 130130 345134
rect 130366 344898 160850 345134
rect 161086 344898 191570 345134
rect 191806 344898 222290 345134
rect 222526 344898 253010 345134
rect 253246 344898 283730 345134
rect 283966 344898 314450 345134
rect 314686 344898 345170 345134
rect 345406 344898 375890 345134
rect 376126 344898 406610 345134
rect 406846 344898 437330 345134
rect 437566 344898 468050 345134
rect 468286 344898 498770 345134
rect 499006 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 84050 327454
rect 84286 327218 114770 327454
rect 115006 327218 145490 327454
rect 145726 327218 176210 327454
rect 176446 327218 206930 327454
rect 207166 327218 237650 327454
rect 237886 327218 268370 327454
rect 268606 327218 299090 327454
rect 299326 327218 329810 327454
rect 330046 327218 360530 327454
rect 360766 327218 391250 327454
rect 391486 327218 421970 327454
rect 422206 327218 452690 327454
rect 452926 327218 483410 327454
rect 483646 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 84050 327134
rect 84286 326898 114770 327134
rect 115006 326898 145490 327134
rect 145726 326898 176210 327134
rect 176446 326898 206930 327134
rect 207166 326898 237650 327134
rect 237886 326898 268370 327134
rect 268606 326898 299090 327134
rect 299326 326898 329810 327134
rect 330046 326898 360530 327134
rect 360766 326898 391250 327134
rect 391486 326898 421970 327134
rect 422206 326898 452690 327134
rect 452926 326898 483410 327134
rect 483646 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 99410 309454
rect 99646 309218 130130 309454
rect 130366 309218 160850 309454
rect 161086 309218 191570 309454
rect 191806 309218 222290 309454
rect 222526 309218 253010 309454
rect 253246 309218 283730 309454
rect 283966 309218 314450 309454
rect 314686 309218 345170 309454
rect 345406 309218 375890 309454
rect 376126 309218 406610 309454
rect 406846 309218 437330 309454
rect 437566 309218 468050 309454
rect 468286 309218 498770 309454
rect 499006 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 99410 309134
rect 99646 308898 130130 309134
rect 130366 308898 160850 309134
rect 161086 308898 191570 309134
rect 191806 308898 222290 309134
rect 222526 308898 253010 309134
rect 253246 308898 283730 309134
rect 283966 308898 314450 309134
rect 314686 308898 345170 309134
rect 345406 308898 375890 309134
rect 376126 308898 406610 309134
rect 406846 308898 437330 309134
rect 437566 308898 468050 309134
rect 468286 308898 498770 309134
rect 499006 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 84050 291454
rect 84286 291218 114770 291454
rect 115006 291218 145490 291454
rect 145726 291218 176210 291454
rect 176446 291218 206930 291454
rect 207166 291218 237650 291454
rect 237886 291218 268370 291454
rect 268606 291218 299090 291454
rect 299326 291218 329810 291454
rect 330046 291218 360530 291454
rect 360766 291218 391250 291454
rect 391486 291218 421970 291454
rect 422206 291218 452690 291454
rect 452926 291218 483410 291454
rect 483646 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 84050 291134
rect 84286 290898 114770 291134
rect 115006 290898 145490 291134
rect 145726 290898 176210 291134
rect 176446 290898 206930 291134
rect 207166 290898 237650 291134
rect 237886 290898 268370 291134
rect 268606 290898 299090 291134
rect 299326 290898 329810 291134
rect 330046 290898 360530 291134
rect 360766 290898 391250 291134
rect 391486 290898 421970 291134
rect 422206 290898 452690 291134
rect 452926 290898 483410 291134
rect 483646 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 99410 273454
rect 99646 273218 130130 273454
rect 130366 273218 160850 273454
rect 161086 273218 191570 273454
rect 191806 273218 222290 273454
rect 222526 273218 253010 273454
rect 253246 273218 283730 273454
rect 283966 273218 314450 273454
rect 314686 273218 345170 273454
rect 345406 273218 375890 273454
rect 376126 273218 406610 273454
rect 406846 273218 437330 273454
rect 437566 273218 468050 273454
rect 468286 273218 498770 273454
rect 499006 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 99410 273134
rect 99646 272898 130130 273134
rect 130366 272898 160850 273134
rect 161086 272898 191570 273134
rect 191806 272898 222290 273134
rect 222526 272898 253010 273134
rect 253246 272898 283730 273134
rect 283966 272898 314450 273134
rect 314686 272898 345170 273134
rect 345406 272898 375890 273134
rect 376126 272898 406610 273134
rect 406846 272898 437330 273134
rect 437566 272898 468050 273134
rect 468286 272898 498770 273134
rect 499006 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 84050 255454
rect 84286 255218 114770 255454
rect 115006 255218 145490 255454
rect 145726 255218 176210 255454
rect 176446 255218 206930 255454
rect 207166 255218 237650 255454
rect 237886 255218 268370 255454
rect 268606 255218 299090 255454
rect 299326 255218 329810 255454
rect 330046 255218 360530 255454
rect 360766 255218 391250 255454
rect 391486 255218 421970 255454
rect 422206 255218 452690 255454
rect 452926 255218 483410 255454
rect 483646 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 84050 255134
rect 84286 254898 114770 255134
rect 115006 254898 145490 255134
rect 145726 254898 176210 255134
rect 176446 254898 206930 255134
rect 207166 254898 237650 255134
rect 237886 254898 268370 255134
rect 268606 254898 299090 255134
rect 299326 254898 329810 255134
rect 330046 254898 360530 255134
rect 360766 254898 391250 255134
rect 391486 254898 421970 255134
rect 422206 254898 452690 255134
rect 452926 254898 483410 255134
rect 483646 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 99410 237454
rect 99646 237218 130130 237454
rect 130366 237218 160850 237454
rect 161086 237218 191570 237454
rect 191806 237218 222290 237454
rect 222526 237218 253010 237454
rect 253246 237218 283730 237454
rect 283966 237218 314450 237454
rect 314686 237218 345170 237454
rect 345406 237218 375890 237454
rect 376126 237218 406610 237454
rect 406846 237218 437330 237454
rect 437566 237218 468050 237454
rect 468286 237218 498770 237454
rect 499006 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 99410 237134
rect 99646 236898 130130 237134
rect 130366 236898 160850 237134
rect 161086 236898 191570 237134
rect 191806 236898 222290 237134
rect 222526 236898 253010 237134
rect 253246 236898 283730 237134
rect 283966 236898 314450 237134
rect 314686 236898 345170 237134
rect 345406 236898 375890 237134
rect 376126 236898 406610 237134
rect 406846 236898 437330 237134
rect 437566 236898 468050 237134
rect 468286 236898 498770 237134
rect 499006 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 84050 219454
rect 84286 219218 114770 219454
rect 115006 219218 145490 219454
rect 145726 219218 176210 219454
rect 176446 219218 206930 219454
rect 207166 219218 237650 219454
rect 237886 219218 268370 219454
rect 268606 219218 299090 219454
rect 299326 219218 329810 219454
rect 330046 219218 360530 219454
rect 360766 219218 391250 219454
rect 391486 219218 421970 219454
rect 422206 219218 452690 219454
rect 452926 219218 483410 219454
rect 483646 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 84050 219134
rect 84286 218898 114770 219134
rect 115006 218898 145490 219134
rect 145726 218898 176210 219134
rect 176446 218898 206930 219134
rect 207166 218898 237650 219134
rect 237886 218898 268370 219134
rect 268606 218898 299090 219134
rect 299326 218898 329810 219134
rect 330046 218898 360530 219134
rect 360766 218898 391250 219134
rect 391486 218898 421970 219134
rect 422206 218898 452690 219134
rect 452926 218898 483410 219134
rect 483646 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 99410 201454
rect 99646 201218 130130 201454
rect 130366 201218 160850 201454
rect 161086 201218 191570 201454
rect 191806 201218 222290 201454
rect 222526 201218 253010 201454
rect 253246 201218 283730 201454
rect 283966 201218 314450 201454
rect 314686 201218 345170 201454
rect 345406 201218 375890 201454
rect 376126 201218 406610 201454
rect 406846 201218 437330 201454
rect 437566 201218 468050 201454
rect 468286 201218 498770 201454
rect 499006 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 99410 201134
rect 99646 200898 130130 201134
rect 130366 200898 160850 201134
rect 161086 200898 191570 201134
rect 191806 200898 222290 201134
rect 222526 200898 253010 201134
rect 253246 200898 283730 201134
rect 283966 200898 314450 201134
rect 314686 200898 345170 201134
rect 345406 200898 375890 201134
rect 376126 200898 406610 201134
rect 406846 200898 437330 201134
rect 437566 200898 468050 201134
rect 468286 200898 498770 201134
rect 499006 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 84050 183454
rect 84286 183218 114770 183454
rect 115006 183218 145490 183454
rect 145726 183218 176210 183454
rect 176446 183218 206930 183454
rect 207166 183218 237650 183454
rect 237886 183218 268370 183454
rect 268606 183218 299090 183454
rect 299326 183218 329810 183454
rect 330046 183218 360530 183454
rect 360766 183218 391250 183454
rect 391486 183218 421970 183454
rect 422206 183218 452690 183454
rect 452926 183218 483410 183454
rect 483646 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 84050 183134
rect 84286 182898 114770 183134
rect 115006 182898 145490 183134
rect 145726 182898 176210 183134
rect 176446 182898 206930 183134
rect 207166 182898 237650 183134
rect 237886 182898 268370 183134
rect 268606 182898 299090 183134
rect 299326 182898 329810 183134
rect 330046 182898 360530 183134
rect 360766 182898 391250 183134
rect 391486 182898 421970 183134
rect 422206 182898 452690 183134
rect 452926 182898 483410 183134
rect 483646 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 99410 165454
rect 99646 165218 130130 165454
rect 130366 165218 160850 165454
rect 161086 165218 191570 165454
rect 191806 165218 222290 165454
rect 222526 165218 253010 165454
rect 253246 165218 283730 165454
rect 283966 165218 314450 165454
rect 314686 165218 345170 165454
rect 345406 165218 375890 165454
rect 376126 165218 406610 165454
rect 406846 165218 437330 165454
rect 437566 165218 468050 165454
rect 468286 165218 498770 165454
rect 499006 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 99410 165134
rect 99646 164898 130130 165134
rect 130366 164898 160850 165134
rect 161086 164898 191570 165134
rect 191806 164898 222290 165134
rect 222526 164898 253010 165134
rect 253246 164898 283730 165134
rect 283966 164898 314450 165134
rect 314686 164898 345170 165134
rect 345406 164898 375890 165134
rect 376126 164898 406610 165134
rect 406846 164898 437330 165134
rect 437566 164898 468050 165134
rect 468286 164898 498770 165134
rect 499006 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 84050 147454
rect 84286 147218 114770 147454
rect 115006 147218 145490 147454
rect 145726 147218 176210 147454
rect 176446 147218 206930 147454
rect 207166 147218 237650 147454
rect 237886 147218 268370 147454
rect 268606 147218 299090 147454
rect 299326 147218 329810 147454
rect 330046 147218 360530 147454
rect 360766 147218 391250 147454
rect 391486 147218 421970 147454
rect 422206 147218 452690 147454
rect 452926 147218 483410 147454
rect 483646 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 84050 147134
rect 84286 146898 114770 147134
rect 115006 146898 145490 147134
rect 145726 146898 176210 147134
rect 176446 146898 206930 147134
rect 207166 146898 237650 147134
rect 237886 146898 268370 147134
rect 268606 146898 299090 147134
rect 299326 146898 329810 147134
rect 330046 146898 360530 147134
rect 360766 146898 391250 147134
rect 391486 146898 421970 147134
rect 422206 146898 452690 147134
rect 452926 146898 483410 147134
rect 483646 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1636617456
transform 1 0 79800 0 1 138600
box 382 0 424551 426704
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 136600 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 567304 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 567304 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 567304 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 567304 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 567304 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 567304 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 567304 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 567304 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 567304 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 567304 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 567304 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 567304 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 136600 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 567304 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 567304 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 567304 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 567304 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 567304 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 567304 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 567304 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 567304 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 567304 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 567304 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 567304 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 567304 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 136600 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 567304 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 567304 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 567304 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 567304 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 567304 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 567304 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 567304 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 567304 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 567304 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 567304 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 567304 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 567304 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 136600 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 567304 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 567304 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 567304 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 567304 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 567304 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 567304 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 567304 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 567304 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 567304 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 567304 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 567304 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 567304 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 136600 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 567304 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 567304 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 567304 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 567304 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 567304 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 567304 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 567304 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 567304 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 567304 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 567304 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 567304 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 567304 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 136600 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 567304 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 567304 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 567304 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 567304 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 567304 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 567304 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 567304 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 567304 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 567304 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 567304 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 567304 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 567304 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 136600 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 567304 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 567304 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 567304 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 567304 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 567304 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 567304 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 567304 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 567304 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 567304 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 567304 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 567304 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 567304 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 136600 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 567304 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 567304 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 567304 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 567304 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 567304 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 567304 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 567304 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 567304 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 567304 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 567304 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 567304 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 567304 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
