magic
tech sky130A
magscale 1 2
timestamp 1635436522
<< obsli1 >>
rect 1104 1377 446016 445009
<< obsm1 >>
rect 382 76 446738 445120
<< metal2 >>
rect 1950 446400 2006 447200
rect 5814 446400 5870 447200
rect 9770 446400 9826 447200
rect 13634 446400 13690 447200
rect 17590 446400 17646 447200
rect 21546 446400 21602 447200
rect 25410 446400 25466 447200
rect 29366 446400 29422 447200
rect 33322 446400 33378 447200
rect 37186 446400 37242 447200
rect 41142 446400 41198 447200
rect 45098 446400 45154 447200
rect 48962 446400 49018 447200
rect 52918 446400 52974 447200
rect 56782 446400 56838 447200
rect 60738 446400 60794 447200
rect 64694 446400 64750 447200
rect 68558 446400 68614 447200
rect 72514 446400 72570 447200
rect 76470 446400 76526 447200
rect 80334 446400 80390 447200
rect 84290 446400 84346 447200
rect 88246 446400 88302 447200
rect 92110 446400 92166 447200
rect 96066 446400 96122 447200
rect 100022 446400 100078 447200
rect 103886 446400 103942 447200
rect 107842 446400 107898 447200
rect 111706 446400 111762 447200
rect 115662 446400 115718 447200
rect 119618 446400 119674 447200
rect 123482 446400 123538 447200
rect 127438 446400 127494 447200
rect 131394 446400 131450 447200
rect 135258 446400 135314 447200
rect 139214 446400 139270 447200
rect 143170 446400 143226 447200
rect 147034 446400 147090 447200
rect 150990 446400 151046 447200
rect 154854 446400 154910 447200
rect 158810 446400 158866 447200
rect 162766 446400 162822 447200
rect 166630 446400 166686 447200
rect 170586 446400 170642 447200
rect 174542 446400 174598 447200
rect 178406 446400 178462 447200
rect 182362 446400 182418 447200
rect 186318 446400 186374 447200
rect 190182 446400 190238 447200
rect 194138 446400 194194 447200
rect 198094 446400 198150 447200
rect 201958 446400 202014 447200
rect 205914 446400 205970 447200
rect 209778 446400 209834 447200
rect 213734 446400 213790 447200
rect 217690 446400 217746 447200
rect 221554 446400 221610 447200
rect 225510 446400 225566 447200
rect 229466 446400 229522 447200
rect 233330 446400 233386 447200
rect 237286 446400 237342 447200
rect 241242 446400 241298 447200
rect 245106 446400 245162 447200
rect 249062 446400 249118 447200
rect 252926 446400 252982 447200
rect 256882 446400 256938 447200
rect 260838 446400 260894 447200
rect 264702 446400 264758 447200
rect 268658 446400 268714 447200
rect 272614 446400 272670 447200
rect 276478 446400 276534 447200
rect 280434 446400 280490 447200
rect 284390 446400 284446 447200
rect 288254 446400 288310 447200
rect 292210 446400 292266 447200
rect 296166 446400 296222 447200
rect 300030 446400 300086 447200
rect 303986 446400 304042 447200
rect 307850 446400 307906 447200
rect 311806 446400 311862 447200
rect 315762 446400 315818 447200
rect 319626 446400 319682 447200
rect 323582 446400 323638 447200
rect 327538 446400 327594 447200
rect 331402 446400 331458 447200
rect 335358 446400 335414 447200
rect 339314 446400 339370 447200
rect 343178 446400 343234 447200
rect 347134 446400 347190 447200
rect 350998 446400 351054 447200
rect 354954 446400 355010 447200
rect 358910 446400 358966 447200
rect 362774 446400 362830 447200
rect 366730 446400 366786 447200
rect 370686 446400 370742 447200
rect 374550 446400 374606 447200
rect 378506 446400 378562 447200
rect 382462 446400 382518 447200
rect 386326 446400 386382 447200
rect 390282 446400 390338 447200
rect 394238 446400 394294 447200
rect 398102 446400 398158 447200
rect 402058 446400 402114 447200
rect 405922 446400 405978 447200
rect 409878 446400 409934 447200
rect 413834 446400 413890 447200
rect 417698 446400 417754 447200
rect 421654 446400 421710 447200
rect 425610 446400 425666 447200
rect 429474 446400 429530 447200
rect 433430 446400 433486 447200
rect 437386 446400 437442 447200
rect 441250 446400 441306 447200
rect 445206 446400 445262 447200
rect 386 0 442 800
rect 1214 0 1270 800
rect 2134 0 2190 800
rect 3054 0 3110 800
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15750 0 15806 800
rect 16670 0 16726 800
rect 17590 0 17646 800
rect 18510 0 18566 800
rect 19430 0 19486 800
rect 20258 0 20314 800
rect 21178 0 21234 800
rect 22098 0 22154 800
rect 23018 0 23074 800
rect 23938 0 23994 800
rect 24858 0 24914 800
rect 25778 0 25834 800
rect 26606 0 26662 800
rect 27526 0 27582 800
rect 28446 0 28502 800
rect 29366 0 29422 800
rect 30286 0 30342 800
rect 31206 0 31262 800
rect 32126 0 32182 800
rect 32954 0 33010 800
rect 33874 0 33930 800
rect 34794 0 34850 800
rect 35714 0 35770 800
rect 36634 0 36690 800
rect 37554 0 37610 800
rect 38474 0 38530 800
rect 39302 0 39358 800
rect 40222 0 40278 800
rect 41142 0 41198 800
rect 42062 0 42118 800
rect 42982 0 43038 800
rect 43902 0 43958 800
rect 44822 0 44878 800
rect 45742 0 45798 800
rect 46570 0 46626 800
rect 47490 0 47546 800
rect 48410 0 48466 800
rect 49330 0 49386 800
rect 50250 0 50306 800
rect 51170 0 51226 800
rect 52090 0 52146 800
rect 52918 0 52974 800
rect 53838 0 53894 800
rect 54758 0 54814 800
rect 55678 0 55734 800
rect 56598 0 56654 800
rect 57518 0 57574 800
rect 58438 0 58494 800
rect 59266 0 59322 800
rect 60186 0 60242 800
rect 61106 0 61162 800
rect 62026 0 62082 800
rect 62946 0 63002 800
rect 63866 0 63922 800
rect 64786 0 64842 800
rect 65614 0 65670 800
rect 66534 0 66590 800
rect 67454 0 67510 800
rect 68374 0 68430 800
rect 69294 0 69350 800
rect 70214 0 70270 800
rect 71134 0 71190 800
rect 71962 0 72018 800
rect 72882 0 72938 800
rect 73802 0 73858 800
rect 74722 0 74778 800
rect 75642 0 75698 800
rect 76562 0 76618 800
rect 77482 0 77538 800
rect 78310 0 78366 800
rect 79230 0 79286 800
rect 80150 0 80206 800
rect 81070 0 81126 800
rect 81990 0 82046 800
rect 82910 0 82966 800
rect 83830 0 83886 800
rect 84658 0 84714 800
rect 85578 0 85634 800
rect 86498 0 86554 800
rect 87418 0 87474 800
rect 88338 0 88394 800
rect 89258 0 89314 800
rect 90178 0 90234 800
rect 91098 0 91154 800
rect 91926 0 91982 800
rect 92846 0 92902 800
rect 93766 0 93822 800
rect 94686 0 94742 800
rect 95606 0 95662 800
rect 96526 0 96582 800
rect 97446 0 97502 800
rect 98274 0 98330 800
rect 99194 0 99250 800
rect 100114 0 100170 800
rect 101034 0 101090 800
rect 101954 0 102010 800
rect 102874 0 102930 800
rect 103794 0 103850 800
rect 104622 0 104678 800
rect 105542 0 105598 800
rect 106462 0 106518 800
rect 107382 0 107438 800
rect 108302 0 108358 800
rect 109222 0 109278 800
rect 110142 0 110198 800
rect 110970 0 111026 800
rect 111890 0 111946 800
rect 112810 0 112866 800
rect 113730 0 113786 800
rect 114650 0 114706 800
rect 115570 0 115626 800
rect 116490 0 116546 800
rect 117318 0 117374 800
rect 118238 0 118294 800
rect 119158 0 119214 800
rect 120078 0 120134 800
rect 120998 0 121054 800
rect 121918 0 121974 800
rect 122838 0 122894 800
rect 123666 0 123722 800
rect 124586 0 124642 800
rect 125506 0 125562 800
rect 126426 0 126482 800
rect 127346 0 127402 800
rect 128266 0 128322 800
rect 129186 0 129242 800
rect 130014 0 130070 800
rect 130934 0 130990 800
rect 131854 0 131910 800
rect 132774 0 132830 800
rect 133694 0 133750 800
rect 134614 0 134670 800
rect 135534 0 135590 800
rect 136454 0 136510 800
rect 137282 0 137338 800
rect 138202 0 138258 800
rect 139122 0 139178 800
rect 140042 0 140098 800
rect 140962 0 141018 800
rect 141882 0 141938 800
rect 142802 0 142858 800
rect 143630 0 143686 800
rect 144550 0 144606 800
rect 145470 0 145526 800
rect 146390 0 146446 800
rect 147310 0 147366 800
rect 148230 0 148286 800
rect 149150 0 149206 800
rect 149978 0 150034 800
rect 150898 0 150954 800
rect 151818 0 151874 800
rect 152738 0 152794 800
rect 153658 0 153714 800
rect 154578 0 154634 800
rect 155498 0 155554 800
rect 156326 0 156382 800
rect 157246 0 157302 800
rect 158166 0 158222 800
rect 159086 0 159142 800
rect 160006 0 160062 800
rect 160926 0 160982 800
rect 161846 0 161902 800
rect 162674 0 162730 800
rect 163594 0 163650 800
rect 164514 0 164570 800
rect 165434 0 165490 800
rect 166354 0 166410 800
rect 167274 0 167330 800
rect 168194 0 168250 800
rect 169022 0 169078 800
rect 169942 0 169998 800
rect 170862 0 170918 800
rect 171782 0 171838 800
rect 172702 0 172758 800
rect 173622 0 173678 800
rect 174542 0 174598 800
rect 175370 0 175426 800
rect 176290 0 176346 800
rect 177210 0 177266 800
rect 178130 0 178186 800
rect 179050 0 179106 800
rect 179970 0 180026 800
rect 180890 0 180946 800
rect 181810 0 181866 800
rect 182638 0 182694 800
rect 183558 0 183614 800
rect 184478 0 184534 800
rect 185398 0 185454 800
rect 186318 0 186374 800
rect 187238 0 187294 800
rect 188158 0 188214 800
rect 188986 0 189042 800
rect 189906 0 189962 800
rect 190826 0 190882 800
rect 191746 0 191802 800
rect 192666 0 192722 800
rect 193586 0 193642 800
rect 194506 0 194562 800
rect 195334 0 195390 800
rect 196254 0 196310 800
rect 197174 0 197230 800
rect 198094 0 198150 800
rect 199014 0 199070 800
rect 199934 0 199990 800
rect 200854 0 200910 800
rect 201682 0 201738 800
rect 202602 0 202658 800
rect 203522 0 203578 800
rect 204442 0 204498 800
rect 205362 0 205418 800
rect 206282 0 206338 800
rect 207202 0 207258 800
rect 208030 0 208086 800
rect 208950 0 209006 800
rect 209870 0 209926 800
rect 210790 0 210846 800
rect 211710 0 211766 800
rect 212630 0 212686 800
rect 213550 0 213606 800
rect 214378 0 214434 800
rect 215298 0 215354 800
rect 216218 0 216274 800
rect 217138 0 217194 800
rect 218058 0 218114 800
rect 218978 0 219034 800
rect 219898 0 219954 800
rect 220726 0 220782 800
rect 221646 0 221702 800
rect 222566 0 222622 800
rect 223486 0 223542 800
rect 224406 0 224462 800
rect 225326 0 225382 800
rect 226246 0 226302 800
rect 227166 0 227222 800
rect 227994 0 228050 800
rect 228914 0 228970 800
rect 229834 0 229890 800
rect 230754 0 230810 800
rect 231674 0 231730 800
rect 232594 0 232650 800
rect 233514 0 233570 800
rect 234342 0 234398 800
rect 235262 0 235318 800
rect 236182 0 236238 800
rect 237102 0 237158 800
rect 238022 0 238078 800
rect 238942 0 238998 800
rect 239862 0 239918 800
rect 240690 0 240746 800
rect 241610 0 241666 800
rect 242530 0 242586 800
rect 243450 0 243506 800
rect 244370 0 244426 800
rect 245290 0 245346 800
rect 246210 0 246266 800
rect 247038 0 247094 800
rect 247958 0 248014 800
rect 248878 0 248934 800
rect 249798 0 249854 800
rect 250718 0 250774 800
rect 251638 0 251694 800
rect 252558 0 252614 800
rect 253386 0 253442 800
rect 254306 0 254362 800
rect 255226 0 255282 800
rect 256146 0 256202 800
rect 257066 0 257122 800
rect 257986 0 258042 800
rect 258906 0 258962 800
rect 259734 0 259790 800
rect 260654 0 260710 800
rect 261574 0 261630 800
rect 262494 0 262550 800
rect 263414 0 263470 800
rect 264334 0 264390 800
rect 265254 0 265310 800
rect 266082 0 266138 800
rect 267002 0 267058 800
rect 267922 0 267978 800
rect 268842 0 268898 800
rect 269762 0 269818 800
rect 270682 0 270738 800
rect 271602 0 271658 800
rect 272522 0 272578 800
rect 273350 0 273406 800
rect 274270 0 274326 800
rect 275190 0 275246 800
rect 276110 0 276166 800
rect 277030 0 277086 800
rect 277950 0 278006 800
rect 278870 0 278926 800
rect 279698 0 279754 800
rect 280618 0 280674 800
rect 281538 0 281594 800
rect 282458 0 282514 800
rect 283378 0 283434 800
rect 284298 0 284354 800
rect 285218 0 285274 800
rect 286046 0 286102 800
rect 286966 0 287022 800
rect 287886 0 287942 800
rect 288806 0 288862 800
rect 289726 0 289782 800
rect 290646 0 290702 800
rect 291566 0 291622 800
rect 292394 0 292450 800
rect 293314 0 293370 800
rect 294234 0 294290 800
rect 295154 0 295210 800
rect 296074 0 296130 800
rect 296994 0 297050 800
rect 297914 0 297970 800
rect 298742 0 298798 800
rect 299662 0 299718 800
rect 300582 0 300638 800
rect 301502 0 301558 800
rect 302422 0 302478 800
rect 303342 0 303398 800
rect 304262 0 304318 800
rect 305090 0 305146 800
rect 306010 0 306066 800
rect 306930 0 306986 800
rect 307850 0 307906 800
rect 308770 0 308826 800
rect 309690 0 309746 800
rect 310610 0 310666 800
rect 311438 0 311494 800
rect 312358 0 312414 800
rect 313278 0 313334 800
rect 314198 0 314254 800
rect 315118 0 315174 800
rect 316038 0 316094 800
rect 316958 0 317014 800
rect 317878 0 317934 800
rect 318706 0 318762 800
rect 319626 0 319682 800
rect 320546 0 320602 800
rect 321466 0 321522 800
rect 322386 0 322442 800
rect 323306 0 323362 800
rect 324226 0 324282 800
rect 325054 0 325110 800
rect 325974 0 326030 800
rect 326894 0 326950 800
rect 327814 0 327870 800
rect 328734 0 328790 800
rect 329654 0 329710 800
rect 330574 0 330630 800
rect 331402 0 331458 800
rect 332322 0 332378 800
rect 333242 0 333298 800
rect 334162 0 334218 800
rect 335082 0 335138 800
rect 336002 0 336058 800
rect 336922 0 336978 800
rect 337750 0 337806 800
rect 338670 0 338726 800
rect 339590 0 339646 800
rect 340510 0 340566 800
rect 341430 0 341486 800
rect 342350 0 342406 800
rect 343270 0 343326 800
rect 344098 0 344154 800
rect 345018 0 345074 800
rect 345938 0 345994 800
rect 346858 0 346914 800
rect 347778 0 347834 800
rect 348698 0 348754 800
rect 349618 0 349674 800
rect 350446 0 350502 800
rect 351366 0 351422 800
rect 352286 0 352342 800
rect 353206 0 353262 800
rect 354126 0 354182 800
rect 355046 0 355102 800
rect 355966 0 356022 800
rect 356794 0 356850 800
rect 357714 0 357770 800
rect 358634 0 358690 800
rect 359554 0 359610 800
rect 360474 0 360530 800
rect 361394 0 361450 800
rect 362314 0 362370 800
rect 363234 0 363290 800
rect 364062 0 364118 800
rect 364982 0 365038 800
rect 365902 0 365958 800
rect 366822 0 366878 800
rect 367742 0 367798 800
rect 368662 0 368718 800
rect 369582 0 369638 800
rect 370410 0 370466 800
rect 371330 0 371386 800
rect 372250 0 372306 800
rect 373170 0 373226 800
rect 374090 0 374146 800
rect 375010 0 375066 800
rect 375930 0 375986 800
rect 376758 0 376814 800
rect 377678 0 377734 800
rect 378598 0 378654 800
rect 379518 0 379574 800
rect 380438 0 380494 800
rect 381358 0 381414 800
rect 382278 0 382334 800
rect 383106 0 383162 800
rect 384026 0 384082 800
rect 384946 0 385002 800
rect 385866 0 385922 800
rect 386786 0 386842 800
rect 387706 0 387762 800
rect 388626 0 388682 800
rect 389454 0 389510 800
rect 390374 0 390430 800
rect 391294 0 391350 800
rect 392214 0 392270 800
rect 393134 0 393190 800
rect 394054 0 394110 800
rect 394974 0 395030 800
rect 395802 0 395858 800
rect 396722 0 396778 800
rect 397642 0 397698 800
rect 398562 0 398618 800
rect 399482 0 399538 800
rect 400402 0 400458 800
rect 401322 0 401378 800
rect 402150 0 402206 800
rect 403070 0 403126 800
rect 403990 0 404046 800
rect 404910 0 404966 800
rect 405830 0 405886 800
rect 406750 0 406806 800
rect 407670 0 407726 800
rect 408590 0 408646 800
rect 409418 0 409474 800
rect 410338 0 410394 800
rect 411258 0 411314 800
rect 412178 0 412234 800
rect 413098 0 413154 800
rect 414018 0 414074 800
rect 414938 0 414994 800
rect 415766 0 415822 800
rect 416686 0 416742 800
rect 417606 0 417662 800
rect 418526 0 418582 800
rect 419446 0 419502 800
rect 420366 0 420422 800
rect 421286 0 421342 800
rect 422114 0 422170 800
rect 423034 0 423090 800
rect 423954 0 424010 800
rect 424874 0 424930 800
rect 425794 0 425850 800
rect 426714 0 426770 800
rect 427634 0 427690 800
rect 428462 0 428518 800
rect 429382 0 429438 800
rect 430302 0 430358 800
rect 431222 0 431278 800
rect 432142 0 432198 800
rect 433062 0 433118 800
rect 433982 0 434038 800
rect 434810 0 434866 800
rect 435730 0 435786 800
rect 436650 0 436706 800
rect 437570 0 437626 800
rect 438490 0 438546 800
rect 439410 0 439466 800
rect 440330 0 440386 800
rect 441158 0 441214 800
rect 442078 0 442134 800
rect 442998 0 443054 800
rect 443918 0 443974 800
rect 444838 0 444894 800
rect 445758 0 445814 800
rect 446678 0 446734 800
<< obsm2 >>
rect 388 446344 1894 446434
rect 2062 446344 5758 446434
rect 5926 446344 9714 446434
rect 9882 446344 13578 446434
rect 13746 446344 17534 446434
rect 17702 446344 21490 446434
rect 21658 446344 25354 446434
rect 25522 446344 29310 446434
rect 29478 446344 33266 446434
rect 33434 446344 37130 446434
rect 37298 446344 41086 446434
rect 41254 446344 45042 446434
rect 45210 446344 48906 446434
rect 49074 446344 52862 446434
rect 53030 446344 56726 446434
rect 56894 446344 60682 446434
rect 60850 446344 64638 446434
rect 64806 446344 68502 446434
rect 68670 446344 72458 446434
rect 72626 446344 76414 446434
rect 76582 446344 80278 446434
rect 80446 446344 84234 446434
rect 84402 446344 88190 446434
rect 88358 446344 92054 446434
rect 92222 446344 96010 446434
rect 96178 446344 99966 446434
rect 100134 446344 103830 446434
rect 103998 446344 107786 446434
rect 107954 446344 111650 446434
rect 111818 446344 115606 446434
rect 115774 446344 119562 446434
rect 119730 446344 123426 446434
rect 123594 446344 127382 446434
rect 127550 446344 131338 446434
rect 131506 446344 135202 446434
rect 135370 446344 139158 446434
rect 139326 446344 143114 446434
rect 143282 446344 146978 446434
rect 147146 446344 150934 446434
rect 151102 446344 154798 446434
rect 154966 446344 158754 446434
rect 158922 446344 162710 446434
rect 162878 446344 166574 446434
rect 166742 446344 170530 446434
rect 170698 446344 174486 446434
rect 174654 446344 178350 446434
rect 178518 446344 182306 446434
rect 182474 446344 186262 446434
rect 186430 446344 190126 446434
rect 190294 446344 194082 446434
rect 194250 446344 198038 446434
rect 198206 446344 201902 446434
rect 202070 446344 205858 446434
rect 206026 446344 209722 446434
rect 209890 446344 213678 446434
rect 213846 446344 217634 446434
rect 217802 446344 221498 446434
rect 221666 446344 225454 446434
rect 225622 446344 229410 446434
rect 229578 446344 233274 446434
rect 233442 446344 237230 446434
rect 237398 446344 241186 446434
rect 241354 446344 245050 446434
rect 245218 446344 249006 446434
rect 249174 446344 252870 446434
rect 253038 446344 256826 446434
rect 256994 446344 260782 446434
rect 260950 446344 264646 446434
rect 264814 446344 268602 446434
rect 268770 446344 272558 446434
rect 272726 446344 276422 446434
rect 276590 446344 280378 446434
rect 280546 446344 284334 446434
rect 284502 446344 288198 446434
rect 288366 446344 292154 446434
rect 292322 446344 296110 446434
rect 296278 446344 299974 446434
rect 300142 446344 303930 446434
rect 304098 446344 307794 446434
rect 307962 446344 311750 446434
rect 311918 446344 315706 446434
rect 315874 446344 319570 446434
rect 319738 446344 323526 446434
rect 323694 446344 327482 446434
rect 327650 446344 331346 446434
rect 331514 446344 335302 446434
rect 335470 446344 339258 446434
rect 339426 446344 343122 446434
rect 343290 446344 347078 446434
rect 347246 446344 350942 446434
rect 351110 446344 354898 446434
rect 355066 446344 358854 446434
rect 359022 446344 362718 446434
rect 362886 446344 366674 446434
rect 366842 446344 370630 446434
rect 370798 446344 374494 446434
rect 374662 446344 378450 446434
rect 378618 446344 382406 446434
rect 382574 446344 386270 446434
rect 386438 446344 390226 446434
rect 390394 446344 394182 446434
rect 394350 446344 398046 446434
rect 398214 446344 402002 446434
rect 402170 446344 405866 446434
rect 406034 446344 409822 446434
rect 409990 446344 413778 446434
rect 413946 446344 417642 446434
rect 417810 446344 421598 446434
rect 421766 446344 425554 446434
rect 425722 446344 429418 446434
rect 429586 446344 433374 446434
rect 433542 446344 437330 446434
rect 437498 446344 441194 446434
rect 441362 446344 445150 446434
rect 445318 446344 446732 446434
rect 388 856 446732 446344
rect 498 70 1158 856
rect 1326 70 2078 856
rect 2246 70 2998 856
rect 3166 70 3918 856
rect 4086 70 4838 856
rect 5006 70 5758 856
rect 5926 70 6678 856
rect 6846 70 7506 856
rect 7674 70 8426 856
rect 8594 70 9346 856
rect 9514 70 10266 856
rect 10434 70 11186 856
rect 11354 70 12106 856
rect 12274 70 13026 856
rect 13194 70 13854 856
rect 14022 70 14774 856
rect 14942 70 15694 856
rect 15862 70 16614 856
rect 16782 70 17534 856
rect 17702 70 18454 856
rect 18622 70 19374 856
rect 19542 70 20202 856
rect 20370 70 21122 856
rect 21290 70 22042 856
rect 22210 70 22962 856
rect 23130 70 23882 856
rect 24050 70 24802 856
rect 24970 70 25722 856
rect 25890 70 26550 856
rect 26718 70 27470 856
rect 27638 70 28390 856
rect 28558 70 29310 856
rect 29478 70 30230 856
rect 30398 70 31150 856
rect 31318 70 32070 856
rect 32238 70 32898 856
rect 33066 70 33818 856
rect 33986 70 34738 856
rect 34906 70 35658 856
rect 35826 70 36578 856
rect 36746 70 37498 856
rect 37666 70 38418 856
rect 38586 70 39246 856
rect 39414 70 40166 856
rect 40334 70 41086 856
rect 41254 70 42006 856
rect 42174 70 42926 856
rect 43094 70 43846 856
rect 44014 70 44766 856
rect 44934 70 45686 856
rect 45854 70 46514 856
rect 46682 70 47434 856
rect 47602 70 48354 856
rect 48522 70 49274 856
rect 49442 70 50194 856
rect 50362 70 51114 856
rect 51282 70 52034 856
rect 52202 70 52862 856
rect 53030 70 53782 856
rect 53950 70 54702 856
rect 54870 70 55622 856
rect 55790 70 56542 856
rect 56710 70 57462 856
rect 57630 70 58382 856
rect 58550 70 59210 856
rect 59378 70 60130 856
rect 60298 70 61050 856
rect 61218 70 61970 856
rect 62138 70 62890 856
rect 63058 70 63810 856
rect 63978 70 64730 856
rect 64898 70 65558 856
rect 65726 70 66478 856
rect 66646 70 67398 856
rect 67566 70 68318 856
rect 68486 70 69238 856
rect 69406 70 70158 856
rect 70326 70 71078 856
rect 71246 70 71906 856
rect 72074 70 72826 856
rect 72994 70 73746 856
rect 73914 70 74666 856
rect 74834 70 75586 856
rect 75754 70 76506 856
rect 76674 70 77426 856
rect 77594 70 78254 856
rect 78422 70 79174 856
rect 79342 70 80094 856
rect 80262 70 81014 856
rect 81182 70 81934 856
rect 82102 70 82854 856
rect 83022 70 83774 856
rect 83942 70 84602 856
rect 84770 70 85522 856
rect 85690 70 86442 856
rect 86610 70 87362 856
rect 87530 70 88282 856
rect 88450 70 89202 856
rect 89370 70 90122 856
rect 90290 70 91042 856
rect 91210 70 91870 856
rect 92038 70 92790 856
rect 92958 70 93710 856
rect 93878 70 94630 856
rect 94798 70 95550 856
rect 95718 70 96470 856
rect 96638 70 97390 856
rect 97558 70 98218 856
rect 98386 70 99138 856
rect 99306 70 100058 856
rect 100226 70 100978 856
rect 101146 70 101898 856
rect 102066 70 102818 856
rect 102986 70 103738 856
rect 103906 70 104566 856
rect 104734 70 105486 856
rect 105654 70 106406 856
rect 106574 70 107326 856
rect 107494 70 108246 856
rect 108414 70 109166 856
rect 109334 70 110086 856
rect 110254 70 110914 856
rect 111082 70 111834 856
rect 112002 70 112754 856
rect 112922 70 113674 856
rect 113842 70 114594 856
rect 114762 70 115514 856
rect 115682 70 116434 856
rect 116602 70 117262 856
rect 117430 70 118182 856
rect 118350 70 119102 856
rect 119270 70 120022 856
rect 120190 70 120942 856
rect 121110 70 121862 856
rect 122030 70 122782 856
rect 122950 70 123610 856
rect 123778 70 124530 856
rect 124698 70 125450 856
rect 125618 70 126370 856
rect 126538 70 127290 856
rect 127458 70 128210 856
rect 128378 70 129130 856
rect 129298 70 129958 856
rect 130126 70 130878 856
rect 131046 70 131798 856
rect 131966 70 132718 856
rect 132886 70 133638 856
rect 133806 70 134558 856
rect 134726 70 135478 856
rect 135646 70 136398 856
rect 136566 70 137226 856
rect 137394 70 138146 856
rect 138314 70 139066 856
rect 139234 70 139986 856
rect 140154 70 140906 856
rect 141074 70 141826 856
rect 141994 70 142746 856
rect 142914 70 143574 856
rect 143742 70 144494 856
rect 144662 70 145414 856
rect 145582 70 146334 856
rect 146502 70 147254 856
rect 147422 70 148174 856
rect 148342 70 149094 856
rect 149262 70 149922 856
rect 150090 70 150842 856
rect 151010 70 151762 856
rect 151930 70 152682 856
rect 152850 70 153602 856
rect 153770 70 154522 856
rect 154690 70 155442 856
rect 155610 70 156270 856
rect 156438 70 157190 856
rect 157358 70 158110 856
rect 158278 70 159030 856
rect 159198 70 159950 856
rect 160118 70 160870 856
rect 161038 70 161790 856
rect 161958 70 162618 856
rect 162786 70 163538 856
rect 163706 70 164458 856
rect 164626 70 165378 856
rect 165546 70 166298 856
rect 166466 70 167218 856
rect 167386 70 168138 856
rect 168306 70 168966 856
rect 169134 70 169886 856
rect 170054 70 170806 856
rect 170974 70 171726 856
rect 171894 70 172646 856
rect 172814 70 173566 856
rect 173734 70 174486 856
rect 174654 70 175314 856
rect 175482 70 176234 856
rect 176402 70 177154 856
rect 177322 70 178074 856
rect 178242 70 178994 856
rect 179162 70 179914 856
rect 180082 70 180834 856
rect 181002 70 181754 856
rect 181922 70 182582 856
rect 182750 70 183502 856
rect 183670 70 184422 856
rect 184590 70 185342 856
rect 185510 70 186262 856
rect 186430 70 187182 856
rect 187350 70 188102 856
rect 188270 70 188930 856
rect 189098 70 189850 856
rect 190018 70 190770 856
rect 190938 70 191690 856
rect 191858 70 192610 856
rect 192778 70 193530 856
rect 193698 70 194450 856
rect 194618 70 195278 856
rect 195446 70 196198 856
rect 196366 70 197118 856
rect 197286 70 198038 856
rect 198206 70 198958 856
rect 199126 70 199878 856
rect 200046 70 200798 856
rect 200966 70 201626 856
rect 201794 70 202546 856
rect 202714 70 203466 856
rect 203634 70 204386 856
rect 204554 70 205306 856
rect 205474 70 206226 856
rect 206394 70 207146 856
rect 207314 70 207974 856
rect 208142 70 208894 856
rect 209062 70 209814 856
rect 209982 70 210734 856
rect 210902 70 211654 856
rect 211822 70 212574 856
rect 212742 70 213494 856
rect 213662 70 214322 856
rect 214490 70 215242 856
rect 215410 70 216162 856
rect 216330 70 217082 856
rect 217250 70 218002 856
rect 218170 70 218922 856
rect 219090 70 219842 856
rect 220010 70 220670 856
rect 220838 70 221590 856
rect 221758 70 222510 856
rect 222678 70 223430 856
rect 223598 70 224350 856
rect 224518 70 225270 856
rect 225438 70 226190 856
rect 226358 70 227110 856
rect 227278 70 227938 856
rect 228106 70 228858 856
rect 229026 70 229778 856
rect 229946 70 230698 856
rect 230866 70 231618 856
rect 231786 70 232538 856
rect 232706 70 233458 856
rect 233626 70 234286 856
rect 234454 70 235206 856
rect 235374 70 236126 856
rect 236294 70 237046 856
rect 237214 70 237966 856
rect 238134 70 238886 856
rect 239054 70 239806 856
rect 239974 70 240634 856
rect 240802 70 241554 856
rect 241722 70 242474 856
rect 242642 70 243394 856
rect 243562 70 244314 856
rect 244482 70 245234 856
rect 245402 70 246154 856
rect 246322 70 246982 856
rect 247150 70 247902 856
rect 248070 70 248822 856
rect 248990 70 249742 856
rect 249910 70 250662 856
rect 250830 70 251582 856
rect 251750 70 252502 856
rect 252670 70 253330 856
rect 253498 70 254250 856
rect 254418 70 255170 856
rect 255338 70 256090 856
rect 256258 70 257010 856
rect 257178 70 257930 856
rect 258098 70 258850 856
rect 259018 70 259678 856
rect 259846 70 260598 856
rect 260766 70 261518 856
rect 261686 70 262438 856
rect 262606 70 263358 856
rect 263526 70 264278 856
rect 264446 70 265198 856
rect 265366 70 266026 856
rect 266194 70 266946 856
rect 267114 70 267866 856
rect 268034 70 268786 856
rect 268954 70 269706 856
rect 269874 70 270626 856
rect 270794 70 271546 856
rect 271714 70 272466 856
rect 272634 70 273294 856
rect 273462 70 274214 856
rect 274382 70 275134 856
rect 275302 70 276054 856
rect 276222 70 276974 856
rect 277142 70 277894 856
rect 278062 70 278814 856
rect 278982 70 279642 856
rect 279810 70 280562 856
rect 280730 70 281482 856
rect 281650 70 282402 856
rect 282570 70 283322 856
rect 283490 70 284242 856
rect 284410 70 285162 856
rect 285330 70 285990 856
rect 286158 70 286910 856
rect 287078 70 287830 856
rect 287998 70 288750 856
rect 288918 70 289670 856
rect 289838 70 290590 856
rect 290758 70 291510 856
rect 291678 70 292338 856
rect 292506 70 293258 856
rect 293426 70 294178 856
rect 294346 70 295098 856
rect 295266 70 296018 856
rect 296186 70 296938 856
rect 297106 70 297858 856
rect 298026 70 298686 856
rect 298854 70 299606 856
rect 299774 70 300526 856
rect 300694 70 301446 856
rect 301614 70 302366 856
rect 302534 70 303286 856
rect 303454 70 304206 856
rect 304374 70 305034 856
rect 305202 70 305954 856
rect 306122 70 306874 856
rect 307042 70 307794 856
rect 307962 70 308714 856
rect 308882 70 309634 856
rect 309802 70 310554 856
rect 310722 70 311382 856
rect 311550 70 312302 856
rect 312470 70 313222 856
rect 313390 70 314142 856
rect 314310 70 315062 856
rect 315230 70 315982 856
rect 316150 70 316902 856
rect 317070 70 317822 856
rect 317990 70 318650 856
rect 318818 70 319570 856
rect 319738 70 320490 856
rect 320658 70 321410 856
rect 321578 70 322330 856
rect 322498 70 323250 856
rect 323418 70 324170 856
rect 324338 70 324998 856
rect 325166 70 325918 856
rect 326086 70 326838 856
rect 327006 70 327758 856
rect 327926 70 328678 856
rect 328846 70 329598 856
rect 329766 70 330518 856
rect 330686 70 331346 856
rect 331514 70 332266 856
rect 332434 70 333186 856
rect 333354 70 334106 856
rect 334274 70 335026 856
rect 335194 70 335946 856
rect 336114 70 336866 856
rect 337034 70 337694 856
rect 337862 70 338614 856
rect 338782 70 339534 856
rect 339702 70 340454 856
rect 340622 70 341374 856
rect 341542 70 342294 856
rect 342462 70 343214 856
rect 343382 70 344042 856
rect 344210 70 344962 856
rect 345130 70 345882 856
rect 346050 70 346802 856
rect 346970 70 347722 856
rect 347890 70 348642 856
rect 348810 70 349562 856
rect 349730 70 350390 856
rect 350558 70 351310 856
rect 351478 70 352230 856
rect 352398 70 353150 856
rect 353318 70 354070 856
rect 354238 70 354990 856
rect 355158 70 355910 856
rect 356078 70 356738 856
rect 356906 70 357658 856
rect 357826 70 358578 856
rect 358746 70 359498 856
rect 359666 70 360418 856
rect 360586 70 361338 856
rect 361506 70 362258 856
rect 362426 70 363178 856
rect 363346 70 364006 856
rect 364174 70 364926 856
rect 365094 70 365846 856
rect 366014 70 366766 856
rect 366934 70 367686 856
rect 367854 70 368606 856
rect 368774 70 369526 856
rect 369694 70 370354 856
rect 370522 70 371274 856
rect 371442 70 372194 856
rect 372362 70 373114 856
rect 373282 70 374034 856
rect 374202 70 374954 856
rect 375122 70 375874 856
rect 376042 70 376702 856
rect 376870 70 377622 856
rect 377790 70 378542 856
rect 378710 70 379462 856
rect 379630 70 380382 856
rect 380550 70 381302 856
rect 381470 70 382222 856
rect 382390 70 383050 856
rect 383218 70 383970 856
rect 384138 70 384890 856
rect 385058 70 385810 856
rect 385978 70 386730 856
rect 386898 70 387650 856
rect 387818 70 388570 856
rect 388738 70 389398 856
rect 389566 70 390318 856
rect 390486 70 391238 856
rect 391406 70 392158 856
rect 392326 70 393078 856
rect 393246 70 393998 856
rect 394166 70 394918 856
rect 395086 70 395746 856
rect 395914 70 396666 856
rect 396834 70 397586 856
rect 397754 70 398506 856
rect 398674 70 399426 856
rect 399594 70 400346 856
rect 400514 70 401266 856
rect 401434 70 402094 856
rect 402262 70 403014 856
rect 403182 70 403934 856
rect 404102 70 404854 856
rect 405022 70 405774 856
rect 405942 70 406694 856
rect 406862 70 407614 856
rect 407782 70 408534 856
rect 408702 70 409362 856
rect 409530 70 410282 856
rect 410450 70 411202 856
rect 411370 70 412122 856
rect 412290 70 413042 856
rect 413210 70 413962 856
rect 414130 70 414882 856
rect 415050 70 415710 856
rect 415878 70 416630 856
rect 416798 70 417550 856
rect 417718 70 418470 856
rect 418638 70 419390 856
rect 419558 70 420310 856
rect 420478 70 421230 856
rect 421398 70 422058 856
rect 422226 70 422978 856
rect 423146 70 423898 856
rect 424066 70 424818 856
rect 424986 70 425738 856
rect 425906 70 426658 856
rect 426826 70 427578 856
rect 427746 70 428406 856
rect 428574 70 429326 856
rect 429494 70 430246 856
rect 430414 70 431166 856
rect 431334 70 432086 856
rect 432254 70 433006 856
rect 433174 70 433926 856
rect 434094 70 434754 856
rect 434922 70 435674 856
rect 435842 70 436594 856
rect 436762 70 437514 856
rect 437682 70 438434 856
rect 438602 70 439354 856
rect 439522 70 440274 856
rect 440442 70 441102 856
rect 441270 70 442022 856
rect 442190 70 442942 856
rect 443110 70 443862 856
rect 444030 70 444782 856
rect 444950 70 445702 856
rect 445870 70 446622 856
<< obsm3 >>
rect 4208 579 434608 445025
<< metal4 >>
rect 4208 2128 4528 445040
rect 19568 2128 19888 445040
rect 34928 2128 35248 445040
rect 50288 2128 50608 445040
rect 65648 2128 65968 445040
rect 81008 2128 81328 445040
rect 96368 2128 96688 445040
rect 111728 2128 112048 445040
rect 127088 2128 127408 445040
rect 142448 2128 142768 445040
rect 157808 2128 158128 445040
rect 173168 2128 173488 445040
rect 188528 2128 188848 445040
rect 203888 2128 204208 445040
rect 219248 2128 219568 445040
rect 234608 2128 234928 445040
rect 249968 2128 250288 445040
rect 265328 2128 265648 445040
rect 280688 2128 281008 445040
rect 296048 2128 296368 445040
rect 311408 2128 311728 445040
rect 326768 2128 327088 445040
rect 342128 2128 342448 445040
rect 357488 2128 357808 445040
rect 372848 2128 373168 445040
rect 388208 2128 388528 445040
rect 403568 2128 403888 445040
rect 418928 2128 419248 445040
rect 434288 2128 434608 445040
<< obsm4 >>
rect 58019 2075 65568 328405
rect 66048 2075 80928 328405
rect 81408 2075 96288 328405
rect 96768 2075 111648 328405
rect 112128 2075 127008 328405
rect 127488 2075 142368 328405
rect 142848 2075 157728 328405
rect 158208 2075 173088 328405
rect 173568 2075 188448 328405
rect 188928 2075 203808 328405
rect 204288 2075 219168 328405
rect 219648 2075 234528 328405
rect 235008 2075 249888 328405
rect 250368 2075 265248 328405
rect 265728 2075 280608 328405
rect 281088 2075 295968 328405
rect 296448 2075 311328 328405
rect 311808 2075 326688 328405
rect 327168 2075 342048 328405
rect 342528 2075 357408 328405
rect 357888 2075 367205 328405
<< labels >>
rlabel metal2 s 1950 446400 2006 447200 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 119618 446400 119674 447200 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 131394 446400 131450 447200 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 143170 446400 143226 447200 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 154854 446400 154910 447200 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 166630 446400 166686 447200 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 178406 446400 178462 447200 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 190182 446400 190238 447200 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 201958 446400 202014 447200 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 213734 446400 213790 447200 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 225510 446400 225566 447200 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 13634 446400 13690 447200 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 237286 446400 237342 447200 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 249062 446400 249118 447200 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 260838 446400 260894 447200 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 272614 446400 272670 447200 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 284390 446400 284446 447200 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 296166 446400 296222 447200 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 307850 446400 307906 447200 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 319626 446400 319682 447200 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 331402 446400 331458 447200 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 343178 446400 343234 447200 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 25410 446400 25466 447200 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 354954 446400 355010 447200 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 366730 446400 366786 447200 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 378506 446400 378562 447200 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 390282 446400 390338 447200 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 402058 446400 402114 447200 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 413834 446400 413890 447200 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 425610 446400 425666 447200 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 437386 446400 437442 447200 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 37186 446400 37242 447200 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 48962 446400 49018 447200 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 60738 446400 60794 447200 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 72514 446400 72570 447200 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 84290 446400 84346 447200 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 96066 446400 96122 447200 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 107842 446400 107898 447200 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5814 446400 5870 447200 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 123482 446400 123538 447200 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 135258 446400 135314 447200 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 147034 446400 147090 447200 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 158810 446400 158866 447200 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 170586 446400 170642 447200 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 182362 446400 182418 447200 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 194138 446400 194194 447200 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 205914 446400 205970 447200 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 217690 446400 217746 447200 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 229466 446400 229522 447200 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 17590 446400 17646 447200 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 241242 446400 241298 447200 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 252926 446400 252982 447200 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 264702 446400 264758 447200 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 276478 446400 276534 447200 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 288254 446400 288310 447200 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 300030 446400 300086 447200 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 311806 446400 311862 447200 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 323582 446400 323638 447200 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 335358 446400 335414 447200 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 347134 446400 347190 447200 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 29366 446400 29422 447200 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 358910 446400 358966 447200 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 370686 446400 370742 447200 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 382462 446400 382518 447200 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 394238 446400 394294 447200 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 405922 446400 405978 447200 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 417698 446400 417754 447200 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 429474 446400 429530 447200 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 441250 446400 441306 447200 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 41142 446400 41198 447200 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 52918 446400 52974 447200 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 64694 446400 64750 447200 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 76470 446400 76526 447200 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 88246 446400 88302 447200 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 100022 446400 100078 447200 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 111706 446400 111762 447200 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9770 446400 9826 447200 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 127438 446400 127494 447200 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 139214 446400 139270 447200 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 150990 446400 151046 447200 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 162766 446400 162822 447200 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 174542 446400 174598 447200 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 186318 446400 186374 447200 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 198094 446400 198150 447200 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 209778 446400 209834 447200 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 221554 446400 221610 447200 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 233330 446400 233386 447200 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 21546 446400 21602 447200 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 245106 446400 245162 447200 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 256882 446400 256938 447200 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 268658 446400 268714 447200 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 280434 446400 280490 447200 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 292210 446400 292266 447200 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 303986 446400 304042 447200 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 315762 446400 315818 447200 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 327538 446400 327594 447200 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 339314 446400 339370 447200 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 350998 446400 351054 447200 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 33322 446400 33378 447200 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 362774 446400 362830 447200 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 374550 446400 374606 447200 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 386326 446400 386382 447200 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 398102 446400 398158 447200 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 409878 446400 409934 447200 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 421654 446400 421710 447200 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 433430 446400 433486 447200 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 445206 446400 445262 447200 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 45098 446400 45154 447200 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 56782 446400 56838 447200 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 68558 446400 68614 447200 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 80334 446400 80390 447200 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 92110 446400 92166 447200 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 103886 446400 103942 447200 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 115662 446400 115718 447200 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 444838 0 444894 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 445758 0 445814 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 446678 0 446734 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 368662 0 368718 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 371330 0 371386 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 374090 0 374146 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 376758 0 376814 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 379518 0 379574 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 382278 0 382334 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 384946 0 385002 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 387706 0 387762 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 390374 0 390430 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 393134 0 393190 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 395802 0 395858 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 398562 0 398618 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 401322 0 401378 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 403990 0 404046 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 406750 0 406806 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 409418 0 409474 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 412178 0 412234 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 414938 0 414994 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 417606 0 417662 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 420366 0 420422 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 423034 0 423090 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 425794 0 425850 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 428462 0 428518 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 431222 0 431278 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 433982 0 434038 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 436650 0 436706 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 439410 0 439466 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 442078 0 442134 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 172702 0 172758 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 180890 0 180946 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 188986 0 189042 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 191746 0 191802 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 197174 0 197230 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 205362 0 205418 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 213550 0 213606 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 216218 0 216274 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 218978 0 219034 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 224406 0 224462 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 227166 0 227222 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 229834 0 229890 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 232594 0 232650 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 235262 0 235318 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 240690 0 240746 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 243450 0 243506 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 246210 0 246266 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 248878 0 248934 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 251638 0 251694 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 254306 0 254362 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 257066 0 257122 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 259734 0 259790 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 262494 0 262550 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 265254 0 265310 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 267922 0 267978 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 270682 0 270738 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 273350 0 273406 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 276110 0 276166 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 278870 0 278926 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 281538 0 281594 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 284298 0 284354 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 286966 0 287022 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 289726 0 289782 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 292394 0 292450 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 295154 0 295210 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 297914 0 297970 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 300582 0 300638 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 303342 0 303398 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 306010 0 306066 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 308770 0 308826 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 311438 0 311494 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 314198 0 314254 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 316958 0 317014 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 319626 0 319682 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 322386 0 322442 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 325054 0 325110 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 327814 0 327870 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 330574 0 330630 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 333242 0 333298 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 336002 0 336058 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 338670 0 338726 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 341430 0 341486 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 344098 0 344154 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 346858 0 346914 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 349618 0 349674 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 352286 0 352342 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 355046 0 355102 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 357714 0 357770 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 360474 0 360530 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 363234 0 363290 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 365902 0 365958 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 369582 0 369638 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 372250 0 372306 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 375010 0 375066 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 377678 0 377734 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 380438 0 380494 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 383106 0 383162 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 385866 0 385922 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 388626 0 388682 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 391294 0 391350 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 394054 0 394110 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 396722 0 396778 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 399482 0 399538 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 402150 0 402206 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 404910 0 404966 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 407670 0 407726 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 410338 0 410394 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 413098 0 413154 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 415766 0 415822 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 418526 0 418582 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 421286 0 421342 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 127346 0 127402 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 423954 0 424010 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 426714 0 426770 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 429382 0 429438 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 432142 0 432198 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 434810 0 434866 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 437570 0 437626 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 440330 0 440386 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 442998 0 443054 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 130014 0 130070 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 146390 0 146446 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 160006 0 160062 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 165434 0 165490 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 168194 0 168250 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 173622 0 173678 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 176290 0 176346 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 181810 0 181866 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 184478 0 184534 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 187238 0 187294 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 192666 0 192722 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 195334 0 195390 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 198094 0 198150 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 200854 0 200910 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 203522 0 203578 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 206282 0 206338 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 208950 0 209006 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 211710 0 211766 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 214378 0 214434 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 217138 0 217194 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 222566 0 222622 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 225326 0 225382 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 227994 0 228050 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 230754 0 230810 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 233514 0 233570 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 236182 0 236238 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 238942 0 238998 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 241610 0 241666 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 244370 0 244426 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 247038 0 247094 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 249798 0 249854 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 252558 0 252614 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 255226 0 255282 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 257986 0 258042 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 260654 0 260710 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 263414 0 263470 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 266082 0 266138 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 268842 0 268898 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 271602 0 271658 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 274270 0 274326 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 277030 0 277086 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 279698 0 279754 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 282458 0 282514 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 285218 0 285274 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 287886 0 287942 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 290646 0 290702 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 293314 0 293370 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 296074 0 296130 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 298742 0 298798 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 301502 0 301558 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 304262 0 304318 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 306930 0 306986 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 309690 0 309746 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 312358 0 312414 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 315118 0 315174 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 317878 0 317934 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 320546 0 320602 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 323306 0 323362 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 325974 0 326030 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 328734 0 328790 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 331402 0 331458 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 334162 0 334218 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 336922 0 336978 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 339590 0 339646 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 342350 0 342406 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 345018 0 345074 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 347778 0 347834 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 350446 0 350502 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 353206 0 353262 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 355966 0 356022 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 358634 0 358690 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 361394 0 361450 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 364062 0 364118 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 366822 0 366878 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 370410 0 370466 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 373170 0 373226 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 375930 0 375986 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 378598 0 378654 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 381358 0 381414 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 384026 0 384082 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 386786 0 386842 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 389454 0 389510 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 392214 0 392270 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 394974 0 395030 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 397642 0 397698 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 400402 0 400458 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 403070 0 403126 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 405830 0 405886 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 408590 0 408646 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 411258 0 411314 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 414018 0 414074 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 416686 0 416742 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 419446 0 419502 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 422114 0 422170 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 424874 0 424930 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 427634 0 427690 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 430302 0 430358 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 433062 0 433118 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 435730 0 435786 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 438490 0 438546 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 441158 0 441214 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 443918 0 443974 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 179970 0 180026 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 193586 0 193642 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 196254 0 196310 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 199014 0 199070 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 201682 0 201738 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 204442 0 204498 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 212630 0 212686 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 215298 0 215354 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 223486 0 223542 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 226246 0 226302 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 228914 0 228970 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 231674 0 231730 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 234342 0 234398 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 237102 0 237158 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 239862 0 239918 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 242530 0 242586 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 245290 0 245346 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 250718 0 250774 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 256146 0 256202 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 258906 0 258962 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 261574 0 261630 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 264334 0 264390 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 267002 0 267058 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 269762 0 269818 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 272522 0 272578 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 275190 0 275246 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 277950 0 278006 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 280618 0 280674 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 283378 0 283434 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 286046 0 286102 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 288806 0 288862 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 294234 0 294290 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 299662 0 299718 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 302422 0 302478 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 305090 0 305146 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 310610 0 310666 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 313278 0 313334 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 316038 0 316094 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 318706 0 318762 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 321466 0 321522 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 324226 0 324282 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 326894 0 326950 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 329654 0 329710 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 332322 0 332378 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 335082 0 335138 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 337750 0 337806 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 340510 0 340566 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 343270 0 343326 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 345938 0 345994 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 348698 0 348754 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 351366 0 351422 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 354126 0 354182 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 356794 0 356850 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 359554 0 359610 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 362314 0 362370 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 364982 0 365038 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 367742 0 367798 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 434288 2128 434608 445040 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 445040 6 vssd1
port 503 nsew ground input
rlabel metal4 s 418928 2128 419248 445040 6 vssd1
port 503 nsew ground input
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 447200 447200
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 213557260
string GDS_START 1475556
<< end >>

