magic
tech sky130A
magscale 1 2
timestamp 1636386767
<< obsli1 >>
rect 1104 85 424551 424337
<< obsm1 >>
rect 382 8 424471 424516
<< metal2 >>
rect 1858 425904 1914 426704
rect 5538 425904 5594 426704
rect 9218 425904 9274 426704
rect 12990 425904 13046 426704
rect 16670 425904 16726 426704
rect 20442 425904 20498 426704
rect 24122 425904 24178 426704
rect 27894 425904 27950 426704
rect 31574 425904 31630 426704
rect 35346 425904 35402 426704
rect 39026 425904 39082 426704
rect 42798 425904 42854 426704
rect 46478 425904 46534 426704
rect 50250 425904 50306 426704
rect 53930 425904 53986 426704
rect 57702 425904 57758 426704
rect 61382 425904 61438 426704
rect 65154 425904 65210 426704
rect 68834 425904 68890 426704
rect 72606 425904 72662 426704
rect 76286 425904 76342 426704
rect 80058 425904 80114 426704
rect 83738 425904 83794 426704
rect 87510 425904 87566 426704
rect 91190 425904 91246 426704
rect 94962 425904 95018 426704
rect 98642 425904 98698 426704
rect 102414 425904 102470 426704
rect 106094 425904 106150 426704
rect 109774 425904 109830 426704
rect 113546 425904 113602 426704
rect 117226 425904 117282 426704
rect 120998 425904 121054 426704
rect 124678 425904 124734 426704
rect 128450 425904 128506 426704
rect 132130 425904 132186 426704
rect 135902 425904 135958 426704
rect 139582 425904 139638 426704
rect 143354 425904 143410 426704
rect 147034 425904 147090 426704
rect 150806 425904 150862 426704
rect 154486 425904 154542 426704
rect 158258 425904 158314 426704
rect 161938 425904 161994 426704
rect 165710 425904 165766 426704
rect 169390 425904 169446 426704
rect 173162 425904 173218 426704
rect 176842 425904 176898 426704
rect 180614 425904 180670 426704
rect 184294 425904 184350 426704
rect 188066 425904 188122 426704
rect 191746 425904 191802 426704
rect 195518 425904 195574 426704
rect 199198 425904 199254 426704
rect 202970 425904 203026 426704
rect 206650 425904 206706 426704
rect 210422 425904 210478 426704
rect 214102 425904 214158 426704
rect 217782 425904 217838 426704
rect 221554 425904 221610 426704
rect 225234 425904 225290 426704
rect 229006 425904 229062 426704
rect 232686 425904 232742 426704
rect 236458 425904 236514 426704
rect 240138 425904 240194 426704
rect 243910 425904 243966 426704
rect 247590 425904 247646 426704
rect 251362 425904 251418 426704
rect 255042 425904 255098 426704
rect 258814 425904 258870 426704
rect 262494 425904 262550 426704
rect 266266 425904 266322 426704
rect 269946 425904 270002 426704
rect 273718 425904 273774 426704
rect 277398 425904 277454 426704
rect 281170 425904 281226 426704
rect 284850 425904 284906 426704
rect 288622 425904 288678 426704
rect 292302 425904 292358 426704
rect 296074 425904 296130 426704
rect 299754 425904 299810 426704
rect 303526 425904 303582 426704
rect 307206 425904 307262 426704
rect 310978 425904 311034 426704
rect 314658 425904 314714 426704
rect 318430 425904 318486 426704
rect 322110 425904 322166 426704
rect 325790 425904 325846 426704
rect 329562 425904 329618 426704
rect 333242 425904 333298 426704
rect 337014 425904 337070 426704
rect 340694 425904 340750 426704
rect 344466 425904 344522 426704
rect 348146 425904 348202 426704
rect 351918 425904 351974 426704
rect 355598 425904 355654 426704
rect 359370 425904 359426 426704
rect 363050 425904 363106 426704
rect 366822 425904 366878 426704
rect 370502 425904 370558 426704
rect 374274 425904 374330 426704
rect 377954 425904 378010 426704
rect 381726 425904 381782 426704
rect 385406 425904 385462 426704
rect 389178 425904 389234 426704
rect 392858 425904 392914 426704
rect 396630 425904 396686 426704
rect 400310 425904 400366 426704
rect 404082 425904 404138 426704
rect 407762 425904 407818 426704
rect 411534 425904 411590 426704
rect 415214 425904 415270 426704
rect 418986 425904 419042 426704
rect 422666 425904 422722 426704
rect 386 0 442 800
rect 1214 0 1270 800
rect 2042 0 2098 800
rect 2962 0 3018 800
rect 3790 0 3846 800
rect 4618 0 4674 800
rect 5538 0 5594 800
rect 6366 0 6422 800
rect 7194 0 7250 800
rect 8114 0 8170 800
rect 8942 0 8998 800
rect 9770 0 9826 800
rect 10690 0 10746 800
rect 11518 0 11574 800
rect 12438 0 12494 800
rect 13266 0 13322 800
rect 14094 0 14150 800
rect 15014 0 15070 800
rect 15842 0 15898 800
rect 16670 0 16726 800
rect 17590 0 17646 800
rect 18418 0 18474 800
rect 19246 0 19302 800
rect 20166 0 20222 800
rect 20994 0 21050 800
rect 21914 0 21970 800
rect 22742 0 22798 800
rect 23570 0 23626 800
rect 24490 0 24546 800
rect 25318 0 25374 800
rect 26146 0 26202 800
rect 27066 0 27122 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29642 0 29698 800
rect 30470 0 30526 800
rect 31298 0 31354 800
rect 32218 0 32274 800
rect 33046 0 33102 800
rect 33966 0 34022 800
rect 34794 0 34850 800
rect 35622 0 35678 800
rect 36542 0 36598 800
rect 37370 0 37426 800
rect 38198 0 38254 800
rect 39118 0 39174 800
rect 39946 0 40002 800
rect 40774 0 40830 800
rect 41694 0 41750 800
rect 42522 0 42578 800
rect 43442 0 43498 800
rect 44270 0 44326 800
rect 45098 0 45154 800
rect 46018 0 46074 800
rect 46846 0 46902 800
rect 47674 0 47730 800
rect 48594 0 48650 800
rect 49422 0 49478 800
rect 50250 0 50306 800
rect 51170 0 51226 800
rect 51998 0 52054 800
rect 52918 0 52974 800
rect 53746 0 53802 800
rect 54574 0 54630 800
rect 55494 0 55550 800
rect 56322 0 56378 800
rect 57150 0 57206 800
rect 58070 0 58126 800
rect 58898 0 58954 800
rect 59726 0 59782 800
rect 60646 0 60702 800
rect 61474 0 61530 800
rect 62302 0 62358 800
rect 63222 0 63278 800
rect 64050 0 64106 800
rect 64970 0 65026 800
rect 65798 0 65854 800
rect 66626 0 66682 800
rect 67546 0 67602 800
rect 68374 0 68430 800
rect 69202 0 69258 800
rect 70122 0 70178 800
rect 70950 0 71006 800
rect 71778 0 71834 800
rect 72698 0 72754 800
rect 73526 0 73582 800
rect 74446 0 74502 800
rect 75274 0 75330 800
rect 76102 0 76158 800
rect 77022 0 77078 800
rect 77850 0 77906 800
rect 78678 0 78734 800
rect 79598 0 79654 800
rect 80426 0 80482 800
rect 81254 0 81310 800
rect 82174 0 82230 800
rect 83002 0 83058 800
rect 83922 0 83978 800
rect 84750 0 84806 800
rect 85578 0 85634 800
rect 86498 0 86554 800
rect 87326 0 87382 800
rect 88154 0 88210 800
rect 89074 0 89130 800
rect 89902 0 89958 800
rect 90730 0 90786 800
rect 91650 0 91706 800
rect 92478 0 92534 800
rect 93306 0 93362 800
rect 94226 0 94282 800
rect 95054 0 95110 800
rect 95974 0 96030 800
rect 96802 0 96858 800
rect 97630 0 97686 800
rect 98550 0 98606 800
rect 99378 0 99434 800
rect 100206 0 100262 800
rect 101126 0 101182 800
rect 101954 0 102010 800
rect 102782 0 102838 800
rect 103702 0 103758 800
rect 104530 0 104586 800
rect 105450 0 105506 800
rect 106278 0 106334 800
rect 107106 0 107162 800
rect 108026 0 108082 800
rect 108854 0 108910 800
rect 109682 0 109738 800
rect 110602 0 110658 800
rect 111430 0 111486 800
rect 112258 0 112314 800
rect 113178 0 113234 800
rect 114006 0 114062 800
rect 114926 0 114982 800
rect 115754 0 115810 800
rect 116582 0 116638 800
rect 117502 0 117558 800
rect 118330 0 118386 800
rect 119158 0 119214 800
rect 120078 0 120134 800
rect 120906 0 120962 800
rect 121734 0 121790 800
rect 122654 0 122710 800
rect 123482 0 123538 800
rect 124310 0 124366 800
rect 125230 0 125286 800
rect 126058 0 126114 800
rect 126978 0 127034 800
rect 127806 0 127862 800
rect 128634 0 128690 800
rect 129554 0 129610 800
rect 130382 0 130438 800
rect 131210 0 131266 800
rect 132130 0 132186 800
rect 132958 0 133014 800
rect 133786 0 133842 800
rect 134706 0 134762 800
rect 135534 0 135590 800
rect 136454 0 136510 800
rect 137282 0 137338 800
rect 138110 0 138166 800
rect 139030 0 139086 800
rect 139858 0 139914 800
rect 140686 0 140742 800
rect 141606 0 141662 800
rect 142434 0 142490 800
rect 143262 0 143318 800
rect 144182 0 144238 800
rect 145010 0 145066 800
rect 145930 0 145986 800
rect 146758 0 146814 800
rect 147586 0 147642 800
rect 148506 0 148562 800
rect 149334 0 149390 800
rect 150162 0 150218 800
rect 151082 0 151138 800
rect 151910 0 151966 800
rect 152738 0 152794 800
rect 153658 0 153714 800
rect 154486 0 154542 800
rect 155314 0 155370 800
rect 156234 0 156290 800
rect 157062 0 157118 800
rect 157982 0 158038 800
rect 158810 0 158866 800
rect 159638 0 159694 800
rect 160558 0 160614 800
rect 161386 0 161442 800
rect 162214 0 162270 800
rect 163134 0 163190 800
rect 163962 0 164018 800
rect 164790 0 164846 800
rect 165710 0 165766 800
rect 166538 0 166594 800
rect 167458 0 167514 800
rect 168286 0 168342 800
rect 169114 0 169170 800
rect 170034 0 170090 800
rect 170862 0 170918 800
rect 171690 0 171746 800
rect 172610 0 172666 800
rect 173438 0 173494 800
rect 174266 0 174322 800
rect 175186 0 175242 800
rect 176014 0 176070 800
rect 176934 0 176990 800
rect 177762 0 177818 800
rect 178590 0 178646 800
rect 179510 0 179566 800
rect 180338 0 180394 800
rect 181166 0 181222 800
rect 182086 0 182142 800
rect 182914 0 182970 800
rect 183742 0 183798 800
rect 184662 0 184718 800
rect 185490 0 185546 800
rect 186318 0 186374 800
rect 187238 0 187294 800
rect 188066 0 188122 800
rect 188986 0 189042 800
rect 189814 0 189870 800
rect 190642 0 190698 800
rect 191562 0 191618 800
rect 192390 0 192446 800
rect 193218 0 193274 800
rect 194138 0 194194 800
rect 194966 0 195022 800
rect 195794 0 195850 800
rect 196714 0 196770 800
rect 197542 0 197598 800
rect 198462 0 198518 800
rect 199290 0 199346 800
rect 200118 0 200174 800
rect 201038 0 201094 800
rect 201866 0 201922 800
rect 202694 0 202750 800
rect 203614 0 203670 800
rect 204442 0 204498 800
rect 205270 0 205326 800
rect 206190 0 206246 800
rect 207018 0 207074 800
rect 207938 0 207994 800
rect 208766 0 208822 800
rect 209594 0 209650 800
rect 210514 0 210570 800
rect 211342 0 211398 800
rect 212170 0 212226 800
rect 213090 0 213146 800
rect 213918 0 213974 800
rect 214746 0 214802 800
rect 215666 0 215722 800
rect 216494 0 216550 800
rect 217322 0 217378 800
rect 218242 0 218298 800
rect 219070 0 219126 800
rect 219990 0 220046 800
rect 220818 0 220874 800
rect 221646 0 221702 800
rect 222566 0 222622 800
rect 223394 0 223450 800
rect 224222 0 224278 800
rect 225142 0 225198 800
rect 225970 0 226026 800
rect 226798 0 226854 800
rect 227718 0 227774 800
rect 228546 0 228602 800
rect 229466 0 229522 800
rect 230294 0 230350 800
rect 231122 0 231178 800
rect 232042 0 232098 800
rect 232870 0 232926 800
rect 233698 0 233754 800
rect 234618 0 234674 800
rect 235446 0 235502 800
rect 236274 0 236330 800
rect 237194 0 237250 800
rect 238022 0 238078 800
rect 238942 0 238998 800
rect 239770 0 239826 800
rect 240598 0 240654 800
rect 241518 0 241574 800
rect 242346 0 242402 800
rect 243174 0 243230 800
rect 244094 0 244150 800
rect 244922 0 244978 800
rect 245750 0 245806 800
rect 246670 0 246726 800
rect 247498 0 247554 800
rect 248326 0 248382 800
rect 249246 0 249302 800
rect 250074 0 250130 800
rect 250994 0 251050 800
rect 251822 0 251878 800
rect 252650 0 252706 800
rect 253570 0 253626 800
rect 254398 0 254454 800
rect 255226 0 255282 800
rect 256146 0 256202 800
rect 256974 0 257030 800
rect 257802 0 257858 800
rect 258722 0 258778 800
rect 259550 0 259606 800
rect 260470 0 260526 800
rect 261298 0 261354 800
rect 262126 0 262182 800
rect 263046 0 263102 800
rect 263874 0 263930 800
rect 264702 0 264758 800
rect 265622 0 265678 800
rect 266450 0 266506 800
rect 267278 0 267334 800
rect 268198 0 268254 800
rect 269026 0 269082 800
rect 269946 0 270002 800
rect 270774 0 270830 800
rect 271602 0 271658 800
rect 272522 0 272578 800
rect 273350 0 273406 800
rect 274178 0 274234 800
rect 275098 0 275154 800
rect 275926 0 275982 800
rect 276754 0 276810 800
rect 277674 0 277730 800
rect 278502 0 278558 800
rect 279330 0 279386 800
rect 280250 0 280306 800
rect 281078 0 281134 800
rect 281998 0 282054 800
rect 282826 0 282882 800
rect 283654 0 283710 800
rect 284574 0 284630 800
rect 285402 0 285458 800
rect 286230 0 286286 800
rect 287150 0 287206 800
rect 287978 0 288034 800
rect 288806 0 288862 800
rect 289726 0 289782 800
rect 290554 0 290610 800
rect 291474 0 291530 800
rect 292302 0 292358 800
rect 293130 0 293186 800
rect 294050 0 294106 800
rect 294878 0 294934 800
rect 295706 0 295762 800
rect 296626 0 296682 800
rect 297454 0 297510 800
rect 298282 0 298338 800
rect 299202 0 299258 800
rect 300030 0 300086 800
rect 300950 0 301006 800
rect 301778 0 301834 800
rect 302606 0 302662 800
rect 303526 0 303582 800
rect 304354 0 304410 800
rect 305182 0 305238 800
rect 306102 0 306158 800
rect 306930 0 306986 800
rect 307758 0 307814 800
rect 308678 0 308734 800
rect 309506 0 309562 800
rect 310334 0 310390 800
rect 311254 0 311310 800
rect 312082 0 312138 800
rect 313002 0 313058 800
rect 313830 0 313886 800
rect 314658 0 314714 800
rect 315578 0 315634 800
rect 316406 0 316462 800
rect 317234 0 317290 800
rect 318154 0 318210 800
rect 318982 0 319038 800
rect 319810 0 319866 800
rect 320730 0 320786 800
rect 321558 0 321614 800
rect 322478 0 322534 800
rect 323306 0 323362 800
rect 324134 0 324190 800
rect 325054 0 325110 800
rect 325882 0 325938 800
rect 326710 0 326766 800
rect 327630 0 327686 800
rect 328458 0 328514 800
rect 329286 0 329342 800
rect 330206 0 330262 800
rect 331034 0 331090 800
rect 331954 0 332010 800
rect 332782 0 332838 800
rect 333610 0 333666 800
rect 334530 0 334586 800
rect 335358 0 335414 800
rect 336186 0 336242 800
rect 337106 0 337162 800
rect 337934 0 337990 800
rect 338762 0 338818 800
rect 339682 0 339738 800
rect 340510 0 340566 800
rect 341338 0 341394 800
rect 342258 0 342314 800
rect 343086 0 343142 800
rect 344006 0 344062 800
rect 344834 0 344890 800
rect 345662 0 345718 800
rect 346582 0 346638 800
rect 347410 0 347466 800
rect 348238 0 348294 800
rect 349158 0 349214 800
rect 349986 0 350042 800
rect 350814 0 350870 800
rect 351734 0 351790 800
rect 352562 0 352618 800
rect 353482 0 353538 800
rect 354310 0 354366 800
rect 355138 0 355194 800
rect 356058 0 356114 800
rect 356886 0 356942 800
rect 357714 0 357770 800
rect 358634 0 358690 800
rect 359462 0 359518 800
rect 360290 0 360346 800
rect 361210 0 361266 800
rect 362038 0 362094 800
rect 362958 0 363014 800
rect 363786 0 363842 800
rect 364614 0 364670 800
rect 365534 0 365590 800
rect 366362 0 366418 800
rect 367190 0 367246 800
rect 368110 0 368166 800
rect 368938 0 368994 800
rect 369766 0 369822 800
rect 370686 0 370742 800
rect 371514 0 371570 800
rect 372342 0 372398 800
rect 373262 0 373318 800
rect 374090 0 374146 800
rect 375010 0 375066 800
rect 375838 0 375894 800
rect 376666 0 376722 800
rect 377586 0 377642 800
rect 378414 0 378470 800
rect 379242 0 379298 800
rect 380162 0 380218 800
rect 380990 0 381046 800
rect 381818 0 381874 800
rect 382738 0 382794 800
rect 383566 0 383622 800
rect 384486 0 384542 800
rect 385314 0 385370 800
rect 386142 0 386198 800
rect 387062 0 387118 800
rect 387890 0 387946 800
rect 388718 0 388774 800
rect 389638 0 389694 800
rect 390466 0 390522 800
rect 391294 0 391350 800
rect 392214 0 392270 800
rect 393042 0 393098 800
rect 393962 0 394018 800
rect 394790 0 394846 800
rect 395618 0 395674 800
rect 396538 0 396594 800
rect 397366 0 397422 800
rect 398194 0 398250 800
rect 399114 0 399170 800
rect 399942 0 399998 800
rect 400770 0 400826 800
rect 401690 0 401746 800
rect 402518 0 402574 800
rect 403346 0 403402 800
rect 404266 0 404322 800
rect 405094 0 405150 800
rect 406014 0 406070 800
rect 406842 0 406898 800
rect 407670 0 407726 800
rect 408590 0 408646 800
rect 409418 0 409474 800
rect 410246 0 410302 800
rect 411166 0 411222 800
rect 411994 0 412050 800
rect 412822 0 412878 800
rect 413742 0 413798 800
rect 414570 0 414626 800
rect 415490 0 415546 800
rect 416318 0 416374 800
rect 417146 0 417202 800
rect 418066 0 418122 800
rect 418894 0 418950 800
rect 419722 0 419778 800
rect 420642 0 420698 800
rect 421470 0 421526 800
rect 422298 0 422354 800
rect 423218 0 423274 800
rect 424046 0 424102 800
<< obsm2 >>
rect 388 425848 1802 425904
rect 1970 425848 5482 425904
rect 5650 425848 9162 425904
rect 9330 425848 12934 425904
rect 13102 425848 16614 425904
rect 16782 425848 20386 425904
rect 20554 425848 24066 425904
rect 24234 425848 27838 425904
rect 28006 425848 31518 425904
rect 31686 425848 35290 425904
rect 35458 425848 38970 425904
rect 39138 425848 42742 425904
rect 42910 425848 46422 425904
rect 46590 425848 50194 425904
rect 50362 425848 53874 425904
rect 54042 425848 57646 425904
rect 57814 425848 61326 425904
rect 61494 425848 65098 425904
rect 65266 425848 68778 425904
rect 68946 425848 72550 425904
rect 72718 425848 76230 425904
rect 76398 425848 80002 425904
rect 80170 425848 83682 425904
rect 83850 425848 87454 425904
rect 87622 425848 91134 425904
rect 91302 425848 94906 425904
rect 95074 425848 98586 425904
rect 98754 425848 102358 425904
rect 102526 425848 106038 425904
rect 106206 425848 109718 425904
rect 109886 425848 113490 425904
rect 113658 425848 117170 425904
rect 117338 425848 120942 425904
rect 121110 425848 124622 425904
rect 124790 425848 128394 425904
rect 128562 425848 132074 425904
rect 132242 425848 135846 425904
rect 136014 425848 139526 425904
rect 139694 425848 143298 425904
rect 143466 425848 146978 425904
rect 147146 425848 150750 425904
rect 150918 425848 154430 425904
rect 154598 425848 158202 425904
rect 158370 425848 161882 425904
rect 162050 425848 165654 425904
rect 165822 425848 169334 425904
rect 169502 425848 173106 425904
rect 173274 425848 176786 425904
rect 176954 425848 180558 425904
rect 180726 425848 184238 425904
rect 184406 425848 188010 425904
rect 188178 425848 191690 425904
rect 191858 425848 195462 425904
rect 195630 425848 199142 425904
rect 199310 425848 202914 425904
rect 203082 425848 206594 425904
rect 206762 425848 210366 425904
rect 210534 425848 214046 425904
rect 214214 425848 217726 425904
rect 217894 425848 221498 425904
rect 221666 425848 225178 425904
rect 225346 425848 228950 425904
rect 229118 425848 232630 425904
rect 232798 425848 236402 425904
rect 236570 425848 240082 425904
rect 240250 425848 243854 425904
rect 244022 425848 247534 425904
rect 247702 425848 251306 425904
rect 251474 425848 254986 425904
rect 255154 425848 258758 425904
rect 258926 425848 262438 425904
rect 262606 425848 266210 425904
rect 266378 425848 269890 425904
rect 270058 425848 273662 425904
rect 273830 425848 277342 425904
rect 277510 425848 281114 425904
rect 281282 425848 284794 425904
rect 284962 425848 288566 425904
rect 288734 425848 292246 425904
rect 292414 425848 296018 425904
rect 296186 425848 299698 425904
rect 299866 425848 303470 425904
rect 303638 425848 307150 425904
rect 307318 425848 310922 425904
rect 311090 425848 314602 425904
rect 314770 425848 318374 425904
rect 318542 425848 322054 425904
rect 322222 425848 325734 425904
rect 325902 425848 329506 425904
rect 329674 425848 333186 425904
rect 333354 425848 336958 425904
rect 337126 425848 340638 425904
rect 340806 425848 344410 425904
rect 344578 425848 348090 425904
rect 348258 425848 351862 425904
rect 352030 425848 355542 425904
rect 355710 425848 359314 425904
rect 359482 425848 362994 425904
rect 363162 425848 366766 425904
rect 366934 425848 370446 425904
rect 370614 425848 374218 425904
rect 374386 425848 377898 425904
rect 378066 425848 381670 425904
rect 381838 425848 385350 425904
rect 385518 425848 389122 425904
rect 389290 425848 392802 425904
rect 392970 425848 396574 425904
rect 396742 425848 400254 425904
rect 400422 425848 404026 425904
rect 404194 425848 407706 425904
rect 407874 425848 411478 425904
rect 411646 425848 415158 425904
rect 415326 425848 418930 425904
rect 419098 425848 422610 425904
rect 422778 425848 424378 425904
rect 388 856 424378 425848
rect 498 2 1158 856
rect 1326 2 1986 856
rect 2154 2 2906 856
rect 3074 2 3734 856
rect 3902 2 4562 856
rect 4730 2 5482 856
rect 5650 2 6310 856
rect 6478 2 7138 856
rect 7306 2 8058 856
rect 8226 2 8886 856
rect 9054 2 9714 856
rect 9882 2 10634 856
rect 10802 2 11462 856
rect 11630 2 12382 856
rect 12550 2 13210 856
rect 13378 2 14038 856
rect 14206 2 14958 856
rect 15126 2 15786 856
rect 15954 2 16614 856
rect 16782 2 17534 856
rect 17702 2 18362 856
rect 18530 2 19190 856
rect 19358 2 20110 856
rect 20278 2 20938 856
rect 21106 2 21858 856
rect 22026 2 22686 856
rect 22854 2 23514 856
rect 23682 2 24434 856
rect 24602 2 25262 856
rect 25430 2 26090 856
rect 26258 2 27010 856
rect 27178 2 27838 856
rect 28006 2 28666 856
rect 28834 2 29586 856
rect 29754 2 30414 856
rect 30582 2 31242 856
rect 31410 2 32162 856
rect 32330 2 32990 856
rect 33158 2 33910 856
rect 34078 2 34738 856
rect 34906 2 35566 856
rect 35734 2 36486 856
rect 36654 2 37314 856
rect 37482 2 38142 856
rect 38310 2 39062 856
rect 39230 2 39890 856
rect 40058 2 40718 856
rect 40886 2 41638 856
rect 41806 2 42466 856
rect 42634 2 43386 856
rect 43554 2 44214 856
rect 44382 2 45042 856
rect 45210 2 45962 856
rect 46130 2 46790 856
rect 46958 2 47618 856
rect 47786 2 48538 856
rect 48706 2 49366 856
rect 49534 2 50194 856
rect 50362 2 51114 856
rect 51282 2 51942 856
rect 52110 2 52862 856
rect 53030 2 53690 856
rect 53858 2 54518 856
rect 54686 2 55438 856
rect 55606 2 56266 856
rect 56434 2 57094 856
rect 57262 2 58014 856
rect 58182 2 58842 856
rect 59010 2 59670 856
rect 59838 2 60590 856
rect 60758 2 61418 856
rect 61586 2 62246 856
rect 62414 2 63166 856
rect 63334 2 63994 856
rect 64162 2 64914 856
rect 65082 2 65742 856
rect 65910 2 66570 856
rect 66738 2 67490 856
rect 67658 2 68318 856
rect 68486 2 69146 856
rect 69314 2 70066 856
rect 70234 2 70894 856
rect 71062 2 71722 856
rect 71890 2 72642 856
rect 72810 2 73470 856
rect 73638 2 74390 856
rect 74558 2 75218 856
rect 75386 2 76046 856
rect 76214 2 76966 856
rect 77134 2 77794 856
rect 77962 2 78622 856
rect 78790 2 79542 856
rect 79710 2 80370 856
rect 80538 2 81198 856
rect 81366 2 82118 856
rect 82286 2 82946 856
rect 83114 2 83866 856
rect 84034 2 84694 856
rect 84862 2 85522 856
rect 85690 2 86442 856
rect 86610 2 87270 856
rect 87438 2 88098 856
rect 88266 2 89018 856
rect 89186 2 89846 856
rect 90014 2 90674 856
rect 90842 2 91594 856
rect 91762 2 92422 856
rect 92590 2 93250 856
rect 93418 2 94170 856
rect 94338 2 94998 856
rect 95166 2 95918 856
rect 96086 2 96746 856
rect 96914 2 97574 856
rect 97742 2 98494 856
rect 98662 2 99322 856
rect 99490 2 100150 856
rect 100318 2 101070 856
rect 101238 2 101898 856
rect 102066 2 102726 856
rect 102894 2 103646 856
rect 103814 2 104474 856
rect 104642 2 105394 856
rect 105562 2 106222 856
rect 106390 2 107050 856
rect 107218 2 107970 856
rect 108138 2 108798 856
rect 108966 2 109626 856
rect 109794 2 110546 856
rect 110714 2 111374 856
rect 111542 2 112202 856
rect 112370 2 113122 856
rect 113290 2 113950 856
rect 114118 2 114870 856
rect 115038 2 115698 856
rect 115866 2 116526 856
rect 116694 2 117446 856
rect 117614 2 118274 856
rect 118442 2 119102 856
rect 119270 2 120022 856
rect 120190 2 120850 856
rect 121018 2 121678 856
rect 121846 2 122598 856
rect 122766 2 123426 856
rect 123594 2 124254 856
rect 124422 2 125174 856
rect 125342 2 126002 856
rect 126170 2 126922 856
rect 127090 2 127750 856
rect 127918 2 128578 856
rect 128746 2 129498 856
rect 129666 2 130326 856
rect 130494 2 131154 856
rect 131322 2 132074 856
rect 132242 2 132902 856
rect 133070 2 133730 856
rect 133898 2 134650 856
rect 134818 2 135478 856
rect 135646 2 136398 856
rect 136566 2 137226 856
rect 137394 2 138054 856
rect 138222 2 138974 856
rect 139142 2 139802 856
rect 139970 2 140630 856
rect 140798 2 141550 856
rect 141718 2 142378 856
rect 142546 2 143206 856
rect 143374 2 144126 856
rect 144294 2 144954 856
rect 145122 2 145874 856
rect 146042 2 146702 856
rect 146870 2 147530 856
rect 147698 2 148450 856
rect 148618 2 149278 856
rect 149446 2 150106 856
rect 150274 2 151026 856
rect 151194 2 151854 856
rect 152022 2 152682 856
rect 152850 2 153602 856
rect 153770 2 154430 856
rect 154598 2 155258 856
rect 155426 2 156178 856
rect 156346 2 157006 856
rect 157174 2 157926 856
rect 158094 2 158754 856
rect 158922 2 159582 856
rect 159750 2 160502 856
rect 160670 2 161330 856
rect 161498 2 162158 856
rect 162326 2 163078 856
rect 163246 2 163906 856
rect 164074 2 164734 856
rect 164902 2 165654 856
rect 165822 2 166482 856
rect 166650 2 167402 856
rect 167570 2 168230 856
rect 168398 2 169058 856
rect 169226 2 169978 856
rect 170146 2 170806 856
rect 170974 2 171634 856
rect 171802 2 172554 856
rect 172722 2 173382 856
rect 173550 2 174210 856
rect 174378 2 175130 856
rect 175298 2 175958 856
rect 176126 2 176878 856
rect 177046 2 177706 856
rect 177874 2 178534 856
rect 178702 2 179454 856
rect 179622 2 180282 856
rect 180450 2 181110 856
rect 181278 2 182030 856
rect 182198 2 182858 856
rect 183026 2 183686 856
rect 183854 2 184606 856
rect 184774 2 185434 856
rect 185602 2 186262 856
rect 186430 2 187182 856
rect 187350 2 188010 856
rect 188178 2 188930 856
rect 189098 2 189758 856
rect 189926 2 190586 856
rect 190754 2 191506 856
rect 191674 2 192334 856
rect 192502 2 193162 856
rect 193330 2 194082 856
rect 194250 2 194910 856
rect 195078 2 195738 856
rect 195906 2 196658 856
rect 196826 2 197486 856
rect 197654 2 198406 856
rect 198574 2 199234 856
rect 199402 2 200062 856
rect 200230 2 200982 856
rect 201150 2 201810 856
rect 201978 2 202638 856
rect 202806 2 203558 856
rect 203726 2 204386 856
rect 204554 2 205214 856
rect 205382 2 206134 856
rect 206302 2 206962 856
rect 207130 2 207882 856
rect 208050 2 208710 856
rect 208878 2 209538 856
rect 209706 2 210458 856
rect 210626 2 211286 856
rect 211454 2 212114 856
rect 212282 2 213034 856
rect 213202 2 213862 856
rect 214030 2 214690 856
rect 214858 2 215610 856
rect 215778 2 216438 856
rect 216606 2 217266 856
rect 217434 2 218186 856
rect 218354 2 219014 856
rect 219182 2 219934 856
rect 220102 2 220762 856
rect 220930 2 221590 856
rect 221758 2 222510 856
rect 222678 2 223338 856
rect 223506 2 224166 856
rect 224334 2 225086 856
rect 225254 2 225914 856
rect 226082 2 226742 856
rect 226910 2 227662 856
rect 227830 2 228490 856
rect 228658 2 229410 856
rect 229578 2 230238 856
rect 230406 2 231066 856
rect 231234 2 231986 856
rect 232154 2 232814 856
rect 232982 2 233642 856
rect 233810 2 234562 856
rect 234730 2 235390 856
rect 235558 2 236218 856
rect 236386 2 237138 856
rect 237306 2 237966 856
rect 238134 2 238886 856
rect 239054 2 239714 856
rect 239882 2 240542 856
rect 240710 2 241462 856
rect 241630 2 242290 856
rect 242458 2 243118 856
rect 243286 2 244038 856
rect 244206 2 244866 856
rect 245034 2 245694 856
rect 245862 2 246614 856
rect 246782 2 247442 856
rect 247610 2 248270 856
rect 248438 2 249190 856
rect 249358 2 250018 856
rect 250186 2 250938 856
rect 251106 2 251766 856
rect 251934 2 252594 856
rect 252762 2 253514 856
rect 253682 2 254342 856
rect 254510 2 255170 856
rect 255338 2 256090 856
rect 256258 2 256918 856
rect 257086 2 257746 856
rect 257914 2 258666 856
rect 258834 2 259494 856
rect 259662 2 260414 856
rect 260582 2 261242 856
rect 261410 2 262070 856
rect 262238 2 262990 856
rect 263158 2 263818 856
rect 263986 2 264646 856
rect 264814 2 265566 856
rect 265734 2 266394 856
rect 266562 2 267222 856
rect 267390 2 268142 856
rect 268310 2 268970 856
rect 269138 2 269890 856
rect 270058 2 270718 856
rect 270886 2 271546 856
rect 271714 2 272466 856
rect 272634 2 273294 856
rect 273462 2 274122 856
rect 274290 2 275042 856
rect 275210 2 275870 856
rect 276038 2 276698 856
rect 276866 2 277618 856
rect 277786 2 278446 856
rect 278614 2 279274 856
rect 279442 2 280194 856
rect 280362 2 281022 856
rect 281190 2 281942 856
rect 282110 2 282770 856
rect 282938 2 283598 856
rect 283766 2 284518 856
rect 284686 2 285346 856
rect 285514 2 286174 856
rect 286342 2 287094 856
rect 287262 2 287922 856
rect 288090 2 288750 856
rect 288918 2 289670 856
rect 289838 2 290498 856
rect 290666 2 291418 856
rect 291586 2 292246 856
rect 292414 2 293074 856
rect 293242 2 293994 856
rect 294162 2 294822 856
rect 294990 2 295650 856
rect 295818 2 296570 856
rect 296738 2 297398 856
rect 297566 2 298226 856
rect 298394 2 299146 856
rect 299314 2 299974 856
rect 300142 2 300894 856
rect 301062 2 301722 856
rect 301890 2 302550 856
rect 302718 2 303470 856
rect 303638 2 304298 856
rect 304466 2 305126 856
rect 305294 2 306046 856
rect 306214 2 306874 856
rect 307042 2 307702 856
rect 307870 2 308622 856
rect 308790 2 309450 856
rect 309618 2 310278 856
rect 310446 2 311198 856
rect 311366 2 312026 856
rect 312194 2 312946 856
rect 313114 2 313774 856
rect 313942 2 314602 856
rect 314770 2 315522 856
rect 315690 2 316350 856
rect 316518 2 317178 856
rect 317346 2 318098 856
rect 318266 2 318926 856
rect 319094 2 319754 856
rect 319922 2 320674 856
rect 320842 2 321502 856
rect 321670 2 322422 856
rect 322590 2 323250 856
rect 323418 2 324078 856
rect 324246 2 324998 856
rect 325166 2 325826 856
rect 325994 2 326654 856
rect 326822 2 327574 856
rect 327742 2 328402 856
rect 328570 2 329230 856
rect 329398 2 330150 856
rect 330318 2 330978 856
rect 331146 2 331898 856
rect 332066 2 332726 856
rect 332894 2 333554 856
rect 333722 2 334474 856
rect 334642 2 335302 856
rect 335470 2 336130 856
rect 336298 2 337050 856
rect 337218 2 337878 856
rect 338046 2 338706 856
rect 338874 2 339626 856
rect 339794 2 340454 856
rect 340622 2 341282 856
rect 341450 2 342202 856
rect 342370 2 343030 856
rect 343198 2 343950 856
rect 344118 2 344778 856
rect 344946 2 345606 856
rect 345774 2 346526 856
rect 346694 2 347354 856
rect 347522 2 348182 856
rect 348350 2 349102 856
rect 349270 2 349930 856
rect 350098 2 350758 856
rect 350926 2 351678 856
rect 351846 2 352506 856
rect 352674 2 353426 856
rect 353594 2 354254 856
rect 354422 2 355082 856
rect 355250 2 356002 856
rect 356170 2 356830 856
rect 356998 2 357658 856
rect 357826 2 358578 856
rect 358746 2 359406 856
rect 359574 2 360234 856
rect 360402 2 361154 856
rect 361322 2 361982 856
rect 362150 2 362902 856
rect 363070 2 363730 856
rect 363898 2 364558 856
rect 364726 2 365478 856
rect 365646 2 366306 856
rect 366474 2 367134 856
rect 367302 2 368054 856
rect 368222 2 368882 856
rect 369050 2 369710 856
rect 369878 2 370630 856
rect 370798 2 371458 856
rect 371626 2 372286 856
rect 372454 2 373206 856
rect 373374 2 374034 856
rect 374202 2 374954 856
rect 375122 2 375782 856
rect 375950 2 376610 856
rect 376778 2 377530 856
rect 377698 2 378358 856
rect 378526 2 379186 856
rect 379354 2 380106 856
rect 380274 2 380934 856
rect 381102 2 381762 856
rect 381930 2 382682 856
rect 382850 2 383510 856
rect 383678 2 384430 856
rect 384598 2 385258 856
rect 385426 2 386086 856
rect 386254 2 387006 856
rect 387174 2 387834 856
rect 388002 2 388662 856
rect 388830 2 389582 856
rect 389750 2 390410 856
rect 390578 2 391238 856
rect 391406 2 392158 856
rect 392326 2 392986 856
rect 393154 2 393906 856
rect 394074 2 394734 856
rect 394902 2 395562 856
rect 395730 2 396482 856
rect 396650 2 397310 856
rect 397478 2 398138 856
rect 398306 2 399058 856
rect 399226 2 399886 856
rect 400054 2 400714 856
rect 400882 2 401634 856
rect 401802 2 402462 856
rect 402630 2 403290 856
rect 403458 2 404210 856
rect 404378 2 405038 856
rect 405206 2 405958 856
rect 406126 2 406786 856
rect 406954 2 407614 856
rect 407782 2 408534 856
rect 408702 2 409362 856
rect 409530 2 410190 856
rect 410358 2 411110 856
rect 411278 2 411938 856
rect 412106 2 412766 856
rect 412934 2 413686 856
rect 413854 2 414514 856
rect 414682 2 415434 856
rect 415602 2 416262 856
rect 416430 2 417090 856
rect 417258 2 418010 856
rect 418178 2 418838 856
rect 419006 2 419666 856
rect 419834 2 420586 856
rect 420754 2 421414 856
rect 421582 2 422242 856
rect 422410 2 423162 856
rect 423330 2 423990 856
rect 424158 2 424378 856
<< obsm3 >>
rect 2681 171 424383 424353
<< metal4 >>
rect 4208 2128 4528 424368
rect 19568 2128 19888 424368
rect 34928 2128 35248 424368
rect 50288 2128 50608 424368
rect 65648 2128 65968 424368
rect 81008 2128 81328 424368
rect 96368 2128 96688 424368
rect 111728 2128 112048 424368
rect 127088 2128 127408 424368
rect 142448 2128 142768 424368
rect 157808 2128 158128 424368
rect 173168 2128 173488 424368
rect 188528 2128 188848 424368
rect 203888 2128 204208 424368
rect 219248 2128 219568 424368
rect 234608 2128 234928 424368
rect 249968 2128 250288 424368
rect 265328 2128 265648 424368
rect 280688 2128 281008 424368
rect 296048 2128 296368 424368
rect 311408 2128 311728 424368
rect 326768 2128 327088 424368
rect 342128 2128 342448 424368
rect 357488 2128 357808 424368
rect 372848 2128 373168 424368
rect 388208 2128 388528 424368
rect 403568 2128 403888 424368
rect 418928 2128 419248 424368
<< obsm4 >>
rect 19011 2048 19488 424149
rect 19968 2048 34848 424149
rect 35328 2048 50208 424149
rect 50688 2048 65568 424149
rect 66048 2048 80928 424149
rect 81408 2048 96288 424149
rect 96768 2048 111648 424149
rect 112128 2048 127008 424149
rect 127488 2048 142368 424149
rect 142848 2048 157728 424149
rect 158208 2048 173088 424149
rect 173568 2048 188448 424149
rect 188928 2048 203808 424149
rect 204288 2048 219168 424149
rect 219648 2048 234528 424149
rect 235008 2048 249888 424149
rect 250368 2048 265248 424149
rect 265728 2048 280608 424149
rect 281088 2048 295968 424149
rect 296448 2048 311328 424149
rect 311808 2048 326688 424149
rect 327168 2048 342048 424149
rect 342528 2048 357408 424149
rect 357888 2048 372768 424149
rect 373248 2048 388128 424149
rect 388608 2048 403488 424149
rect 403968 2048 418848 424149
rect 419328 2048 422773 424149
rect 19011 1531 422773 2048
<< labels >>
rlabel metal2 s 1858 425904 1914 426704 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 113546 425904 113602 426704 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 124678 425904 124734 426704 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 135902 425904 135958 426704 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 147034 425904 147090 426704 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 158258 425904 158314 426704 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 169390 425904 169446 426704 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 180614 425904 180670 426704 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 191746 425904 191802 426704 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 202970 425904 203026 426704 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 214102 425904 214158 426704 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 12990 425904 13046 426704 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 225234 425904 225290 426704 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 236458 425904 236514 426704 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 247590 425904 247646 426704 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 258814 425904 258870 426704 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 269946 425904 270002 426704 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 281170 425904 281226 426704 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 292302 425904 292358 426704 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 303526 425904 303582 426704 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 314658 425904 314714 426704 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 325790 425904 325846 426704 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 24122 425904 24178 426704 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 337014 425904 337070 426704 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 348146 425904 348202 426704 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 359370 425904 359426 426704 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 370502 425904 370558 426704 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 381726 425904 381782 426704 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 392858 425904 392914 426704 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 404082 425904 404138 426704 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 415214 425904 415270 426704 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 35346 425904 35402 426704 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 46478 425904 46534 426704 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 57702 425904 57758 426704 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 68834 425904 68890 426704 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 80058 425904 80114 426704 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 91190 425904 91246 426704 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 102414 425904 102470 426704 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5538 425904 5594 426704 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 117226 425904 117282 426704 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 128450 425904 128506 426704 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 139582 425904 139638 426704 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 150806 425904 150862 426704 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 161938 425904 161994 426704 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 173162 425904 173218 426704 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 184294 425904 184350 426704 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 195518 425904 195574 426704 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 206650 425904 206706 426704 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 217782 425904 217838 426704 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 16670 425904 16726 426704 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 229006 425904 229062 426704 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 240138 425904 240194 426704 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 251362 425904 251418 426704 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 262494 425904 262550 426704 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 273718 425904 273774 426704 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 284850 425904 284906 426704 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 296074 425904 296130 426704 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 307206 425904 307262 426704 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 318430 425904 318486 426704 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 329562 425904 329618 426704 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 27894 425904 27950 426704 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 340694 425904 340750 426704 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 351918 425904 351974 426704 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 363050 425904 363106 426704 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 374274 425904 374330 426704 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 385406 425904 385462 426704 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 396630 425904 396686 426704 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 407762 425904 407818 426704 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 418986 425904 419042 426704 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 39026 425904 39082 426704 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 50250 425904 50306 426704 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 61382 425904 61438 426704 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 72606 425904 72662 426704 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 83738 425904 83794 426704 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 94962 425904 95018 426704 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 106094 425904 106150 426704 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9218 425904 9274 426704 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 120998 425904 121054 426704 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 132130 425904 132186 426704 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 143354 425904 143410 426704 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 154486 425904 154542 426704 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 165710 425904 165766 426704 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 176842 425904 176898 426704 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 188066 425904 188122 426704 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 199198 425904 199254 426704 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 210422 425904 210478 426704 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 221554 425904 221610 426704 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 20442 425904 20498 426704 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 232686 425904 232742 426704 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 243910 425904 243966 426704 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 255042 425904 255098 426704 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 266266 425904 266322 426704 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 277398 425904 277454 426704 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 288622 425904 288678 426704 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 299754 425904 299810 426704 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 310978 425904 311034 426704 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 322110 425904 322166 426704 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 333242 425904 333298 426704 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 31574 425904 31630 426704 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 344466 425904 344522 426704 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 355598 425904 355654 426704 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 366822 425904 366878 426704 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 377954 425904 378010 426704 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 389178 425904 389234 426704 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 400310 425904 400366 426704 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 411534 425904 411590 426704 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 422666 425904 422722 426704 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 42798 425904 42854 426704 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 53930 425904 53986 426704 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 65154 425904 65210 426704 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 76286 425904 76342 426704 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 87510 425904 87566 426704 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 98642 425904 98698 426704 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 109774 425904 109830 426704 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 422298 0 422354 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 423218 0 423274 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 424046 0 424102 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 349986 0 350042 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 352562 0 352618 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 355138 0 355194 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 357714 0 357770 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 360290 0 360346 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 362958 0 363014 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 365534 0 365590 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 368110 0 368166 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 370686 0 370742 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 373262 0 373318 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 375838 0 375894 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 378414 0 378470 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 380990 0 381046 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 383566 0 383622 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 386142 0 386198 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 388718 0 388774 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 391294 0 391350 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 393962 0 394018 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 396538 0 396594 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 399114 0 399170 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 401690 0 401746 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 404266 0 404322 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 406842 0 406898 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 409418 0 409474 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 411994 0 412050 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 414570 0 414626 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 417146 0 417202 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 419722 0 419778 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 179510 0 179566 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 184662 0 184718 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 192390 0 192446 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 200118 0 200174 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 202694 0 202750 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 207938 0 207994 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 213090 0 213146 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 220818 0 220874 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 223394 0 223450 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 228546 0 228602 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 233698 0 233754 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 236274 0 236330 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 238942 0 238998 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 241518 0 241574 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 249246 0 249302 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 251822 0 251878 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 256974 0 257030 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 264702 0 264758 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 267278 0 267334 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 269946 0 270002 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 272522 0 272578 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 275098 0 275154 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 277674 0 277730 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 285402 0 285458 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 287978 0 288034 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 290554 0 290610 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 293130 0 293186 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 295706 0 295762 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 298282 0 298338 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 300950 0 301006 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 303526 0 303582 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 306102 0 306158 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 308678 0 308734 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 311254 0 311310 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 313830 0 313886 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 316406 0 316462 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 318982 0 319038 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 321558 0 321614 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 324134 0 324190 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 326710 0 326766 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 329286 0 329342 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 331954 0 332010 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 334530 0 334586 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 337106 0 337162 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 339682 0 339738 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 342258 0 342314 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 344834 0 344890 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 347410 0 347466 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 350814 0 350870 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 353482 0 353538 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 356058 0 356114 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 358634 0 358690 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 361210 0 361266 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 363786 0 363842 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 366362 0 366418 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 368938 0 368994 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 371514 0 371570 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 374090 0 374146 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 376666 0 376722 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 379242 0 379298 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 381818 0 381874 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 384486 0 384542 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 387062 0 387118 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 389638 0 389694 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 392214 0 392270 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 394790 0 394846 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 397366 0 397422 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 399942 0 399998 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 402518 0 402574 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 405094 0 405150 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 407670 0 407726 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 410246 0 410302 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 412822 0 412878 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 415490 0 415546 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 418066 0 418122 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 420642 0 420698 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 133786 0 133842 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 136454 0 136510 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 139030 0 139086 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 144182 0 144238 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 162214 0 162270 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 170034 0 170090 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 177762 0 177818 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 180338 0 180394 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 182914 0 182970 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 188066 0 188122 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 190642 0 190698 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 198462 0 198518 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 203614 0 203670 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 206190 0 206246 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 208766 0 208822 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 211342 0 211398 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 213918 0 213974 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 216494 0 216550 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 219070 0 219126 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 221646 0 221702 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 224222 0 224278 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 226798 0 226854 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 229466 0 229522 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 232042 0 232098 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 234618 0 234674 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 237194 0 237250 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 239770 0 239826 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 242346 0 242402 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 244922 0 244978 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 247498 0 247554 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 250074 0 250130 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 252650 0 252706 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 255226 0 255282 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 257802 0 257858 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 263046 0 263102 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 265622 0 265678 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 268198 0 268254 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 270774 0 270830 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 273350 0 273406 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 275926 0 275982 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 278502 0 278558 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 281078 0 281134 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 283654 0 283710 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 286230 0 286286 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 288806 0 288862 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 291474 0 291530 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 294050 0 294106 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 296626 0 296682 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 299202 0 299258 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 301778 0 301834 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 304354 0 304410 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 306930 0 306986 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 309506 0 309562 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 312082 0 312138 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 314658 0 314714 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 317234 0 317290 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 319810 0 319866 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 322478 0 322534 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 113178 0 113234 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 325054 0 325110 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 327630 0 327686 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 330206 0 330262 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 332782 0 332838 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 335358 0 335414 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 337934 0 337990 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 340510 0 340566 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 343086 0 343142 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 345662 0 345718 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 348238 0 348294 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 115754 0 115810 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 351734 0 351790 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 354310 0 354366 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 356886 0 356942 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 359462 0 359518 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 362038 0 362094 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 364614 0 364670 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 367190 0 367246 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 369766 0 369822 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 372342 0 372398 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 375010 0 375066 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 377586 0 377642 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 380162 0 380218 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 382738 0 382794 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 385314 0 385370 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 387890 0 387946 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 390466 0 390522 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 393042 0 393098 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 395618 0 395674 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 398194 0 398250 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 400770 0 400826 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 403346 0 403402 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 406014 0 406070 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 408590 0 408646 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 411166 0 411222 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 413742 0 413798 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 416318 0 416374 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 418894 0 418950 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 421470 0 421526 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 170862 0 170918 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 176014 0 176070 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 181166 0 181222 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 188986 0 189042 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 196714 0 196770 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 201866 0 201922 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 204442 0 204498 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 212170 0 212226 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 214746 0 214802 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 217322 0 217378 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 219990 0 220046 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 222566 0 222622 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 227718 0 227774 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 230294 0 230350 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 232870 0 232926 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 240598 0 240654 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 243174 0 243230 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 245750 0 245806 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 248326 0 248382 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 250994 0 251050 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 253570 0 253626 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 256146 0 256202 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 258722 0 258778 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 261298 0 261354 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 263874 0 263930 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 266450 0 266506 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 269026 0 269082 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 271602 0 271658 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 274178 0 274234 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 276754 0 276810 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 279330 0 279386 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 281998 0 282054 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 287150 0 287206 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 289726 0 289782 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 292302 0 292358 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 294878 0 294934 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 297454 0 297510 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 300030 0 300086 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 302606 0 302662 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 305182 0 305238 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 307758 0 307814 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 310334 0 310390 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 313002 0 313058 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 315578 0 315634 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 318154 0 318210 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 320730 0 320786 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 323306 0 323362 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 325882 0 325938 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 328458 0 328514 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 331034 0 331090 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 333610 0 333666 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 336186 0 336242 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 338762 0 338818 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 341338 0 341394 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 344006 0 344062 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 346582 0 346638 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 349158 0 349214 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 424368 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 424368 6 vssd1
port 503 nsew ground input
rlabel metal4 s 418928 2128 419248 424368 6 vssd1
port 503 nsew ground input
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 424560 426704
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 467978368
string GDS_START 1813940
<< end >>

