magic
tech sky130A
magscale 1 2
timestamp 1635447575
<< locali >>
rect 289955 578085 290105 578119
rect 109877 574311 109911 574889
rect 117697 574107 117731 574889
rect 145021 574583 145055 574889
rect 164801 574379 164835 574889
rect 176577 574515 176611 574889
rect 180441 574651 180475 574889
rect 391857 574855 391891 575025
rect 403449 574719 403483 575025
rect 415409 574447 415443 575025
rect 438869 574243 438903 575025
rect 450553 574787 450587 575025
rect 462329 574175 462363 575025
rect 175933 126803 175967 126905
rect 176025 126055 176059 126769
rect 484777 126599 484811 126701
rect 493057 126463 493091 126701
rect 214573 125851 214607 126361
rect 465733 126123 465767 126429
rect 496001 126259 496035 126429
rect 512745 125851 512779 126225
rect 514033 125919 514067 126837
rect 53297 4743 53331 4981
rect 485053 4607 485087 5253
rect 88993 3927 89027 4097
rect 88901 3655 88935 3893
rect 35265 3315 35299 3621
rect 74825 3621 75135 3655
rect 83047 3621 83197 3655
rect 74825 3587 74859 3621
rect 75101 3587 75135 3621
rect 75101 3553 76205 3587
rect 74917 3451 74951 3553
rect 89085 3451 89119 4097
rect 91661 3723 91695 4097
rect 91569 3451 91603 3689
rect 52469 3043 52503 3349
rect 95433 3247 95467 4097
rect 432923 4029 433073 4063
rect 437305 3995 437339 4097
rect 95525 3179 95559 3893
rect 102149 3315 102183 3621
rect 123401 3451 123435 3689
rect 132877 3519 132911 3689
rect 142353 3315 142387 3689
rect 149069 3315 149103 3485
rect 125977 2975 126011 3077
rect 172989 2975 173023 3757
rect 173081 3519 173115 3757
rect 173725 3519 173759 3553
rect 187065 3519 187099 3621
rect 173725 3485 173909 3519
rect 200129 3383 200163 3553
rect 407313 3247 407347 3689
rect 412097 3247 412131 3689
rect 417157 3689 417651 3723
rect 417157 3587 417191 3689
rect 417617 3655 417651 3689
rect 417249 3451 417283 3553
rect 125977 2941 126161 2975
rect 412005 2839 412039 3213
rect 417341 3179 417375 3417
rect 417433 3043 417467 3145
rect 417525 3043 417559 3621
rect 417985 3519 418019 3689
rect 419089 2907 419123 3621
rect 421665 3519 421699 3689
rect 424793 3417 425069 3451
rect 424793 3179 424827 3417
rect 426265 2975 426299 3417
rect 427093 2975 427127 3145
rect 427185 3043 427219 3553
rect 436937 3383 436971 3961
rect 428565 3179 428599 3349
rect 428657 3043 428691 3145
rect 436753 3111 436787 3281
rect 436695 3077 436787 3111
rect 436845 3043 436879 3349
rect 427277 2975 427311 3009
rect 427093 2941 427311 2975
<< viali >>
rect 289921 578085 289955 578119
rect 290105 578085 290139 578119
rect 391857 575025 391891 575059
rect 109877 574889 109911 574923
rect 109877 574277 109911 574311
rect 117697 574889 117731 574923
rect 145021 574889 145055 574923
rect 145021 574549 145055 574583
rect 164801 574889 164835 574923
rect 176577 574889 176611 574923
rect 180441 574889 180475 574923
rect 391857 574821 391891 574855
rect 403449 575025 403483 575059
rect 403449 574685 403483 574719
rect 415409 575025 415443 575059
rect 180441 574617 180475 574651
rect 176577 574481 176611 574515
rect 415409 574413 415443 574447
rect 438869 575025 438903 575059
rect 164801 574345 164835 574379
rect 450553 575025 450587 575059
rect 450553 574753 450587 574787
rect 462329 575025 462363 575059
rect 438869 574209 438903 574243
rect 462329 574141 462363 574175
rect 117697 574073 117731 574107
rect 175933 126905 175967 126939
rect 514033 126837 514067 126871
rect 175933 126769 175967 126803
rect 176025 126769 176059 126803
rect 484777 126701 484811 126735
rect 484777 126565 484811 126599
rect 493057 126701 493091 126735
rect 465733 126429 465767 126463
rect 493057 126429 493091 126463
rect 496001 126429 496035 126463
rect 176025 126021 176059 126055
rect 214573 126361 214607 126395
rect 496001 126225 496035 126259
rect 512745 126225 512779 126259
rect 465733 126089 465767 126123
rect 214573 125817 214607 125851
rect 514033 125885 514067 125919
rect 512745 125817 512779 125851
rect 485053 5253 485087 5287
rect 53297 4981 53331 5015
rect 53297 4709 53331 4743
rect 485053 4573 485087 4607
rect 88993 4097 89027 4131
rect 88901 3893 88935 3927
rect 88993 3893 89027 3927
rect 89085 4097 89119 4131
rect 35265 3621 35299 3655
rect 83013 3621 83047 3655
rect 83197 3621 83231 3655
rect 88901 3621 88935 3655
rect 74825 3553 74859 3587
rect 74917 3553 74951 3587
rect 76205 3553 76239 3587
rect 74917 3417 74951 3451
rect 91661 4097 91695 4131
rect 89085 3417 89119 3451
rect 91569 3689 91603 3723
rect 91661 3689 91695 3723
rect 95433 4097 95467 4131
rect 91569 3417 91603 3451
rect 35265 3281 35299 3315
rect 52469 3349 52503 3383
rect 437305 4097 437339 4131
rect 432889 4029 432923 4063
rect 433073 4029 433107 4063
rect 436937 3961 436971 3995
rect 437305 3961 437339 3995
rect 95433 3213 95467 3247
rect 95525 3893 95559 3927
rect 172989 3757 173023 3791
rect 123401 3689 123435 3723
rect 102149 3621 102183 3655
rect 132877 3689 132911 3723
rect 132877 3485 132911 3519
rect 142353 3689 142387 3723
rect 123401 3417 123435 3451
rect 102149 3281 102183 3315
rect 142353 3281 142387 3315
rect 149069 3485 149103 3519
rect 149069 3281 149103 3315
rect 95525 3145 95559 3179
rect 52469 3009 52503 3043
rect 125977 3077 126011 3111
rect 173081 3757 173115 3791
rect 407313 3689 407347 3723
rect 187065 3621 187099 3655
rect 173081 3485 173115 3519
rect 173725 3553 173759 3587
rect 173909 3485 173943 3519
rect 187065 3485 187099 3519
rect 200129 3553 200163 3587
rect 200129 3349 200163 3383
rect 412097 3689 412131 3723
rect 417525 3621 417559 3655
rect 417617 3621 417651 3655
rect 417985 3689 418019 3723
rect 417157 3553 417191 3587
rect 417249 3553 417283 3587
rect 417249 3417 417283 3451
rect 417341 3417 417375 3451
rect 407313 3213 407347 3247
rect 412005 3213 412039 3247
rect 412097 3213 412131 3247
rect 126161 2941 126195 2975
rect 172989 2941 173023 2975
rect 417341 3145 417375 3179
rect 417433 3145 417467 3179
rect 417433 3009 417467 3043
rect 421665 3689 421699 3723
rect 417985 3485 418019 3519
rect 419089 3621 419123 3655
rect 417525 3009 417559 3043
rect 421665 3485 421699 3519
rect 427185 3553 427219 3587
rect 425069 3417 425103 3451
rect 426265 3417 426299 3451
rect 424793 3145 424827 3179
rect 426265 2941 426299 2975
rect 427093 3145 427127 3179
rect 428565 3349 428599 3383
rect 436845 3349 436879 3383
rect 436937 3349 436971 3383
rect 436753 3281 436787 3315
rect 428565 3145 428599 3179
rect 428657 3145 428691 3179
rect 436661 3077 436695 3111
rect 427185 3009 427219 3043
rect 427277 3009 427311 3043
rect 428657 3009 428691 3043
rect 436845 3009 436879 3043
rect 419089 2873 419123 2907
rect 412005 2805 412039 2839
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 324314 700992 324320 701004
rect 154172 700964 324320 700992
rect 154172 700952 154178 700964
rect 324314 700952 324320 700964
rect 324372 700952 324378 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 320174 700924 320180 700936
rect 137888 700896 320180 700924
rect 137888 700884 137894 700896
rect 320174 700884 320180 700896
rect 320232 700884 320238 700936
rect 263502 700816 263508 700868
rect 263560 700856 263566 700868
rect 462314 700856 462320 700868
rect 263560 700828 462320 700856
rect 263560 700816 263566 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 267642 700748 267648 700800
rect 267700 700788 267706 700800
rect 478506 700788 478512 700800
rect 267700 700760 478512 700788
rect 267700 700748 267706 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 336734 700720 336740 700732
rect 89220 700692 336740 700720
rect 89220 700680 89226 700692
rect 336734 700680 336740 700692
rect 336792 700680 336798 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 332594 700652 332600 700664
rect 73028 700624 332600 700652
rect 73028 700612 73034 700624
rect 332594 700612 332600 700624
rect 332652 700612 332658 700664
rect 251082 700544 251088 700596
rect 251140 700584 251146 700596
rect 527174 700584 527180 700596
rect 251140 700556 527180 700584
rect 251140 700544 251146 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 255222 700476 255228 700528
rect 255280 700516 255286 700528
rect 543458 700516 543464 700528
rect 255280 700488 543464 700516
rect 255280 700476 255286 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 340874 700448 340880 700460
rect 40552 700420 340880 700448
rect 40552 700408 40558 700420
rect 340874 700408 340880 700420
rect 340932 700408 340938 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 347774 700380 347780 700392
rect 24360 700352 347780 700380
rect 24360 700340 24366 700352
rect 347774 700340 347780 700352
rect 347832 700340 347838 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 343634 700312 343640 700324
rect 8168 700284 343640 700312
rect 8168 700272 8174 700284
rect 343634 700272 343640 700284
rect 343692 700272 343698 700324
rect 278682 700204 278688 700256
rect 278740 700244 278746 700256
rect 413646 700244 413652 700256
rect 278740 700216 413652 700244
rect 278740 700204 278746 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 274542 700136 274548 700188
rect 274600 700176 274606 700188
rect 397454 700176 397460 700188
rect 274600 700148 397460 700176
rect 274600 700136 274606 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 309134 700108 309140 700120
rect 202840 700080 309140 700108
rect 202840 700068 202846 700080
rect 309134 700068 309140 700080
rect 309192 700068 309198 700120
rect 218974 700000 218980 700052
rect 219032 700040 219038 700052
rect 313274 700040 313280 700052
rect 219032 700012 313280 700040
rect 219032 700000 219038 700012
rect 313274 700000 313280 700012
rect 313332 700000 313338 700052
rect 291102 699932 291108 699984
rect 291160 699972 291166 699984
rect 348786 699972 348792 699984
rect 291160 699944 348792 699972
rect 291160 699932 291166 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 286962 699864 286968 699916
rect 287020 699904 287026 699916
rect 332502 699904 332508 699916
rect 287020 699876 332508 699904
rect 287020 699864 287026 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 267550 699796 267556 699848
rect 267608 699836 267614 699848
rect 296714 699836 296720 699848
rect 267608 699808 296720 699836
rect 267608 699796 267614 699808
rect 296714 699796 296720 699808
rect 296772 699796 296778 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 300854 699768 300860 699780
rect 283892 699740 300860 699768
rect 283892 699728 283898 699740
rect 300854 699728 300860 699740
rect 300912 699728 300918 699780
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 240042 696940 240048 696992
rect 240100 696980 240106 696992
rect 580166 696980 580172 696992
rect 240100 696952 580172 696980
rect 240100 696940 240106 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 244182 683204 244188 683256
rect 244240 683244 244246 683256
rect 580166 683244 580172 683256
rect 244240 683216 580172 683244
rect 244240 683204 244246 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 351914 683176 351920 683188
rect 3476 683148 351920 683176
rect 3476 683136 3482 683148
rect 351914 683136 351920 683148
rect 351972 683136 351978 683188
rect 235810 670760 235816 670812
rect 235868 670800 235874 670812
rect 580166 670800 580172 670812
rect 235868 670772 580172 670800
rect 235868 670760 235874 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 360194 670732 360200 670744
rect 3568 670704 360200 670732
rect 3568 670692 3574 670704
rect 360194 670692 360200 670704
rect 360252 670692 360258 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 356054 656928 356060 656940
rect 3476 656900 356060 656928
rect 3476 656888 3482 656900
rect 356054 656888 356060 656900
rect 356112 656888 356118 656940
rect 227622 643084 227628 643136
rect 227680 643124 227686 643136
rect 580166 643124 580172 643136
rect 227680 643096 580172 643124
rect 227680 643084 227686 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 364426 632108 364432 632120
rect 3476 632080 364432 632108
rect 3476 632068 3482 632080
rect 364426 632068 364432 632080
rect 364484 632068 364490 632120
rect 231762 630640 231768 630692
rect 231820 630680 231826 630692
rect 580166 630680 580172 630692
rect 231820 630652 580172 630680
rect 231820 630640 231826 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 371234 618304 371240 618316
rect 3200 618276 371240 618304
rect 3200 618264 3206 618276
rect 371234 618264 371240 618276
rect 371292 618264 371298 618316
rect 223482 616836 223488 616888
rect 223540 616876 223546 616888
rect 580166 616876 580172 616888
rect 223540 616848 580172 616876
rect 223540 616836 223546 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 367094 605860 367100 605872
rect 3292 605832 367100 605860
rect 3292 605820 3298 605832
rect 367094 605820 367100 605832
rect 367152 605820 367158 605872
rect 216582 590656 216588 590708
rect 216640 590696 216646 590708
rect 579798 590696 579804 590708
rect 216640 590668 579804 590696
rect 216640 590656 216646 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 375834 579680 375840 579692
rect 3384 579652 375840 579680
rect 3384 579640 3390 579652
rect 375834 579640 375840 579652
rect 375892 579640 375898 579692
rect 4798 578280 4804 578332
rect 4856 578320 4862 578332
rect 430850 578320 430856 578332
rect 4856 578292 430856 578320
rect 4856 578280 4862 578292
rect 430850 578280 430856 578292
rect 430908 578280 430914 578332
rect 14458 578212 14464 578264
rect 14516 578252 14522 578264
rect 442626 578252 442632 578264
rect 14516 578224 442632 578252
rect 14516 578212 14522 578224
rect 442626 578212 442632 578224
rect 442684 578212 442690 578264
rect 215754 578144 215760 578196
rect 215812 578184 215818 578196
rect 216582 578184 216588 578196
rect 215812 578156 216588 578184
rect 215812 578144 215818 578156
rect 216582 578144 216588 578156
rect 216640 578144 216646 578196
rect 235350 578144 235356 578196
rect 235408 578184 235414 578196
rect 235810 578184 235816 578196
rect 235408 578156 235816 578184
rect 235408 578144 235414 578156
rect 235810 578144 235816 578156
rect 235868 578144 235874 578196
rect 239306 578144 239312 578196
rect 239364 578184 239370 578196
rect 240042 578184 240048 578196
rect 239364 578156 240048 578184
rect 239364 578144 239370 578156
rect 240042 578144 240048 578156
rect 240100 578144 240106 578196
rect 243262 578144 243268 578196
rect 243320 578184 243326 578196
rect 244182 578184 244188 578196
rect 243320 578156 244188 578184
rect 243320 578144 243326 578156
rect 244182 578144 244188 578156
rect 244240 578144 244246 578196
rect 262858 578144 262864 578196
rect 262916 578184 262922 578196
rect 263502 578184 263508 578196
rect 262916 578156 263508 578184
rect 262916 578144 262922 578156
rect 263502 578144 263508 578156
rect 263560 578144 263566 578196
rect 266814 578144 266820 578196
rect 266872 578184 266878 578196
rect 267642 578184 267648 578196
rect 266872 578156 267648 578184
rect 266872 578144 266878 578156
rect 267642 578144 267648 578156
rect 267700 578144 267706 578196
rect 282454 578144 282460 578196
rect 282512 578184 282518 578196
rect 282512 578156 290044 578184
rect 282512 578144 282518 578156
rect 235902 578076 235908 578128
rect 235960 578116 235966 578128
rect 289909 578119 289967 578125
rect 289909 578116 289921 578119
rect 235960 578088 289921 578116
rect 235960 578076 235966 578088
rect 289909 578085 289921 578088
rect 289955 578085 289967 578119
rect 289909 578079 289967 578085
rect 286410 578008 286416 578060
rect 286468 578048 286474 578060
rect 286962 578048 286968 578060
rect 286468 578020 286968 578048
rect 286468 578008 286474 578020
rect 286962 578008 286968 578020
rect 287020 578008 287026 578060
rect 290016 578048 290044 578156
rect 290274 578144 290280 578196
rect 290332 578184 290338 578196
rect 291102 578184 291108 578196
rect 290332 578156 291108 578184
rect 290332 578144 290338 578156
rect 291102 578144 291108 578156
rect 291160 578144 291166 578196
rect 293862 578144 293868 578196
rect 293920 578184 293926 578196
rect 299474 578184 299480 578196
rect 293920 578156 299480 578184
rect 293920 578144 293926 578156
rect 299474 578144 299480 578156
rect 299532 578144 299538 578196
rect 290093 578119 290151 578125
rect 290093 578085 290105 578119
rect 290139 578116 290151 578119
rect 305362 578116 305368 578128
rect 290139 578088 305368 578116
rect 290139 578085 290151 578088
rect 290093 578079 290151 578085
rect 305362 578076 305368 578088
rect 305420 578076 305426 578128
rect 364334 578048 364340 578060
rect 290016 578020 364340 578048
rect 364334 578008 364340 578020
rect 364392 578008 364398 578060
rect 171042 577940 171048 577992
rect 171100 577980 171106 577992
rect 317414 577980 317420 577992
rect 171100 577952 317420 577980
rect 171100 577940 171106 577952
rect 317414 577940 317420 577952
rect 317472 577940 317478 577992
rect 270402 577872 270408 577924
rect 270460 577912 270466 577924
rect 429194 577912 429200 577924
rect 270460 577884 429200 577912
rect 270460 577872 270466 577884
rect 429194 577872 429200 577884
rect 429252 577872 429258 577924
rect 106182 577804 106188 577856
rect 106240 577844 106246 577856
rect 328914 577844 328920 577856
rect 106240 577816 328920 577844
rect 106240 577804 106246 577816
rect 328914 577804 328920 577816
rect 328972 577804 328978 577856
rect 258902 577736 258908 577788
rect 258960 577776 258966 577788
rect 494054 577776 494060 577788
rect 258960 577748 494060 577776
rect 258960 577736 258966 577748
rect 494054 577736 494060 577748
rect 494112 577736 494118 577788
rect 246942 577668 246948 577720
rect 247000 577708 247006 577720
rect 558914 577708 558920 577720
rect 247000 577680 558920 577708
rect 247000 577668 247006 577680
rect 558914 577668 558920 577680
rect 558972 577668 558978 577720
rect 53098 577600 53104 577652
rect 53156 577640 53162 577652
rect 407390 577640 407396 577652
rect 53156 577612 407396 577640
rect 53156 577600 53162 577612
rect 407390 577600 407396 577612
rect 407448 577600 407454 577652
rect 184382 577532 184388 577584
rect 184440 577572 184446 577584
rect 538858 577572 538864 577584
rect 184440 577544 538864 577572
rect 184440 577532 184446 577544
rect 538858 577532 538864 577544
rect 538916 577532 538922 577584
rect 219342 577464 219348 577516
rect 219400 577504 219406 577516
rect 580166 577504 580172 577516
rect 219400 577476 580172 577504
rect 219400 577464 219406 577476
rect 580166 577464 580172 577476
rect 580224 577464 580230 577516
rect 172422 577396 172428 577448
rect 172480 577436 172486 577448
rect 537478 577436 537484 577448
rect 172480 577408 537484 577436
rect 172480 577396 172486 577408
rect 537478 577396 537484 577408
rect 537536 577396 537542 577448
rect 160830 577328 160836 577380
rect 160888 577368 160894 577380
rect 536098 577368 536104 577380
rect 160888 577340 536104 577368
rect 160888 577328 160894 577340
rect 536098 577328 536104 577340
rect 536156 577328 536162 577380
rect 168742 577260 168748 577312
rect 168800 577300 168806 577312
rect 551278 577300 551284 577312
rect 168800 577272 551284 577300
rect 168800 577260 168806 577272
rect 551278 577260 551284 577272
rect 551336 577260 551342 577312
rect 148962 577192 148968 577244
rect 149020 577232 149026 577244
rect 533338 577232 533344 577244
rect 149020 577204 533344 577232
rect 149020 577192 149026 577204
rect 533338 577192 533344 577204
rect 533396 577192 533402 577244
rect 137278 577124 137284 577176
rect 137336 577164 137342 577176
rect 530578 577164 530584 577176
rect 137336 577136 530584 577164
rect 137336 577124 137342 577136
rect 530578 577124 530584 577136
rect 530636 577124 530642 577176
rect 125318 577056 125324 577108
rect 125376 577096 125382 577108
rect 529198 577096 529204 577108
rect 125376 577068 529204 577096
rect 125376 577056 125382 577068
rect 529198 577056 529204 577068
rect 529256 577056 529262 577108
rect 121362 576988 121368 577040
rect 121420 577028 121426 577040
rect 542998 577028 543004 577040
rect 121420 577000 543004 577028
rect 121420 576988 121426 577000
rect 542998 576988 543004 577000
rect 543056 576988 543062 577040
rect 17218 576920 17224 576972
rect 17276 576960 17282 576972
rect 454402 576960 454408 576972
rect 17276 576932 454408 576960
rect 17276 576920 17282 576932
rect 454402 576920 454408 576932
rect 454460 576920 454466 576972
rect 18598 576852 18604 576904
rect 18656 576892 18662 576904
rect 466454 576892 466460 576904
rect 18656 576864 466460 576892
rect 18656 576852 18662 576864
rect 466454 576852 466460 576864
rect 466512 576852 466518 576904
rect 211890 576716 211896 576768
rect 211948 576756 211954 576768
rect 519538 576756 519544 576768
rect 211948 576728 519544 576756
rect 211948 576716 211954 576728
rect 519538 576716 519544 576728
rect 519596 576716 519602 576768
rect 199930 576648 199936 576700
rect 199988 576688 199994 576700
rect 518158 576688 518164 576700
rect 199988 576660 518164 576688
rect 199988 576648 199994 576660
rect 518158 576648 518164 576660
rect 518216 576648 518222 576700
rect 188338 576580 188344 576632
rect 188396 576620 188402 576632
rect 516778 576620 516784 576632
rect 188396 576592 516784 576620
rect 188396 576580 188402 576592
rect 516778 576580 516784 576592
rect 516836 576580 516842 576632
rect 66898 576512 66904 576564
rect 66956 576552 66962 576564
rect 423030 576552 423036 576564
rect 66956 576524 423036 576552
rect 66956 576512 66962 576524
rect 423030 576512 423036 576524
rect 423088 576512 423094 576564
rect 36538 576444 36544 576496
rect 36596 576484 36602 576496
rect 399478 576484 399484 576496
rect 36596 576456 399484 576484
rect 36596 576444 36602 576456
rect 399478 576444 399484 576456
rect 399536 576444 399542 576496
rect 57238 576376 57244 576428
rect 57296 576416 57302 576428
rect 426986 576416 426992 576428
rect 57296 576388 426992 576416
rect 57296 576376 57302 576388
rect 426986 576376 426992 576388
rect 427044 576376 427050 576428
rect 153010 576308 153016 576360
rect 153068 576348 153074 576360
rect 525058 576348 525064 576360
rect 153068 576320 525064 576348
rect 153068 576308 153074 576320
rect 525058 576308 525064 576320
rect 525116 576308 525122 576360
rect 61378 576240 61384 576292
rect 61436 576280 61442 576292
rect 434806 576280 434812 576292
rect 61436 576252 434812 576280
rect 61436 576240 61442 576252
rect 434806 576240 434812 576252
rect 434864 576240 434870 576292
rect 11698 576172 11704 576224
rect 11756 576212 11762 576224
rect 387794 576212 387800 576224
rect 11756 576184 387800 576212
rect 11756 576172 11762 576184
rect 387794 576172 387800 576184
rect 387852 576172 387858 576224
rect 39298 576104 39304 576156
rect 39356 576144 39362 576156
rect 419074 576144 419080 576156
rect 39356 576116 419080 576144
rect 39356 576104 39362 576116
rect 419074 576104 419080 576116
rect 419132 576104 419138 576156
rect 65518 576036 65524 576088
rect 65576 576076 65582 576088
rect 446582 576076 446588 576088
rect 65576 576048 446588 576076
rect 65576 576036 65582 576048
rect 446582 576036 446588 576048
rect 446640 576036 446646 576088
rect 141234 575968 141240 576020
rect 141292 576008 141298 576020
rect 522298 576008 522304 576020
rect 141292 575980 522304 576008
rect 141292 575968 141298 575980
rect 522298 575968 522304 575980
rect 522356 575968 522362 576020
rect 25498 575900 25504 575952
rect 25556 575940 25562 575952
rect 411254 575940 411260 575952
rect 25556 575912 411260 575940
rect 25556 575900 25562 575912
rect 411254 575900 411260 575912
rect 411312 575900 411318 575952
rect 156966 575832 156972 575884
rect 157024 575872 157030 575884
rect 548518 575872 548524 575884
rect 157024 575844 548524 575872
rect 157024 575832 157030 575844
rect 548518 575832 548524 575844
rect 548576 575832 548582 575884
rect 129458 575764 129464 575816
rect 129516 575804 129522 575816
rect 520918 575804 520924 575816
rect 129516 575776 520924 575804
rect 129516 575764 129522 575776
rect 520918 575764 520924 575776
rect 520976 575764 520982 575816
rect 47578 575696 47584 575748
rect 47636 575736 47642 575748
rect 458680 575736 458686 575748
rect 47636 575708 458686 575736
rect 47636 575696 47642 575708
rect 458680 575696 458686 575708
rect 458738 575696 458744 575748
rect 133414 575628 133420 575680
rect 133472 575668 133478 575680
rect 544378 575668 544384 575680
rect 133472 575640 544384 575668
rect 133472 575628 133478 575640
rect 544378 575628 544384 575640
rect 544436 575628 544442 575680
rect 51718 575560 51724 575612
rect 51776 575600 51782 575612
rect 470134 575600 470140 575612
rect 51776 575572 470140 575600
rect 51776 575560 51782 575572
rect 470134 575560 470140 575572
rect 470192 575560 470198 575612
rect 50338 575492 50344 575544
rect 50396 575532 50402 575544
rect 473998 575532 474004 575544
rect 50396 575504 474004 575532
rect 50396 575492 50402 575504
rect 473998 575492 474004 575504
rect 474056 575492 474062 575544
rect 54478 575288 54484 575340
rect 54536 575328 54542 575340
rect 395614 575328 395620 575340
rect 54536 575300 395620 575328
rect 54536 575288 54542 575300
rect 395614 575288 395620 575300
rect 395672 575288 395678 575340
rect 207934 575220 207940 575272
rect 207992 575260 207998 575272
rect 580810 575260 580816 575272
rect 207992 575232 580816 575260
rect 207992 575220 207998 575232
rect 580810 575220 580816 575232
rect 580868 575220 580874 575272
rect 3878 575152 3884 575204
rect 3936 575192 3942 575204
rect 379882 575192 379888 575204
rect 3936 575164 379888 575192
rect 3936 575152 3942 575164
rect 379882 575152 379888 575164
rect 379940 575152 379946 575204
rect 203978 575084 203984 575136
rect 204036 575124 204042 575136
rect 580902 575124 580908 575136
rect 204036 575096 580908 575124
rect 204036 575084 204042 575096
rect 580902 575084 580908 575096
rect 580960 575084 580966 575136
rect 3970 575016 3976 575068
rect 4028 575056 4034 575068
rect 383838 575056 383844 575068
rect 4028 575028 383844 575056
rect 4028 575016 4034 575028
rect 383838 575016 383844 575028
rect 383896 575016 383902 575068
rect 391842 575056 391848 575068
rect 391803 575028 391848 575056
rect 391842 575016 391848 575028
rect 391900 575016 391906 575068
rect 403434 575056 403440 575068
rect 403395 575028 403440 575056
rect 403434 575016 403440 575028
rect 403492 575016 403498 575068
rect 415394 575056 415400 575068
rect 415355 575028 415400 575056
rect 415394 575016 415400 575028
rect 415452 575016 415458 575068
rect 438854 575056 438860 575068
rect 438815 575028 438860 575056
rect 438854 575016 438860 575028
rect 438912 575016 438918 575068
rect 450538 575056 450544 575068
rect 450499 575028 450544 575056
rect 450538 575016 450544 575028
rect 450596 575016 450602 575068
rect 462314 575056 462320 575068
rect 462275 575028 462320 575056
rect 462314 575016 462320 575028
rect 462372 575016 462378 575068
rect 195974 574948 195980 575000
rect 196032 574988 196038 575000
rect 580626 574988 580632 575000
rect 196032 574960 580632 574988
rect 196032 574948 196038 574960
rect 580626 574948 580632 574960
rect 580684 574948 580690 575000
rect 109862 574920 109868 574932
rect 109823 574892 109868 574920
rect 109862 574880 109868 574892
rect 109920 574880 109926 574932
rect 117682 574920 117688 574932
rect 117643 574892 117688 574920
rect 117682 574880 117688 574892
rect 117740 574880 117746 574932
rect 145006 574920 145012 574932
rect 144967 574892 145012 574920
rect 145006 574880 145012 574892
rect 145064 574880 145070 574932
rect 164786 574920 164792 574932
rect 164747 574892 164792 574920
rect 164786 574880 164792 574892
rect 164844 574880 164850 574932
rect 176562 574920 176568 574932
rect 176523 574892 176568 574920
rect 176562 574880 176568 574892
rect 176620 574880 176626 574932
rect 180426 574920 180432 574932
rect 180387 574892 180432 574920
rect 180426 574880 180432 574892
rect 180484 574880 180490 574932
rect 192202 574880 192208 574932
rect 192260 574920 192266 574932
rect 580718 574920 580724 574932
rect 192260 574892 580724 574920
rect 192260 574880 192266 574892
rect 580718 574880 580724 574892
rect 580776 574880 580782 574932
rect 3786 574812 3792 574864
rect 3844 574852 3850 574864
rect 391845 574855 391903 574861
rect 391845 574852 391857 574855
rect 3844 574824 391857 574852
rect 3844 574812 3850 574824
rect 391845 574821 391857 574824
rect 391891 574821 391903 574855
rect 391845 574815 391903 574821
rect 58618 574744 58624 574796
rect 58676 574784 58682 574796
rect 450541 574787 450599 574793
rect 450541 574784 450553 574787
rect 58676 574756 450553 574784
rect 58676 574744 58682 574756
rect 450541 574753 450553 574756
rect 450587 574753 450599 574787
rect 450541 574747 450599 574753
rect 3694 574676 3700 574728
rect 3752 574716 3758 574728
rect 403437 574719 403495 574725
rect 403437 574716 403449 574719
rect 3752 574688 403449 574716
rect 3752 574676 3758 574688
rect 403437 574685 403449 574688
rect 403483 574685 403495 574719
rect 403437 574679 403495 574685
rect 180429 574651 180487 574657
rect 180429 574617 180441 574651
rect 180475 574648 180487 574651
rect 580534 574648 580540 574660
rect 180475 574620 580540 574648
rect 180475 574617 180487 574620
rect 180429 574611 180487 574617
rect 580534 574608 580540 574620
rect 580592 574608 580598 574660
rect 145009 574583 145067 574589
rect 145009 574549 145021 574583
rect 145055 574580 145067 574583
rect 547138 574580 547144 574592
rect 145055 574552 547144 574580
rect 145055 574549 145067 574552
rect 145009 574543 145067 574549
rect 547138 574540 547144 574552
rect 547196 574540 547202 574592
rect 176565 574515 176623 574521
rect 176565 574481 176577 574515
rect 176611 574512 176623 574515
rect 580442 574512 580448 574524
rect 176611 574484 580448 574512
rect 176611 574481 176623 574484
rect 176565 574475 176623 574481
rect 580442 574472 580448 574484
rect 580500 574472 580506 574524
rect 3602 574404 3608 574456
rect 3660 574444 3666 574456
rect 415397 574447 415455 574453
rect 415397 574444 415409 574447
rect 3660 574416 415409 574444
rect 3660 574404 3666 574416
rect 415397 574413 415409 574416
rect 415443 574413 415455 574447
rect 415397 574407 415455 574413
rect 164789 574379 164847 574385
rect 164789 574345 164801 574379
rect 164835 574376 164847 574379
rect 580350 574376 580356 574388
rect 164835 574348 580356 574376
rect 164835 574345 164847 574348
rect 164789 574339 164847 574345
rect 580350 574336 580356 574348
rect 580408 574336 580414 574388
rect 109865 574311 109923 574317
rect 109865 574277 109877 574311
rect 109911 574308 109923 574311
rect 540238 574308 540244 574320
rect 109911 574280 540244 574308
rect 109911 574277 109923 574280
rect 109865 574271 109923 574277
rect 540238 574268 540244 574280
rect 540296 574268 540302 574320
rect 3510 574200 3516 574252
rect 3568 574240 3574 574252
rect 438857 574243 438915 574249
rect 438857 574240 438869 574243
rect 3568 574212 438869 574240
rect 3568 574200 3574 574212
rect 438857 574209 438869 574212
rect 438903 574209 438915 574243
rect 438857 574203 438915 574209
rect 3418 574132 3424 574184
rect 3476 574172 3482 574184
rect 462317 574175 462375 574181
rect 462317 574172 462329 574175
rect 3476 574144 462329 574172
rect 3476 574132 3482 574144
rect 462317 574141 462329 574144
rect 462363 574141 462375 574175
rect 462317 574135 462375 574141
rect 117685 574107 117743 574113
rect 117685 574073 117697 574107
rect 117731 574104 117743 574107
rect 580258 574104 580264 574116
rect 117731 574076 580264 574104
rect 117731 574073 117743 574076
rect 117685 574067 117743 574073
rect 580258 574064 580264 574076
rect 580316 574064 580322 574116
rect 519538 564340 519544 564392
rect 519596 564380 519602 564392
rect 580166 564380 580172 564392
rect 519596 564352 580172 564380
rect 519596 564340 519602 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 3234 528504 3240 528556
rect 3292 528544 3298 528556
rect 11698 528544 11704 528556
rect 3292 528516 11704 528544
rect 3292 528504 3298 528516
rect 11698 528504 11704 528516
rect 11756 528504 11762 528556
rect 3326 516060 3332 516112
rect 3384 516100 3390 516112
rect 54478 516100 54484 516112
rect 3384 516072 54484 516100
rect 3384 516060 3390 516072
rect 54478 516060 54484 516072
rect 54536 516060 54542 516112
rect 518158 511912 518164 511964
rect 518216 511952 518222 511964
rect 580166 511952 580172 511964
rect 518216 511924 580172 511952
rect 518216 511912 518222 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 3326 476008 3332 476060
rect 3384 476048 3390 476060
rect 36538 476048 36544 476060
rect 3384 476020 36544 476048
rect 3384 476008 3390 476020
rect 36538 476008 36544 476020
rect 36596 476008 36602 476060
rect 3326 463632 3332 463684
rect 3384 463672 3390 463684
rect 53098 463672 53104 463684
rect 3384 463644 53104 463672
rect 3384 463632 3390 463644
rect 53098 463632 53104 463644
rect 53156 463632 53162 463684
rect 516778 458124 516784 458176
rect 516836 458164 516842 458176
rect 580166 458164 580172 458176
rect 516836 458136 580172 458164
rect 516836 458124 516842 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 25498 423620 25504 423632
rect 3384 423592 25504 423620
rect 3384 423580 3390 423592
rect 25498 423580 25504 423592
rect 25556 423580 25562 423632
rect 538858 419432 538864 419484
rect 538916 419472 538922 419484
rect 579706 419472 579712 419484
rect 538916 419444 579712 419472
rect 538916 419432 538922 419444
rect 579706 419432 579712 419444
rect 579764 419432 579770 419484
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 39298 411244 39304 411256
rect 3384 411216 39304 411244
rect 3384 411204 3390 411216
rect 39298 411204 39304 411216
rect 39356 411204 39362 411256
rect 551278 379448 551284 379500
rect 551336 379488 551342 379500
rect 580166 379488 580172 379500
rect 551336 379460 580172 379488
rect 551336 379448 551342 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 66898 372552 66904 372564
rect 3384 372524 66904 372552
rect 3384 372512 3390 372524
rect 66898 372512 66904 372524
rect 66956 372512 66962 372564
rect 537478 365644 537484 365696
rect 537536 365684 537542 365696
rect 579982 365684 579988 365696
rect 537536 365656 579988 365684
rect 537536 365644 537542 365656
rect 579982 365644 579988 365656
rect 580040 365644 580046 365696
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 4798 358476 4804 358488
rect 2832 358448 4804 358476
rect 2832 358436 2838 358448
rect 4798 358436 4804 358448
rect 4856 358436 4862 358488
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 57238 346372 57244 346384
rect 3384 346344 57244 346372
rect 3384 346332 3390 346344
rect 57238 346332 57244 346344
rect 57296 346332 57302 346384
rect 548518 325592 548524 325644
rect 548576 325632 548582 325644
rect 579890 325632 579896 325644
rect 548576 325604 579896 325632
rect 548576 325592 548582 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 61378 320124 61384 320136
rect 3384 320096 61384 320124
rect 3384 320084 3390 320096
rect 61378 320084 61384 320096
rect 61436 320084 61442 320136
rect 536098 313216 536104 313268
rect 536156 313256 536162 313268
rect 580166 313256 580172 313268
rect 536156 313228 580172 313256
rect 536156 313216 536162 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 14458 306320 14464 306332
rect 3384 306292 14464 306320
rect 3384 306280 3390 306292
rect 14458 306280 14464 306292
rect 14516 306280 14522 306332
rect 525058 299412 525064 299464
rect 525116 299452 525122 299464
rect 579614 299452 579620 299464
rect 525116 299424 579620 299452
rect 525116 299412 525122 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 547138 273164 547144 273216
rect 547196 273204 547202 273216
rect 579890 273204 579896 273216
rect 547196 273176 579896 273204
rect 547196 273164 547202 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 65518 267696 65524 267708
rect 3568 267668 65524 267696
rect 3568 267656 3574 267668
rect 65518 267656 65524 267668
rect 65576 267656 65582 267708
rect 533338 259360 533344 259412
rect 533396 259400 533402 259412
rect 579798 259400 579804 259412
rect 533396 259372 579804 259400
rect 533396 259360 533402 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 17218 255252 17224 255264
rect 3200 255224 17224 255252
rect 3200 255212 3206 255224
rect 17218 255212 17224 255224
rect 17276 255212 17282 255264
rect 522298 245556 522304 245608
rect 522356 245596 522362 245608
rect 580166 245596 580172 245608
rect 522356 245568 580172 245596
rect 522356 245556 522362 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 58618 241448 58624 241460
rect 3568 241420 58624 241448
rect 3568 241408 3574 241420
rect 58618 241408 58624 241420
rect 58676 241408 58682 241460
rect 544378 233180 544384 233232
rect 544436 233220 544442 233232
rect 580166 233220 580172 233232
rect 544436 233192 580172 233220
rect 544436 233180 544442 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 530578 219376 530584 219428
rect 530636 219416 530642 219428
rect 579890 219416 579896 219428
rect 530636 219388 579896 219416
rect 530636 219376 530642 219388
rect 579890 219376 579896 219388
rect 579948 219376 579954 219428
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 47578 215268 47584 215280
rect 3384 215240 47584 215268
rect 3384 215228 3390 215240
rect 47578 215228 47584 215240
rect 47636 215228 47642 215280
rect 520918 206932 520924 206984
rect 520976 206972 520982 206984
rect 580166 206972 580172 206984
rect 520976 206944 580172 206972
rect 520976 206932 520982 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 18598 202824 18604 202836
rect 3108 202796 18604 202824
rect 3108 202784 3114 202796
rect 18598 202784 18604 202796
rect 18656 202784 18662 202836
rect 542998 193128 543004 193180
rect 543056 193168 543062 193180
rect 580166 193168 580172 193180
rect 543056 193140 580172 193168
rect 543056 193128 543062 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 529198 179324 529204 179376
rect 529256 179364 529262 179376
rect 579982 179364 579988 179376
rect 529256 179336 579988 179364
rect 529256 179324 529262 179336
rect 579982 179324 579988 179336
rect 580040 179324 580046 179376
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 51718 164200 51724 164212
rect 3292 164172 51724 164200
rect 3292 164160 3298 164172
rect 51718 164160 51724 164172
rect 51776 164160 51782 164212
rect 540238 153144 540244 153196
rect 540296 153184 540302 153196
rect 580166 153184 580172 153196
rect 540296 153156 580172 153184
rect 540296 153144 540302 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 21358 150396 21364 150408
rect 3476 150368 21364 150396
rect 3476 150356 3482 150368
rect 21358 150356 21364 150368
rect 21416 150356 21422 150408
rect 526438 139340 526444 139392
rect 526496 139380 526502 139392
rect 580166 139380 580172 139392
rect 526496 139352 580172 139380
rect 526496 139340 526502 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 50338 137952 50344 137964
rect 3292 137924 50344 137952
rect 3292 137912 3298 137924
rect 50338 137912 50344 137924
rect 50396 137912 50402 137964
rect 93854 128188 93860 128240
rect 93912 128228 93918 128240
rect 95004 128228 95010 128240
rect 93912 128200 95010 128228
rect 93912 128188 93918 128200
rect 95004 128188 95010 128200
rect 95062 128188 95068 128240
rect 125686 128188 125692 128240
rect 125744 128228 125750 128240
rect 126836 128228 126842 128240
rect 125744 128200 126842 128228
rect 125744 128188 125750 128200
rect 126836 128188 126842 128200
rect 126894 128188 126900 128240
rect 146294 128188 146300 128240
rect 146352 128228 146358 128240
rect 147628 128228 147634 128240
rect 146352 128200 147634 128228
rect 146352 128188 146358 128200
rect 147628 128188 147634 128200
rect 147686 128188 147692 128240
rect 149054 128188 149060 128240
rect 149112 128228 149118 128240
rect 150388 128228 150394 128240
rect 149112 128200 150394 128228
rect 149112 128188 149118 128200
rect 150388 128188 150394 128200
rect 150446 128188 150452 128240
rect 157426 128188 157432 128240
rect 157484 128228 157490 128240
rect 158576 128228 158582 128240
rect 157484 128200 158582 128228
rect 157484 128188 157490 128200
rect 158576 128188 158582 128200
rect 158634 128188 158640 128240
rect 186406 128188 186412 128240
rect 186464 128228 186470 128240
rect 187556 128228 187562 128240
rect 186464 128200 187562 128228
rect 186464 128188 186470 128200
rect 187556 128188 187562 128200
rect 187614 128188 187620 128240
rect 212626 128188 212632 128240
rect 212684 128228 212690 128240
rect 213868 128228 213874 128240
rect 212684 128200 213874 128228
rect 212684 128188 212690 128200
rect 213868 128188 213874 128200
rect 213926 128188 213932 128240
rect 215386 128188 215392 128240
rect 215444 128228 215450 128240
rect 216628 128228 216634 128240
rect 215444 128200 216634 128228
rect 215444 128188 215450 128200
rect 216628 128188 216634 128200
rect 216686 128188 216692 128240
rect 218146 128188 218152 128240
rect 218204 128228 218210 128240
rect 219296 128228 219302 128240
rect 218204 128200 219302 128228
rect 218204 128188 218210 128200
rect 219296 128188 219302 128200
rect 219354 128188 219360 128240
rect 220906 128188 220912 128240
rect 220964 128228 220970 128240
rect 222056 128228 222062 128240
rect 220964 128200 222062 128228
rect 220964 128188 220970 128200
rect 222056 128188 222062 128200
rect 222114 128188 222120 128240
rect 287146 128188 287152 128240
rect 287204 128228 287210 128240
rect 288296 128228 288302 128240
rect 287204 128200 288302 128228
rect 287204 128188 287210 128200
rect 288296 128188 288302 128200
rect 288354 128188 288360 128240
rect 64782 126896 64788 126948
rect 64840 126936 64846 126948
rect 117682 126936 117688 126948
rect 64840 126908 117688 126936
rect 64840 126896 64846 126908
rect 117682 126896 117688 126908
rect 117740 126896 117746 126948
rect 122098 126896 122104 126948
rect 122156 126936 122162 126948
rect 124030 126936 124036 126948
rect 122156 126908 124036 126936
rect 122156 126896 122162 126908
rect 124030 126896 124036 126908
rect 124088 126896 124094 126948
rect 125502 126896 125508 126948
rect 125560 126936 125566 126948
rect 163958 126936 163964 126948
rect 125560 126908 163964 126936
rect 125560 126896 125566 126908
rect 163958 126896 163964 126908
rect 164016 126896 164022 126948
rect 170398 126896 170404 126948
rect 170456 126936 170462 126948
rect 172146 126936 172152 126948
rect 170456 126908 172152 126936
rect 170456 126896 170462 126908
rect 172146 126896 172152 126908
rect 172204 126896 172210 126948
rect 175921 126939 175979 126945
rect 175921 126905 175933 126939
rect 175967 126936 175979 126939
rect 199286 126936 199292 126948
rect 175967 126908 199292 126936
rect 175967 126905 175979 126908
rect 175921 126899 175979 126905
rect 199286 126896 199292 126908
rect 199344 126896 199350 126948
rect 200022 126896 200028 126948
rect 200080 126936 200086 126948
rect 221090 126936 221096 126948
rect 200080 126908 221096 126936
rect 200080 126896 200086 126908
rect 221090 126896 221096 126908
rect 221148 126896 221154 126948
rect 223482 126896 223488 126948
rect 223540 126936 223546 126948
rect 239214 126936 239220 126948
rect 223540 126908 239220 126936
rect 223540 126896 223546 126908
rect 239214 126896 239220 126908
rect 239272 126896 239278 126948
rect 276658 126896 276664 126948
rect 276716 126936 276722 126948
rect 279142 126936 279148 126948
rect 276716 126908 279148 126936
rect 276716 126896 276722 126908
rect 279142 126896 279148 126908
rect 279200 126896 279206 126948
rect 344554 126896 344560 126948
rect 344612 126936 344618 126948
rect 345658 126936 345664 126948
rect 344612 126908 345664 126936
rect 344612 126896 344618 126908
rect 345658 126896 345664 126908
rect 345716 126896 345722 126948
rect 401686 126896 401692 126948
rect 401744 126936 401750 126948
rect 403618 126936 403624 126948
rect 401744 126908 403624 126936
rect 401744 126896 401750 126908
rect 403618 126896 403624 126908
rect 403676 126896 403682 126948
rect 472434 126896 472440 126948
rect 472492 126936 472498 126948
rect 472492 126908 518894 126936
rect 472492 126896 472498 126908
rect 56502 126828 56508 126880
rect 56560 126868 56566 126880
rect 111334 126868 111340 126880
rect 56560 126840 111340 126868
rect 56560 126828 56566 126840
rect 111334 126828 111340 126840
rect 111392 126828 111398 126880
rect 112530 126828 112536 126880
rect 112588 126868 112594 126880
rect 113174 126868 113180 126880
rect 112588 126840 113180 126868
rect 112588 126828 112594 126840
rect 113174 126828 113180 126840
rect 113232 126828 113238 126880
rect 126238 126828 126244 126880
rect 126296 126868 126302 126880
rect 145834 126868 145840 126880
rect 126296 126840 145840 126868
rect 126296 126828 126302 126840
rect 145834 126828 145840 126840
rect 145892 126828 145898 126880
rect 160002 126828 160008 126880
rect 160060 126868 160066 126880
rect 190270 126868 190276 126880
rect 160060 126840 190276 126868
rect 160060 126828 160066 126840
rect 190270 126828 190276 126840
rect 190328 126828 190334 126880
rect 195238 126828 195244 126880
rect 195296 126868 195302 126880
rect 217502 126868 217508 126880
rect 195296 126840 217508 126868
rect 195296 126828 195302 126840
rect 217502 126828 217508 126840
rect 217560 126828 217566 126880
rect 220078 126828 220084 126880
rect 220136 126868 220142 126880
rect 236546 126868 236552 126880
rect 220136 126840 236552 126868
rect 220136 126828 220142 126840
rect 236546 126828 236552 126840
rect 236604 126828 236610 126880
rect 238018 126828 238024 126880
rect 238076 126868 238082 126880
rect 242894 126868 242900 126880
rect 238076 126840 242900 126868
rect 238076 126828 238082 126840
rect 242894 126828 242900 126840
rect 242952 126828 242958 126880
rect 246298 126828 246304 126880
rect 246356 126868 246362 126880
rect 251910 126868 251916 126880
rect 246356 126840 251916 126868
rect 246356 126828 246362 126840
rect 251910 126828 251916 126840
rect 251968 126828 251974 126880
rect 312814 126828 312820 126880
rect 312872 126868 312878 126880
rect 317414 126868 317420 126880
rect 312872 126840 317420 126868
rect 312872 126828 312878 126840
rect 317414 126828 317420 126840
rect 317472 126828 317478 126880
rect 469766 126828 469772 126880
rect 469824 126868 469830 126880
rect 514021 126871 514079 126877
rect 514021 126868 514033 126871
rect 469824 126840 514033 126868
rect 469824 126828 469830 126840
rect 514021 126837 514033 126840
rect 514067 126837 514079 126871
rect 518866 126868 518894 126908
rect 519538 126868 519544 126880
rect 518866 126840 519544 126868
rect 514021 126831 514079 126837
rect 519538 126828 519544 126840
rect 519596 126828 519602 126880
rect 57882 126760 57888 126812
rect 57940 126800 57946 126812
rect 112254 126800 112260 126812
rect 57940 126772 112260 126800
rect 57940 126760 57946 126772
rect 112254 126760 112260 126772
rect 112312 126760 112318 126812
rect 112438 126760 112444 126812
rect 112496 126800 112502 126812
rect 121270 126800 121276 126812
rect 112496 126772 121276 126800
rect 112496 126760 112502 126772
rect 121270 126760 121276 126772
rect 121328 126760 121334 126812
rect 124122 126760 124128 126812
rect 124180 126800 124186 126812
rect 163038 126800 163044 126812
rect 124180 126772 163044 126800
rect 124180 126760 124186 126772
rect 163038 126760 163044 126772
rect 163096 126760 163102 126812
rect 171042 126760 171048 126812
rect 171100 126800 171106 126812
rect 175921 126803 175979 126809
rect 175921 126800 175933 126803
rect 171100 126772 175933 126800
rect 171100 126760 171106 126772
rect 175921 126769 175933 126772
rect 175967 126769 175979 126803
rect 175921 126763 175979 126769
rect 176013 126803 176071 126809
rect 176013 126769 176025 126803
rect 176059 126800 176071 126803
rect 198366 126800 198372 126812
rect 176059 126772 198372 126800
rect 176059 126769 176071 126772
rect 176013 126763 176071 126769
rect 198366 126760 198372 126772
rect 198424 126760 198430 126812
rect 202690 126760 202696 126812
rect 202748 126800 202754 126812
rect 223850 126800 223856 126812
rect 202748 126772 223856 126800
rect 202748 126760 202754 126772
rect 223850 126760 223856 126772
rect 223908 126760 223914 126812
rect 224862 126760 224868 126812
rect 224920 126800 224926 126812
rect 240134 126800 240140 126812
rect 224920 126772 240140 126800
rect 224920 126760 224926 126772
rect 240134 126760 240140 126772
rect 240192 126760 240198 126812
rect 242802 126760 242808 126812
rect 242860 126800 242866 126812
rect 253750 126800 253756 126812
rect 242860 126772 253756 126800
rect 242860 126760 242866 126772
rect 253750 126760 253756 126772
rect 253808 126760 253814 126812
rect 256602 126760 256608 126812
rect 256660 126800 256666 126812
rect 264606 126800 264612 126812
rect 256660 126772 264612 126800
rect 256660 126760 256666 126772
rect 264606 126760 264612 126772
rect 264664 126760 264670 126812
rect 285582 126760 285588 126812
rect 285640 126800 285646 126812
rect 287330 126800 287336 126812
rect 285640 126772 287336 126800
rect 285640 126760 285646 126772
rect 287330 126760 287336 126772
rect 287388 126760 287394 126812
rect 440694 126760 440700 126812
rect 440752 126800 440758 126812
rect 450538 126800 450544 126812
rect 440752 126772 450544 126800
rect 440752 126760 440758 126772
rect 450538 126760 450544 126772
rect 450596 126760 450602 126812
rect 466086 126760 466092 126812
rect 466144 126800 466150 126812
rect 517514 126800 517520 126812
rect 466144 126772 517520 126800
rect 466144 126760 466150 126772
rect 517514 126760 517520 126772
rect 517572 126760 517578 126812
rect 29638 126692 29644 126744
rect 29696 126732 29702 126744
rect 89530 126732 89536 126744
rect 29696 126704 89536 126732
rect 29696 126692 29702 126704
rect 89530 126692 89536 126704
rect 89588 126692 89594 126744
rect 117222 126692 117228 126744
rect 117280 126732 117286 126744
rect 157610 126732 157616 126744
rect 117280 126704 157616 126732
rect 117280 126692 117286 126704
rect 157610 126692 157616 126704
rect 157668 126692 157674 126744
rect 162762 126692 162768 126744
rect 162820 126732 162826 126744
rect 192938 126732 192944 126744
rect 162820 126704 192944 126732
rect 162820 126692 162826 126704
rect 192938 126692 192944 126704
rect 192996 126692 193002 126744
rect 193122 126692 193128 126744
rect 193180 126732 193186 126744
rect 215662 126732 215668 126744
rect 193180 126704 215668 126732
rect 193180 126692 193186 126704
rect 215662 126692 215668 126704
rect 215720 126692 215726 126744
rect 216582 126692 216588 126744
rect 216640 126732 216646 126744
rect 233786 126732 233792 126744
rect 216640 126704 233792 126732
rect 216640 126692 216646 126704
rect 233786 126692 233792 126704
rect 233844 126692 233850 126744
rect 238662 126692 238668 126744
rect 238720 126732 238726 126744
rect 250990 126732 250996 126744
rect 238720 126704 250996 126732
rect 238720 126692 238726 126704
rect 250990 126692 250996 126704
rect 251048 126692 251054 126744
rect 253198 126692 253204 126744
rect 253256 126732 253262 126744
rect 261938 126732 261944 126744
rect 253256 126704 261944 126732
rect 253256 126692 253262 126704
rect 261938 126692 261944 126704
rect 261996 126692 262002 126744
rect 448882 126692 448888 126744
rect 448940 126732 448946 126744
rect 448940 126704 471468 126732
rect 448940 126692 448946 126704
rect 14458 126624 14464 126676
rect 14516 126664 14522 126676
rect 73246 126664 73252 126676
rect 14516 126636 73252 126664
rect 14516 126624 14522 126636
rect 73246 126624 73252 126636
rect 73304 126624 73310 126676
rect 78490 126624 78496 126676
rect 78548 126664 78554 126676
rect 127618 126664 127624 126676
rect 78548 126636 127624 126664
rect 78548 126624 78554 126636
rect 127618 126624 127624 126636
rect 127676 126624 127682 126676
rect 152550 126624 152556 126676
rect 152608 126664 152614 126676
rect 153930 126664 153936 126676
rect 152608 126636 153936 126664
rect 152608 126624 152614 126636
rect 153930 126624 153936 126636
rect 153988 126624 153994 126676
rect 158622 126624 158628 126676
rect 158680 126664 158686 126676
rect 189350 126664 189356 126676
rect 158680 126636 189356 126664
rect 158680 126624 158686 126636
rect 189350 126624 189356 126636
rect 189408 126624 189414 126676
rect 191742 126624 191748 126676
rect 191800 126664 191806 126676
rect 214742 126664 214748 126676
rect 191800 126636 214748 126664
rect 191800 126624 191806 126636
rect 214742 126624 214748 126636
rect 214800 126624 214806 126676
rect 217962 126624 217968 126676
rect 218020 126664 218026 126676
rect 234706 126664 234712 126676
rect 218020 126636 234712 126664
rect 218020 126624 218026 126636
rect 234706 126624 234712 126636
rect 234764 126624 234770 126676
rect 235902 126624 235908 126676
rect 235960 126664 235966 126676
rect 249242 126664 249248 126676
rect 235960 126636 249248 126664
rect 235960 126624 235966 126636
rect 249242 126624 249248 126636
rect 249300 126624 249306 126676
rect 250438 126624 250444 126676
rect 250496 126664 250502 126676
rect 259178 126664 259184 126676
rect 250496 126636 259184 126664
rect 250496 126624 250502 126636
rect 259178 126624 259184 126636
rect 259236 126624 259242 126676
rect 415302 126624 415308 126676
rect 415360 126664 415366 126676
rect 442258 126664 442264 126676
rect 415360 126636 442264 126664
rect 415360 126624 415366 126636
rect 442258 126624 442264 126636
rect 442316 126624 442322 126676
rect 457070 126624 457076 126676
rect 457128 126664 457134 126676
rect 464338 126664 464344 126676
rect 457128 126636 464344 126664
rect 457128 126624 457134 126636
rect 464338 126624 464344 126636
rect 464396 126624 464402 126676
rect 22738 126556 22744 126608
rect 22796 126596 22802 126608
rect 84102 126596 84108 126608
rect 22796 126568 84108 126596
rect 22796 126556 22802 126568
rect 84102 126556 84108 126568
rect 84160 126556 84166 126608
rect 111702 126556 111708 126608
rect 111760 126596 111766 126608
rect 153010 126596 153016 126608
rect 111760 126568 153016 126596
rect 111760 126556 111766 126568
rect 153010 126556 153016 126568
rect 153068 126556 153074 126608
rect 153102 126556 153108 126608
rect 153160 126596 153166 126608
rect 185670 126596 185676 126608
rect 153160 126568 185676 126596
rect 153160 126556 153166 126568
rect 185670 126556 185676 126568
rect 185728 126556 185734 126608
rect 188982 126556 188988 126608
rect 189040 126596 189046 126608
rect 212902 126596 212908 126608
rect 189040 126568 212908 126596
rect 189040 126556 189046 126568
rect 212902 126556 212908 126568
rect 212960 126556 212966 126608
rect 213822 126556 213828 126608
rect 213880 126596 213886 126608
rect 231946 126596 231952 126608
rect 213880 126568 231952 126596
rect 213880 126556 213886 126568
rect 231946 126556 231952 126568
rect 232004 126556 232010 126608
rect 237282 126556 237288 126608
rect 237340 126596 237346 126608
rect 250162 126596 250168 126608
rect 237340 126568 250168 126596
rect 237340 126556 237346 126568
rect 250162 126556 250168 126568
rect 250220 126556 250226 126608
rect 252462 126556 252468 126608
rect 252520 126596 252526 126608
rect 261018 126596 261024 126608
rect 252520 126568 261024 126596
rect 252520 126556 252526 126568
rect 261018 126556 261024 126568
rect 261076 126556 261082 126608
rect 420730 126556 420736 126608
rect 420788 126596 420794 126608
rect 432598 126596 432604 126608
rect 420788 126568 432604 126596
rect 420788 126556 420794 126568
rect 432598 126556 432604 126568
rect 432656 126556 432662 126608
rect 437106 126556 437112 126608
rect 437164 126596 437170 126608
rect 471330 126596 471336 126608
rect 437164 126568 471336 126596
rect 437164 126556 437170 126568
rect 471330 126556 471336 126568
rect 471388 126556 471394 126608
rect 471440 126596 471468 126704
rect 477034 126692 477040 126744
rect 477092 126732 477098 126744
rect 484765 126735 484823 126741
rect 484765 126732 484777 126735
rect 477092 126704 484777 126732
rect 477092 126692 477098 126704
rect 484765 126701 484777 126704
rect 484811 126701 484823 126735
rect 484765 126695 484823 126701
rect 493045 126735 493103 126741
rect 493045 126701 493057 126735
rect 493091 126732 493103 126735
rect 536098 126732 536104 126744
rect 493091 126704 536104 126732
rect 493091 126701 493103 126704
rect 493045 126695 493103 126701
rect 536098 126692 536104 126704
rect 536156 126692 536162 126744
rect 471514 126624 471520 126676
rect 471572 126664 471578 126676
rect 524414 126664 524420 126676
rect 471572 126636 524420 126664
rect 471572 126624 471578 126636
rect 524414 126624 524420 126636
rect 524472 126624 524478 126676
rect 479518 126596 479524 126608
rect 471440 126568 479524 126596
rect 479518 126556 479524 126568
rect 479576 126556 479582 126608
rect 484765 126599 484823 126605
rect 484765 126565 484777 126599
rect 484811 126596 484823 126599
rect 531314 126596 531320 126608
rect 484811 126568 531320 126596
rect 484811 126565 484823 126568
rect 484765 126559 484823 126565
rect 531314 126556 531320 126568
rect 531372 126556 531378 126608
rect 25498 126488 25504 126540
rect 25556 126528 25562 126540
rect 86862 126528 86868 126540
rect 25556 126500 86868 126528
rect 25556 126488 25562 126500
rect 86862 126488 86868 126500
rect 86920 126488 86926 126540
rect 88242 126488 88248 126540
rect 88300 126528 88306 126540
rect 99558 126528 99564 126540
rect 88300 126500 99564 126528
rect 88300 126488 88306 126500
rect 99558 126488 99564 126500
rect 99616 126488 99622 126540
rect 104802 126488 104808 126540
rect 104860 126528 104866 126540
rect 148502 126528 148508 126540
rect 104860 126500 148508 126528
rect 104860 126488 104866 126500
rect 148502 126488 148508 126500
rect 148560 126488 148566 126540
rect 148962 126488 148968 126540
rect 149020 126528 149026 126540
rect 182082 126528 182088 126540
rect 149020 126500 182088 126528
rect 149020 126488 149026 126500
rect 182082 126488 182088 126500
rect 182140 126488 182146 126540
rect 187602 126488 187608 126540
rect 187660 126528 187666 126540
rect 187660 126500 209452 126528
rect 187660 126488 187666 126500
rect 21358 126420 21364 126472
rect 21416 126460 21422 126472
rect 82262 126460 82268 126472
rect 21416 126432 82268 126460
rect 21416 126420 21422 126432
rect 82262 126420 82268 126432
rect 82320 126420 82326 126472
rect 88978 126420 88984 126472
rect 89036 126460 89042 126472
rect 96614 126460 96620 126472
rect 89036 126432 96620 126460
rect 89036 126420 89042 126432
rect 96614 126420 96620 126432
rect 96672 126420 96678 126472
rect 99282 126420 99288 126472
rect 99340 126460 99346 126472
rect 143994 126460 144000 126472
rect 99340 126432 144000 126460
rect 99340 126420 99346 126432
rect 143994 126420 144000 126432
rect 144052 126420 144058 126472
rect 144822 126420 144828 126472
rect 144880 126460 144886 126472
rect 179322 126460 179328 126472
rect 144880 126432 179328 126460
rect 144880 126420 144886 126432
rect 179322 126420 179328 126432
rect 179380 126420 179386 126472
rect 184750 126420 184756 126472
rect 184808 126460 184814 126472
rect 209314 126460 209320 126472
rect 184808 126432 209320 126460
rect 184808 126420 184814 126432
rect 209314 126420 209320 126432
rect 209372 126420 209378 126472
rect 17218 126352 17224 126404
rect 17276 126392 17282 126404
rect 79594 126392 79600 126404
rect 17276 126364 79600 126392
rect 17276 126352 17282 126364
rect 79594 126352 79600 126364
rect 79652 126352 79658 126404
rect 93762 126352 93768 126404
rect 93820 126392 93826 126404
rect 139486 126392 139492 126404
rect 93820 126364 139492 126392
rect 93820 126352 93826 126364
rect 139486 126352 139492 126364
rect 139544 126352 139550 126404
rect 142062 126352 142068 126404
rect 142120 126392 142126 126404
rect 176654 126392 176660 126404
rect 142120 126364 176660 126392
rect 142120 126352 142126 126364
rect 176654 126352 176660 126364
rect 176712 126352 176718 126404
rect 177942 126352 177948 126404
rect 178000 126392 178006 126404
rect 203886 126392 203892 126404
rect 178000 126364 203892 126392
rect 178000 126352 178006 126364
rect 203886 126352 203892 126364
rect 203944 126352 203950 126404
rect 209424 126392 209452 126500
rect 212442 126488 212448 126540
rect 212500 126528 212506 126540
rect 231026 126528 231032 126540
rect 212500 126500 231032 126528
rect 212500 126488 212506 126500
rect 231026 126488 231032 126500
rect 231084 126488 231090 126540
rect 234522 126488 234528 126540
rect 234580 126528 234586 126540
rect 247402 126528 247408 126540
rect 234580 126500 247408 126528
rect 234580 126488 234586 126500
rect 247402 126488 247408 126500
rect 247460 126488 247466 126540
rect 249058 126488 249064 126540
rect 249116 126528 249122 126540
rect 258258 126528 258264 126540
rect 249116 126500 258264 126528
rect 249116 126488 249122 126500
rect 258258 126488 258264 126500
rect 258316 126488 258322 126540
rect 267642 126488 267648 126540
rect 267700 126528 267706 126540
rect 272794 126528 272800 126540
rect 267700 126500 272800 126528
rect 267700 126488 267706 126500
rect 272794 126488 272800 126500
rect 272852 126488 272858 126540
rect 399018 126488 399024 126540
rect 399076 126528 399082 126540
rect 418798 126528 418804 126540
rect 399076 126500 418804 126528
rect 399076 126488 399082 126500
rect 418798 126488 418804 126500
rect 418856 126488 418862 126540
rect 419810 126488 419816 126540
rect 419868 126528 419874 126540
rect 456886 126528 456892 126540
rect 419868 126500 456892 126528
rect 419868 126488 419874 126500
rect 456886 126488 456892 126500
rect 456944 126488 456950 126540
rect 459738 126488 459744 126540
rect 459796 126528 459802 126540
rect 471238 126528 471244 126540
rect 459796 126500 471244 126528
rect 459796 126488 459802 126500
rect 471238 126488 471244 126500
rect 471296 126488 471302 126540
rect 478782 126488 478788 126540
rect 478840 126528 478846 126540
rect 533338 126528 533344 126540
rect 478840 126500 533344 126528
rect 478840 126488 478846 126500
rect 533338 126488 533344 126500
rect 533396 126488 533402 126540
rect 209682 126420 209688 126472
rect 209740 126460 209746 126472
rect 228358 126460 228364 126472
rect 209740 126432 228364 126460
rect 209740 126420 209746 126432
rect 228358 126420 228364 126432
rect 228416 126420 228422 126472
rect 231118 126420 231124 126472
rect 231176 126460 231182 126472
rect 244642 126460 244648 126472
rect 231176 126432 244648 126460
rect 231176 126420 231182 126432
rect 244642 126420 244648 126432
rect 244700 126420 244706 126472
rect 246942 126420 246948 126472
rect 247000 126460 247006 126472
rect 257338 126460 257344 126472
rect 247000 126432 257344 126460
rect 247000 126420 247006 126432
rect 257338 126420 257344 126432
rect 257396 126420 257402 126472
rect 409782 126420 409788 126472
rect 409840 126460 409846 126472
rect 429746 126460 429752 126472
rect 409840 126432 429752 126460
rect 409840 126420 409846 126432
rect 429746 126420 429752 126432
rect 429804 126420 429810 126472
rect 434346 126420 434352 126472
rect 434404 126460 434410 126472
rect 465721 126463 465779 126469
rect 465721 126460 465733 126463
rect 434404 126432 465733 126460
rect 434404 126420 434410 126432
rect 465721 126429 465733 126432
rect 465767 126429 465779 126463
rect 465721 126423 465779 126429
rect 484210 126420 484216 126472
rect 484268 126460 484274 126472
rect 493045 126463 493103 126469
rect 493045 126460 493057 126463
rect 484268 126432 493057 126460
rect 484268 126420 484274 126432
rect 493045 126429 493057 126432
rect 493091 126429 493103 126463
rect 493045 126423 493103 126429
rect 495989 126463 496047 126469
rect 495989 126429 496001 126463
rect 496035 126460 496047 126463
rect 547138 126460 547144 126472
rect 496035 126432 547144 126460
rect 496035 126429 496047 126432
rect 495989 126423 496047 126429
rect 547138 126420 547144 126432
rect 547196 126420 547202 126472
rect 211982 126392 211988 126404
rect 209424 126364 211988 126392
rect 211982 126352 211988 126364
rect 212040 126352 212046 126404
rect 214561 126395 214619 126401
rect 214561 126361 214573 126395
rect 214607 126392 214619 126395
rect 225598 126392 225604 126404
rect 214607 126364 225604 126392
rect 214607 126361 214619 126364
rect 214561 126355 214619 126361
rect 225598 126352 225604 126364
rect 225656 126352 225662 126404
rect 229002 126352 229008 126404
rect 229060 126392 229066 126404
rect 243722 126392 243728 126404
rect 229060 126364 243728 126392
rect 229060 126352 229066 126364
rect 243722 126352 243728 126364
rect 243780 126352 243786 126404
rect 245562 126352 245568 126404
rect 245620 126392 245626 126404
rect 256510 126392 256516 126404
rect 245620 126364 256516 126392
rect 245620 126352 245626 126364
rect 256510 126352 256516 126364
rect 256568 126352 256574 126404
rect 260742 126352 260748 126404
rect 260800 126392 260806 126404
rect 268286 126392 268292 126404
rect 260800 126364 268292 126392
rect 260800 126352 260806 126364
rect 268286 126352 268292 126364
rect 268344 126352 268350 126404
rect 332778 126352 332784 126404
rect 332836 126392 332842 126404
rect 335998 126392 336004 126404
rect 332836 126364 336004 126392
rect 332836 126352 332842 126364
rect 335998 126352 336004 126364
rect 336056 126352 336062 126404
rect 388070 126352 388076 126404
rect 388128 126392 388134 126404
rect 407758 126392 407764 126404
rect 388128 126364 407764 126392
rect 388128 126352 388134 126364
rect 407758 126352 407764 126364
rect 407816 126352 407822 126404
rect 428918 126352 428924 126404
rect 428976 126392 428982 126404
rect 467098 126392 467104 126404
rect 428976 126364 467104 126392
rect 428976 126352 428982 126364
rect 467098 126352 467104 126364
rect 467156 126352 467162 126404
rect 486970 126352 486976 126404
rect 487028 126392 487034 126404
rect 542998 126392 543004 126404
rect 487028 126364 543004 126392
rect 487028 126352 487034 126364
rect 542998 126352 543004 126364
rect 543056 126352 543062 126404
rect 7558 126284 7564 126336
rect 7616 126324 7622 126336
rect 72326 126324 72332 126336
rect 7616 126296 72332 126324
rect 7616 126284 7622 126296
rect 72326 126284 72332 126296
rect 72384 126284 72390 126336
rect 75822 126284 75828 126336
rect 75880 126324 75886 126336
rect 125870 126324 125876 126336
rect 75880 126296 125876 126324
rect 75880 126284 75886 126296
rect 125870 126284 125876 126296
rect 125928 126284 125934 126336
rect 130378 126284 130384 126336
rect 130436 126324 130442 126336
rect 165614 126324 165620 126336
rect 130436 126296 165620 126324
rect 130436 126284 130442 126296
rect 165614 126284 165620 126296
rect 165672 126284 165678 126336
rect 166902 126284 166908 126336
rect 166960 126324 166966 126336
rect 195698 126324 195704 126336
rect 166960 126296 195704 126324
rect 166960 126284 166966 126296
rect 195698 126284 195704 126296
rect 195756 126284 195762 126336
rect 195882 126284 195888 126336
rect 195940 126324 195946 126336
rect 218330 126324 218336 126336
rect 195940 126296 218336 126324
rect 195940 126284 195946 126296
rect 218330 126284 218336 126296
rect 218388 126284 218394 126336
rect 220722 126284 220728 126336
rect 220780 126324 220786 126336
rect 237374 126324 237380 126336
rect 220780 126296 237380 126324
rect 220780 126284 220786 126296
rect 237374 126284 237380 126296
rect 237432 126284 237438 126336
rect 241422 126284 241428 126336
rect 241480 126324 241486 126336
rect 252830 126324 252836 126336
rect 241480 126296 252836 126324
rect 241480 126284 241486 126296
rect 252830 126284 252836 126296
rect 252888 126284 252894 126336
rect 255222 126284 255228 126336
rect 255280 126324 255286 126336
rect 263686 126324 263692 126336
rect 255280 126296 263692 126324
rect 255280 126284 255286 126296
rect 263686 126284 263692 126296
rect 263744 126284 263750 126336
rect 350902 126284 350908 126336
rect 350960 126324 350966 126336
rect 359458 126324 359464 126336
rect 350960 126296 359464 126324
rect 350960 126284 350966 126296
rect 359458 126284 359464 126296
rect 359516 126284 359522 126336
rect 377214 126284 377220 126336
rect 377272 126324 377278 126336
rect 389818 126324 389824 126336
rect 377272 126296 389824 126324
rect 377272 126284 377278 126296
rect 389818 126284 389824 126296
rect 389876 126284 389882 126336
rect 393498 126284 393504 126336
rect 393556 126324 393562 126336
rect 421558 126324 421564 126336
rect 393556 126296 421564 126324
rect 393556 126284 393562 126296
rect 421558 126284 421564 126296
rect 421616 126284 421622 126336
rect 423490 126284 423496 126336
rect 423548 126324 423554 126336
rect 461486 126324 461492 126336
rect 423548 126296 461492 126324
rect 423548 126284 423554 126296
rect 461486 126284 461492 126296
rect 461544 126284 461550 126336
rect 470502 126284 470508 126336
rect 470560 126324 470566 126336
rect 475378 126324 475384 126336
rect 470560 126296 475384 126324
rect 470560 126284 470566 126296
rect 475378 126284 475384 126296
rect 475436 126284 475442 126336
rect 482462 126284 482468 126336
rect 482520 126324 482526 126336
rect 539594 126324 539600 126336
rect 482520 126296 539600 126324
rect 482520 126284 482526 126296
rect 539594 126284 539600 126296
rect 539652 126284 539658 126336
rect 11698 126216 11704 126268
rect 11756 126256 11762 126268
rect 75914 126256 75920 126268
rect 11756 126228 75920 126256
rect 11756 126216 11762 126228
rect 75914 126216 75920 126228
rect 75972 126216 75978 126268
rect 78582 126216 78588 126268
rect 78640 126256 78646 126268
rect 128354 126256 128360 126268
rect 78640 126228 128360 126256
rect 78640 126216 78646 126228
rect 128354 126216 128360 126228
rect 128412 126216 128418 126268
rect 137922 126216 137928 126268
rect 137980 126256 137986 126268
rect 173894 126256 173900 126268
rect 137980 126228 173900 126256
rect 137980 126216 137986 126228
rect 173894 126216 173900 126228
rect 173952 126216 173958 126268
rect 180702 126216 180708 126268
rect 180760 126256 180766 126268
rect 206554 126256 206560 126268
rect 180760 126228 206560 126256
rect 180760 126216 180766 126228
rect 206554 126216 206560 126228
rect 206612 126216 206618 126268
rect 206922 126216 206928 126268
rect 206980 126256 206986 126268
rect 226518 126256 226524 126268
rect 206980 126228 226524 126256
rect 206980 126216 206986 126228
rect 226518 126216 226524 126228
rect 226576 126216 226582 126268
rect 227622 126216 227628 126268
rect 227680 126256 227686 126268
rect 241974 126256 241980 126268
rect 227680 126228 241980 126256
rect 227680 126216 227686 126228
rect 241974 126216 241980 126228
rect 242032 126216 242038 126268
rect 244918 126216 244924 126268
rect 244976 126256 244982 126268
rect 255590 126256 255596 126268
rect 244976 126228 255596 126256
rect 244976 126216 244982 126228
rect 255590 126216 255596 126228
rect 255648 126216 255654 126268
rect 266998 126216 267004 126268
rect 267056 126256 267062 126268
rect 271874 126256 271880 126268
rect 267056 126228 271880 126256
rect 267056 126216 267062 126228
rect 271874 126216 271880 126228
rect 271932 126216 271938 126268
rect 273990 126216 273996 126268
rect 274048 126256 274054 126268
rect 277302 126256 277308 126268
rect 274048 126228 277308 126256
rect 274048 126216 274054 126228
rect 277302 126216 277308 126228
rect 277360 126216 277366 126268
rect 303706 126216 303712 126268
rect 303764 126256 303770 126268
rect 306374 126256 306380 126268
rect 303764 126228 306380 126256
rect 303764 126216 303770 126228
rect 306374 126216 306380 126228
rect 306432 126216 306438 126268
rect 315482 126216 315488 126268
rect 315540 126256 315546 126268
rect 318058 126256 318064 126268
rect 315540 126228 318064 126256
rect 315540 126216 315546 126228
rect 318058 126216 318064 126228
rect 318116 126216 318122 126268
rect 357250 126216 357256 126268
rect 357308 126256 357314 126268
rect 375374 126256 375380 126268
rect 357308 126228 375380 126256
rect 357308 126216 357314 126228
rect 375374 126216 375380 126228
rect 375432 126216 375438 126268
rect 379882 126216 379888 126268
rect 379940 126256 379946 126268
rect 400858 126256 400864 126268
rect 379940 126228 400864 126256
rect 379940 126216 379946 126228
rect 400858 126216 400864 126228
rect 400916 126216 400922 126268
rect 404446 126216 404452 126268
rect 404504 126256 404510 126268
rect 436738 126256 436744 126268
rect 404504 126228 436744 126256
rect 404504 126216 404510 126228
rect 436738 126216 436744 126228
rect 436796 126216 436802 126268
rect 442534 126216 442540 126268
rect 442592 126256 442598 126268
rect 482278 126256 482284 126268
rect 442592 126228 482284 126256
rect 442592 126216 442598 126228
rect 482278 126216 482284 126228
rect 482336 126216 482342 126268
rect 492398 126216 492404 126268
rect 492456 126256 492462 126268
rect 495989 126259 496047 126265
rect 495989 126256 496001 126259
rect 492456 126228 496001 126256
rect 492456 126216 492462 126228
rect 495989 126225 496001 126228
rect 496035 126225 496047 126259
rect 495989 126219 496047 126225
rect 512733 126259 512791 126265
rect 512733 126225 512745 126259
rect 512779 126256 512791 126259
rect 568574 126256 568580 126268
rect 512779 126228 568580 126256
rect 512779 126225 512791 126228
rect 512733 126219 512791 126225
rect 568574 126216 568580 126228
rect 568632 126216 568638 126268
rect 63402 126148 63408 126200
rect 63460 126188 63466 126200
rect 116762 126188 116768 126200
rect 63460 126160 116768 126188
rect 63460 126148 63466 126160
rect 116762 126148 116768 126160
rect 116820 126148 116826 126200
rect 144178 126148 144184 126200
rect 144236 126188 144242 126200
rect 168466 126188 168472 126200
rect 144236 126160 168472 126188
rect 144236 126148 144242 126160
rect 168466 126148 168472 126160
rect 168524 126148 168530 126200
rect 169662 126148 169668 126200
rect 169720 126188 169726 126200
rect 169720 126160 173112 126188
rect 169720 126148 169726 126160
rect 70210 126080 70216 126132
rect 70268 126120 70274 126132
rect 122190 126120 122196 126132
rect 70268 126092 122196 126120
rect 70268 126080 70274 126092
rect 122190 126080 122196 126092
rect 122248 126080 122254 126132
rect 148318 126080 148324 126132
rect 148376 126120 148382 126132
rect 148376 126092 161612 126120
rect 148376 126080 148382 126092
rect 68278 126012 68284 126064
rect 68336 126052 68342 126064
rect 114094 126052 114100 126064
rect 68336 126024 114100 126052
rect 68336 126012 68342 126024
rect 114094 126012 114100 126024
rect 114152 126012 114158 126064
rect 151078 126012 151084 126064
rect 151136 126052 151142 126064
rect 151136 126024 161474 126052
rect 151136 126012 151142 126024
rect 58618 125944 58624 125996
rect 58676 125984 58682 125996
rect 102226 125984 102232 125996
rect 58676 125956 102232 125984
rect 58676 125944 58682 125956
rect 102226 125944 102232 125956
rect 102284 125944 102290 125996
rect 50338 125876 50344 125928
rect 50396 125916 50402 125928
rect 91186 125916 91192 125928
rect 50396 125888 91192 125916
rect 50396 125876 50402 125888
rect 91186 125876 91192 125888
rect 91244 125876 91250 125928
rect 161446 125916 161474 126024
rect 161584 125984 161612 126092
rect 164878 126080 164884 126132
rect 164936 126120 164942 126132
rect 171226 126120 171232 126132
rect 164936 126092 171232 126120
rect 164936 126080 164942 126092
rect 171226 126080 171232 126092
rect 171284 126080 171290 126132
rect 173084 126052 173112 126160
rect 173802 126148 173808 126200
rect 173860 126188 173866 126200
rect 201126 126188 201132 126200
rect 173860 126160 201132 126188
rect 173860 126148 173866 126160
rect 201126 126148 201132 126160
rect 201184 126148 201190 126200
rect 202782 126148 202788 126200
rect 202840 126188 202846 126200
rect 222930 126188 222936 126200
rect 202840 126160 222936 126188
rect 202840 126148 202846 126160
rect 222930 126148 222936 126160
rect 222988 126148 222994 126200
rect 226978 126148 226984 126200
rect 227036 126188 227042 126200
rect 241054 126188 241060 126200
rect 227036 126160 241060 126188
rect 227036 126148 227042 126160
rect 241054 126148 241060 126160
rect 241112 126148 241118 126200
rect 251818 126148 251824 126200
rect 251876 126188 251882 126200
rect 260098 126188 260104 126200
rect 251876 126160 260104 126188
rect 251876 126148 251882 126160
rect 260098 126148 260104 126160
rect 260156 126148 260162 126200
rect 456150 126148 456156 126200
rect 456208 126188 456214 126200
rect 476758 126188 476764 126200
rect 456208 126160 476764 126188
rect 456208 126148 456214 126160
rect 476758 126148 476764 126160
rect 476816 126148 476822 126200
rect 483382 126148 483388 126200
rect 483440 126188 483446 126200
rect 529198 126188 529204 126200
rect 483440 126160 529204 126188
rect 483440 126148 483446 126160
rect 529198 126148 529204 126160
rect 529256 126148 529262 126200
rect 173158 126080 173164 126132
rect 173216 126120 173222 126132
rect 186590 126120 186596 126132
rect 173216 126092 186596 126120
rect 173216 126080 173222 126092
rect 186590 126080 186596 126092
rect 186648 126080 186654 126132
rect 186958 126080 186964 126132
rect 187016 126120 187022 126132
rect 210234 126120 210240 126132
rect 187016 126092 210240 126120
rect 187016 126080 187022 126092
rect 210234 126080 210240 126092
rect 210292 126080 210298 126132
rect 211062 126080 211068 126132
rect 211120 126120 211126 126132
rect 230198 126120 230204 126132
rect 211120 126092 230204 126120
rect 211120 126080 211126 126092
rect 230198 126080 230204 126092
rect 230256 126080 230262 126132
rect 231762 126080 231768 126132
rect 231820 126120 231826 126132
rect 245470 126120 245476 126132
rect 231820 126092 245476 126120
rect 231820 126080 231826 126092
rect 245470 126080 245476 126092
rect 245528 126080 245534 126132
rect 277302 126080 277308 126132
rect 277360 126120 277366 126132
rect 280062 126120 280068 126132
rect 277360 126092 280068 126120
rect 277360 126080 277366 126092
rect 280062 126080 280068 126092
rect 280120 126080 280126 126132
rect 465721 126123 465779 126129
rect 465721 126089 465733 126123
rect 465767 126120 465779 126123
rect 472618 126120 472624 126132
rect 465767 126092 472624 126120
rect 465767 126089 465779 126092
rect 465721 126083 465779 126089
rect 472618 126080 472624 126092
rect 472676 126080 472682 126132
rect 477862 126080 477868 126132
rect 477920 126120 477926 126132
rect 522298 126120 522304 126132
rect 477920 126092 522304 126120
rect 477920 126080 477926 126092
rect 522298 126080 522304 126092
rect 522356 126080 522362 126132
rect 176013 126055 176071 126061
rect 176013 126052 176025 126055
rect 173084 126024 176025 126052
rect 176013 126021 176025 126024
rect 176059 126021 176071 126055
rect 176013 126015 176071 126021
rect 180058 126012 180064 126064
rect 180116 126052 180122 126064
rect 196618 126052 196624 126064
rect 180116 126024 196624 126052
rect 180116 126012 180122 126024
rect 196618 126012 196624 126024
rect 196676 126012 196682 126064
rect 198642 126012 198648 126064
rect 198700 126052 198706 126064
rect 220170 126052 220176 126064
rect 198700 126024 220176 126052
rect 198700 126012 198706 126024
rect 220170 126012 220176 126024
rect 220228 126012 220234 126064
rect 222102 126012 222108 126064
rect 222160 126052 222166 126064
rect 238294 126052 238300 126064
rect 222160 126024 238300 126052
rect 222160 126012 222166 126024
rect 238294 126012 238300 126024
rect 238352 126012 238358 126064
rect 462498 126012 462504 126064
rect 462556 126052 462562 126064
rect 504358 126052 504364 126064
rect 462556 126024 504364 126052
rect 462556 126012 462562 126024
rect 504358 126012 504364 126024
rect 504416 126012 504422 126064
rect 510522 126012 510528 126064
rect 510580 126052 510586 126064
rect 533430 126052 533436 126064
rect 510580 126024 533436 126052
rect 510580 126012 510586 126024
rect 533430 126012 533436 126024
rect 533488 126012 533494 126064
rect 172974 125984 172980 125996
rect 161584 125956 172980 125984
rect 172974 125944 172980 125956
rect 173032 125944 173038 125996
rect 181438 125944 181444 125996
rect 181496 125984 181502 125996
rect 202046 125984 202052 125996
rect 181496 125956 202052 125984
rect 181496 125944 181502 125956
rect 202046 125944 202052 125956
rect 202104 125944 202110 125996
rect 204162 125944 204168 125996
rect 204220 125984 204226 125996
rect 224678 125984 224684 125996
rect 204220 125956 224684 125984
rect 204220 125944 204226 125956
rect 224678 125944 224684 125956
rect 224736 125944 224742 125996
rect 233142 125944 233148 125996
rect 233200 125984 233206 125996
rect 246482 125984 246488 125996
rect 233200 125956 246488 125984
rect 233200 125944 233206 125956
rect 246482 125944 246488 125956
rect 246540 125944 246546 125996
rect 260098 125944 260104 125996
rect 260156 125984 260162 125996
rect 262858 125984 262864 125996
rect 260156 125956 262864 125984
rect 260156 125944 260162 125956
rect 262858 125944 262864 125956
rect 262916 125944 262922 125996
rect 451550 125944 451556 125996
rect 451608 125984 451614 125996
rect 483658 125984 483664 125996
rect 451608 125956 483664 125984
rect 451608 125944 451614 125956
rect 483658 125944 483664 125956
rect 483716 125944 483722 125996
rect 486050 125944 486056 125996
rect 486108 125984 486114 125996
rect 526438 125984 526444 125996
rect 486108 125956 526444 125984
rect 486108 125944 486114 125956
rect 526438 125944 526444 125956
rect 526496 125944 526502 125996
rect 167546 125916 167552 125928
rect 161446 125888 167552 125916
rect 167546 125876 167552 125888
rect 167604 125876 167610 125928
rect 184198 125876 184204 125928
rect 184256 125916 184262 125928
rect 204806 125916 204812 125928
rect 184256 125888 204812 125916
rect 184256 125876 184262 125888
rect 204806 125876 204812 125888
rect 204864 125876 204870 125928
rect 208302 125876 208308 125928
rect 208360 125916 208366 125928
rect 227438 125916 227444 125928
rect 208360 125888 227444 125916
rect 208360 125876 208366 125888
rect 227438 125876 227444 125888
rect 227496 125876 227502 125928
rect 491478 125876 491484 125928
rect 491536 125916 491542 125928
rect 507854 125916 507860 125928
rect 491536 125888 507860 125916
rect 491536 125876 491542 125888
rect 507854 125876 507860 125888
rect 507912 125876 507918 125928
rect 514021 125919 514079 125925
rect 514021 125885 514033 125919
rect 514067 125916 514079 125919
rect 520918 125916 520924 125928
rect 514067 125888 520924 125916
rect 514067 125885 514079 125888
rect 514021 125879 514079 125885
rect 520918 125876 520924 125888
rect 520976 125876 520982 125928
rect 53098 125808 53104 125860
rect 53156 125848 53162 125860
rect 77754 125848 77760 125860
rect 53156 125820 77760 125848
rect 53156 125808 53162 125820
rect 77754 125808 77760 125820
rect 77812 125808 77818 125860
rect 178678 125808 178684 125860
rect 178736 125848 178742 125860
rect 192018 125848 192024 125860
rect 178736 125820 192024 125848
rect 178736 125808 178742 125820
rect 192018 125808 192024 125820
rect 192076 125808 192082 125860
rect 205542 125808 205548 125860
rect 205600 125848 205606 125860
rect 214561 125851 214619 125857
rect 214561 125848 214573 125851
rect 205600 125820 214573 125848
rect 205600 125808 205606 125820
rect 214561 125817 214573 125820
rect 214607 125817 214619 125851
rect 214561 125811 214619 125817
rect 215202 125808 215208 125860
rect 215260 125848 215266 125860
rect 232866 125848 232872 125860
rect 215260 125820 232872 125848
rect 215260 125808 215266 125820
rect 232866 125808 232872 125820
rect 232924 125808 232930 125860
rect 262858 125808 262864 125860
rect 262916 125848 262922 125860
rect 269206 125848 269212 125860
rect 262916 125820 269212 125848
rect 262916 125808 262922 125820
rect 269206 125808 269212 125820
rect 269264 125808 269270 125860
rect 270402 125808 270408 125860
rect 270460 125848 270466 125860
rect 275554 125848 275560 125860
rect 270460 125820 275560 125848
rect 270460 125808 270466 125820
rect 275554 125808 275560 125820
rect 275612 125808 275618 125860
rect 505002 125808 505008 125860
rect 505060 125848 505066 125860
rect 512733 125851 512791 125857
rect 512733 125848 512745 125851
rect 505060 125820 512745 125848
rect 505060 125808 505066 125820
rect 512733 125817 512745 125820
rect 512779 125817 512791 125851
rect 512733 125811 512791 125817
rect 213178 125740 213184 125792
rect 213236 125780 213242 125792
rect 229278 125780 229284 125792
rect 213236 125752 229284 125780
rect 213236 125740 213242 125752
rect 229278 125740 229284 125752
rect 229336 125740 229342 125792
rect 259362 125740 259368 125792
rect 259420 125780 259426 125792
rect 266446 125780 266452 125792
rect 259420 125752 266452 125780
rect 259420 125740 259426 125752
rect 266446 125740 266452 125752
rect 266504 125740 266510 125792
rect 269022 125740 269028 125792
rect 269080 125780 269086 125792
rect 273714 125780 273720 125792
rect 269080 125752 273720 125780
rect 269080 125740 269086 125752
rect 273714 125740 273720 125752
rect 273772 125740 273778 125792
rect 309042 125740 309048 125792
rect 309100 125780 309106 125792
rect 313274 125780 313280 125792
rect 309100 125752 313280 125780
rect 309100 125740 309106 125752
rect 313274 125740 313280 125752
rect 313332 125740 313338 125792
rect 219342 125672 219348 125724
rect 219400 125712 219406 125724
rect 235626 125712 235632 125724
rect 219400 125684 235632 125712
rect 219400 125672 219406 125684
rect 235626 125672 235632 125684
rect 235684 125672 235690 125724
rect 264238 125672 264244 125724
rect 264296 125712 264302 125724
rect 267366 125712 267372 125724
rect 264296 125684 267372 125712
rect 264296 125672 264302 125684
rect 267366 125672 267372 125684
rect 267424 125672 267430 125724
rect 271782 125672 271788 125724
rect 271840 125712 271846 125724
rect 276382 125712 276388 125724
rect 271840 125684 276388 125712
rect 271840 125672 271846 125684
rect 276382 125672 276388 125684
rect 276440 125672 276446 125724
rect 280798 125672 280804 125724
rect 280856 125712 280862 125724
rect 282730 125712 282736 125724
rect 280856 125684 282736 125712
rect 280856 125672 280862 125684
rect 282730 125672 282736 125684
rect 282788 125672 282794 125724
rect 282822 125672 282828 125724
rect 282880 125712 282886 125724
rect 284386 125712 284392 125724
rect 282880 125684 284392 125712
rect 282880 125672 282886 125684
rect 284386 125672 284392 125684
rect 284444 125672 284450 125724
rect 301958 125672 301964 125724
rect 302016 125712 302022 125724
rect 303614 125712 303620 125724
rect 302016 125684 303620 125712
rect 302016 125672 302022 125684
rect 303614 125672 303620 125684
rect 303672 125672 303678 125724
rect 308306 125672 308312 125724
rect 308364 125712 308370 125724
rect 311894 125712 311900 125724
rect 308364 125684 311900 125712
rect 308364 125672 308370 125684
rect 311894 125672 311900 125684
rect 311952 125672 311958 125724
rect 319162 125672 319168 125724
rect 319220 125712 319226 125724
rect 322198 125712 322204 125724
rect 319220 125684 322204 125712
rect 319220 125672 319226 125684
rect 322198 125672 322204 125684
rect 322256 125672 322262 125724
rect 326430 125672 326436 125724
rect 326488 125712 326494 125724
rect 331766 125712 331772 125724
rect 326488 125684 331772 125712
rect 326488 125672 326494 125684
rect 331766 125672 331772 125684
rect 331824 125672 331830 125724
rect 333698 125672 333704 125724
rect 333756 125712 333762 125724
rect 334618 125712 334624 125724
rect 333756 125684 334624 125712
rect 333756 125672 333762 125684
rect 334618 125672 334624 125684
rect 334676 125672 334682 125724
rect 337286 125672 337292 125724
rect 337344 125712 337350 125724
rect 340138 125712 340144 125724
rect 337344 125684 340144 125712
rect 337344 125672 337350 125684
rect 340138 125672 340144 125684
rect 340196 125672 340202 125724
rect 348142 125672 348148 125724
rect 348200 125712 348206 125724
rect 353938 125712 353944 125724
rect 348200 125684 353944 125712
rect 348200 125672 348206 125684
rect 353938 125672 353944 125684
rect 353996 125672 354002 125724
rect 356330 125672 356336 125724
rect 356388 125712 356394 125724
rect 357342 125712 357348 125724
rect 356388 125684 357348 125712
rect 356388 125672 356394 125684
rect 357342 125672 357348 125684
rect 357400 125672 357406 125724
rect 369026 125672 369032 125724
rect 369084 125712 369090 125724
rect 371878 125712 371884 125724
rect 369084 125684 371884 125712
rect 369084 125672 369090 125684
rect 371878 125672 371884 125684
rect 371936 125672 371942 125724
rect 445202 125672 445208 125724
rect 445260 125712 445266 125724
rect 447778 125712 447784 125724
rect 445260 125684 447784 125712
rect 445260 125672 445266 125684
rect 447778 125672 447784 125684
rect 447836 125672 447842 125724
rect 72418 125604 72424 125656
rect 72476 125644 72482 125656
rect 74166 125644 74172 125656
rect 72476 125616 74172 125644
rect 72476 125604 72482 125616
rect 74166 125604 74172 125616
rect 74224 125604 74230 125656
rect 118602 125644 118608 125656
rect 115906 125616 118608 125644
rect 39298 125468 39304 125520
rect 39356 125508 39362 125520
rect 75086 125508 75092 125520
rect 39356 125480 75092 125508
rect 39356 125468 39362 125480
rect 75086 125468 75092 125480
rect 75144 125468 75150 125520
rect 32398 125400 32404 125452
rect 32456 125440 32462 125452
rect 81434 125440 81440 125452
rect 32456 125412 81440 125440
rect 32456 125400 32462 125412
rect 81434 125400 81440 125412
rect 81492 125400 81498 125452
rect 66162 125332 66168 125384
rect 66220 125372 66226 125384
rect 115906 125372 115934 125616
rect 118602 125604 118608 125616
rect 118660 125604 118666 125656
rect 128998 125604 129004 125656
rect 129056 125644 129062 125656
rect 132218 125644 132224 125656
rect 129056 125616 132224 125644
rect 129056 125604 129062 125616
rect 132218 125604 132224 125616
rect 132276 125604 132282 125656
rect 133138 125604 133144 125656
rect 133196 125644 133202 125656
rect 137646 125644 137652 125656
rect 133196 125616 137652 125644
rect 133196 125604 133202 125616
rect 137646 125604 137652 125616
rect 137704 125604 137710 125656
rect 183646 125604 183652 125656
rect 183704 125644 183710 125656
rect 184842 125644 184848 125656
rect 183704 125616 184848 125644
rect 183704 125604 183710 125616
rect 184842 125604 184848 125616
rect 184900 125604 184906 125656
rect 206278 125604 206284 125656
rect 206336 125644 206342 125656
rect 207474 125644 207480 125656
rect 206336 125616 207480 125644
rect 206336 125604 206342 125616
rect 207474 125604 207480 125616
rect 207532 125604 207538 125656
rect 242158 125604 242164 125656
rect 242216 125644 242222 125656
rect 248322 125644 248328 125656
rect 242216 125616 248328 125644
rect 242216 125604 242222 125616
rect 248322 125604 248328 125616
rect 248380 125604 248386 125656
rect 249150 125604 249156 125656
rect 249208 125644 249214 125656
rect 254670 125644 254676 125656
rect 249208 125616 254676 125644
rect 249208 125604 249214 125616
rect 254670 125604 254676 125616
rect 254728 125604 254734 125656
rect 262950 125604 262956 125656
rect 263008 125644 263014 125656
rect 265526 125644 265532 125656
rect 263008 125616 265532 125644
rect 263008 125604 263014 125616
rect 265526 125604 265532 125616
rect 265584 125604 265590 125656
rect 268378 125604 268384 125656
rect 268436 125644 268442 125656
rect 270954 125644 270960 125656
rect 268436 125616 270960 125644
rect 268436 125604 268442 125616
rect 270954 125604 270960 125616
rect 271012 125604 271018 125656
rect 273898 125604 273904 125656
rect 273956 125644 273962 125656
rect 274634 125644 274640 125656
rect 273956 125616 274640 125644
rect 273956 125604 273962 125616
rect 274634 125604 274640 125616
rect 274692 125604 274698 125656
rect 278682 125604 278688 125656
rect 278740 125644 278746 125656
rect 281902 125644 281908 125656
rect 278740 125616 281908 125644
rect 278740 125604 278746 125616
rect 281902 125604 281908 125616
rect 281960 125604 281966 125656
rect 282178 125604 282184 125656
rect 282236 125644 282242 125656
rect 283650 125644 283656 125656
rect 282236 125616 283656 125644
rect 282236 125604 282242 125616
rect 283650 125604 283656 125616
rect 283708 125604 283714 125656
rect 288342 125604 288348 125656
rect 288400 125644 288406 125656
rect 289078 125644 289084 125656
rect 288400 125616 289084 125644
rect 288400 125604 288406 125616
rect 289078 125604 289084 125616
rect 289136 125604 289142 125656
rect 289906 125604 289912 125656
rect 289964 125644 289970 125656
rect 290918 125644 290924 125656
rect 289964 125616 290924 125644
rect 289964 125604 289970 125616
rect 290918 125604 290924 125616
rect 290976 125604 290982 125656
rect 292574 125604 292580 125656
rect 292632 125644 292638 125656
rect 293678 125644 293684 125656
rect 292632 125616 293684 125644
rect 292632 125604 292638 125616
rect 293678 125604 293684 125616
rect 293736 125604 293742 125656
rect 297358 125604 297364 125656
rect 297416 125644 297422 125656
rect 298094 125644 298100 125656
rect 297416 125616 298100 125644
rect 297416 125604 297422 125616
rect 298094 125604 298100 125616
rect 298152 125604 298158 125656
rect 298278 125604 298284 125656
rect 298336 125644 298342 125656
rect 299290 125644 299296 125656
rect 298336 125616 299296 125644
rect 298336 125604 298342 125616
rect 299290 125604 299296 125616
rect 299348 125604 299354 125656
rect 300118 125604 300124 125656
rect 300176 125644 300182 125656
rect 300762 125644 300768 125656
rect 300176 125616 300768 125644
rect 300176 125604 300182 125616
rect 300762 125604 300768 125616
rect 300820 125604 300826 125656
rect 301038 125604 301044 125656
rect 301096 125644 301102 125656
rect 302234 125644 302240 125656
rect 301096 125616 302240 125644
rect 301096 125604 301102 125616
rect 302234 125604 302240 125616
rect 302292 125604 302298 125656
rect 302786 125604 302792 125656
rect 302844 125644 302850 125656
rect 304994 125644 305000 125656
rect 302844 125616 305000 125644
rect 302844 125604 302850 125616
rect 304994 125604 305000 125616
rect 305052 125604 305058 125656
rect 305546 125604 305552 125656
rect 305604 125644 305610 125656
rect 306282 125644 306288 125656
rect 305604 125616 306288 125644
rect 305604 125604 305610 125616
rect 306282 125604 306288 125616
rect 306340 125604 306346 125656
rect 306466 125604 306472 125656
rect 306524 125644 306530 125656
rect 309134 125644 309140 125656
rect 306524 125616 309140 125644
rect 306524 125604 306530 125616
rect 309134 125604 309140 125616
rect 309192 125604 309198 125656
rect 310974 125604 310980 125656
rect 311032 125644 311038 125656
rect 311710 125644 311716 125656
rect 311032 125616 311716 125644
rect 311032 125604 311038 125616
rect 311710 125604 311716 125616
rect 311768 125604 311774 125656
rect 313734 125604 313740 125656
rect 313792 125644 313798 125656
rect 314470 125644 314476 125656
rect 313792 125616 314476 125644
rect 313792 125604 313798 125616
rect 314470 125604 314476 125616
rect 314528 125604 314534 125656
rect 316402 125604 316408 125656
rect 316460 125644 316466 125656
rect 317230 125644 317236 125656
rect 316460 125616 317236 125644
rect 316460 125604 316466 125616
rect 317230 125604 317236 125616
rect 317288 125604 317294 125656
rect 318242 125604 318248 125656
rect 318300 125644 318306 125656
rect 318702 125644 318708 125656
rect 318300 125616 318708 125644
rect 318300 125604 318306 125616
rect 318702 125604 318708 125616
rect 318760 125604 318766 125656
rect 320082 125604 320088 125656
rect 320140 125644 320146 125656
rect 320818 125644 320824 125656
rect 320140 125616 320824 125644
rect 320140 125604 320146 125616
rect 320818 125604 320824 125616
rect 320876 125604 320882 125656
rect 321002 125604 321008 125656
rect 321060 125644 321066 125656
rect 321462 125644 321468 125656
rect 321060 125616 321468 125644
rect 321060 125604 321066 125616
rect 321462 125604 321468 125616
rect 321520 125604 321526 125656
rect 321830 125604 321836 125656
rect 321888 125644 321894 125656
rect 322842 125644 322848 125656
rect 321888 125616 322848 125644
rect 321888 125604 321894 125616
rect 322842 125604 322848 125616
rect 322900 125604 322906 125656
rect 323670 125604 323676 125656
rect 323728 125644 323734 125656
rect 324222 125644 324228 125656
rect 323728 125616 324228 125644
rect 323728 125604 323734 125616
rect 324222 125604 324228 125616
rect 324280 125604 324286 125656
rect 324590 125604 324596 125656
rect 324648 125644 324654 125656
rect 325510 125644 325516 125656
rect 324648 125616 325516 125644
rect 324648 125604 324654 125616
rect 325510 125604 325516 125616
rect 325568 125604 325574 125656
rect 327350 125604 327356 125656
rect 327408 125644 327414 125656
rect 328362 125644 328368 125656
rect 327408 125616 328368 125644
rect 327408 125604 327414 125616
rect 328362 125604 328368 125616
rect 328420 125604 328426 125656
rect 329098 125604 329104 125656
rect 329156 125644 329162 125656
rect 329742 125644 329748 125656
rect 329156 125616 329748 125644
rect 329156 125604 329162 125616
rect 329742 125604 329748 125616
rect 329800 125604 329806 125656
rect 330018 125604 330024 125656
rect 330076 125644 330082 125656
rect 331122 125644 331128 125656
rect 330076 125616 331128 125644
rect 330076 125604 330082 125616
rect 331122 125604 331128 125616
rect 331180 125604 331186 125656
rect 331858 125604 331864 125656
rect 331916 125644 331922 125656
rect 332502 125644 332508 125656
rect 331916 125616 332508 125644
rect 331916 125604 331922 125616
rect 332502 125604 332508 125616
rect 332560 125604 332566 125656
rect 334526 125604 334532 125656
rect 334584 125644 334590 125656
rect 335262 125644 335268 125656
rect 334584 125616 335268 125644
rect 334584 125604 334590 125616
rect 335262 125604 335268 125616
rect 335320 125604 335326 125656
rect 335446 125604 335452 125656
rect 335504 125644 335510 125656
rect 336550 125644 336556 125656
rect 335504 125616 336556 125644
rect 335504 125604 335510 125616
rect 336550 125604 336556 125616
rect 336608 125604 336614 125656
rect 338206 125604 338212 125656
rect 338264 125644 338270 125656
rect 339310 125644 339316 125656
rect 338264 125616 339316 125644
rect 338264 125604 338270 125616
rect 339310 125604 339316 125616
rect 339368 125604 339374 125656
rect 340046 125604 340052 125656
rect 340104 125644 340110 125656
rect 340782 125644 340788 125656
rect 340104 125616 340788 125644
rect 340104 125604 340110 125616
rect 340782 125604 340788 125616
rect 340840 125604 340846 125656
rect 340966 125604 340972 125656
rect 341024 125644 341030 125656
rect 342070 125644 342076 125656
rect 341024 125616 342076 125644
rect 341024 125604 341030 125616
rect 342070 125604 342076 125616
rect 342128 125604 342134 125656
rect 342714 125604 342720 125656
rect 342772 125644 342778 125656
rect 343542 125644 343548 125656
rect 342772 125616 343548 125644
rect 342772 125604 342778 125616
rect 343542 125604 343548 125616
rect 343600 125604 343606 125656
rect 345474 125604 345480 125656
rect 345532 125644 345538 125656
rect 346302 125644 346308 125656
rect 345532 125616 346308 125644
rect 345532 125604 345538 125616
rect 346302 125604 346308 125616
rect 346360 125604 346366 125656
rect 349982 125604 349988 125656
rect 350040 125644 350046 125656
rect 350442 125644 350448 125656
rect 350040 125616 350448 125644
rect 350040 125604 350046 125616
rect 350442 125604 350448 125616
rect 350500 125604 350506 125656
rect 352742 125604 352748 125656
rect 352800 125644 352806 125656
rect 353202 125644 353208 125656
rect 352800 125616 353208 125644
rect 352800 125604 352806 125616
rect 353202 125604 353208 125616
rect 353260 125604 353266 125656
rect 353662 125604 353668 125656
rect 353720 125644 353726 125656
rect 354582 125644 354588 125656
rect 353720 125616 354588 125644
rect 353720 125604 353726 125616
rect 354582 125604 354588 125616
rect 354640 125604 354646 125656
rect 355410 125604 355416 125656
rect 355468 125644 355474 125656
rect 356698 125644 356704 125656
rect 355468 125616 356704 125644
rect 355468 125604 355474 125616
rect 356698 125604 356704 125616
rect 356756 125604 356762 125656
rect 358170 125604 358176 125656
rect 358228 125644 358234 125656
rect 358722 125644 358728 125656
rect 358228 125616 358728 125644
rect 358228 125604 358234 125616
rect 358722 125604 358728 125616
rect 358780 125604 358786 125656
rect 359090 125604 359096 125656
rect 359148 125644 359154 125656
rect 360102 125644 360108 125656
rect 359148 125616 360108 125644
rect 359148 125604 359154 125616
rect 360102 125604 360108 125616
rect 360160 125604 360166 125656
rect 360838 125604 360844 125656
rect 360896 125644 360902 125656
rect 361482 125644 361488 125656
rect 360896 125616 361488 125644
rect 360896 125604 360902 125616
rect 361482 125604 361488 125616
rect 361540 125604 361546 125656
rect 361758 125604 361764 125656
rect 361816 125644 361822 125656
rect 362862 125644 362868 125656
rect 361816 125616 362868 125644
rect 361816 125604 361822 125616
rect 362862 125604 362868 125616
rect 362920 125604 362926 125656
rect 363598 125604 363604 125656
rect 363656 125644 363662 125656
rect 364242 125644 364248 125656
rect 363656 125616 364248 125644
rect 363656 125604 363662 125616
rect 364242 125604 364248 125616
rect 364300 125604 364306 125656
rect 364518 125604 364524 125656
rect 364576 125644 364582 125656
rect 365622 125644 365628 125656
rect 364576 125616 365628 125644
rect 364576 125604 364582 125616
rect 365622 125604 365628 125616
rect 365680 125604 365686 125656
rect 366358 125604 366364 125656
rect 366416 125644 366422 125656
rect 367002 125644 367008 125656
rect 366416 125616 367008 125644
rect 366416 125604 366422 125616
rect 367002 125604 367008 125616
rect 367060 125604 367066 125656
rect 367186 125604 367192 125656
rect 367244 125644 367250 125656
rect 368382 125644 368388 125656
rect 367244 125616 368388 125644
rect 367244 125604 367250 125616
rect 368382 125604 368388 125616
rect 368440 125604 368446 125656
rect 369946 125604 369952 125656
rect 370004 125644 370010 125656
rect 371142 125644 371148 125656
rect 370004 125616 371148 125644
rect 370004 125604 370010 125616
rect 371142 125604 371148 125616
rect 371200 125604 371206 125656
rect 371786 125604 371792 125656
rect 371844 125644 371850 125656
rect 372522 125644 372528 125656
rect 371844 125616 372528 125644
rect 371844 125604 371850 125616
rect 372522 125604 372528 125616
rect 372580 125604 372586 125656
rect 372706 125604 372712 125656
rect 372764 125644 372770 125656
rect 373902 125644 373908 125656
rect 372764 125616 373908 125644
rect 372764 125604 372770 125616
rect 373902 125604 373908 125616
rect 373960 125604 373966 125656
rect 374454 125604 374460 125656
rect 374512 125644 374518 125656
rect 375190 125644 375196 125656
rect 374512 125616 375196 125644
rect 374512 125604 374518 125616
rect 375190 125604 375196 125616
rect 375248 125604 375254 125656
rect 381722 125604 381728 125656
rect 381780 125644 381786 125656
rect 382182 125644 382188 125656
rect 381780 125616 382188 125644
rect 381780 125604 381786 125616
rect 382182 125604 382188 125616
rect 382240 125604 382246 125656
rect 382642 125604 382648 125656
rect 382700 125644 382706 125656
rect 383470 125644 383476 125656
rect 382700 125616 383476 125644
rect 382700 125604 382706 125616
rect 383470 125604 383476 125616
rect 383528 125604 383534 125656
rect 384482 125604 384488 125656
rect 384540 125644 384546 125656
rect 384942 125644 384948 125656
rect 384540 125616 384948 125644
rect 384540 125604 384546 125616
rect 384942 125604 384948 125616
rect 385000 125604 385006 125656
rect 385402 125604 385408 125656
rect 385460 125644 385466 125656
rect 386230 125644 386236 125656
rect 385460 125616 386236 125644
rect 385460 125604 385466 125616
rect 386230 125604 386236 125616
rect 386288 125604 386294 125656
rect 387150 125604 387156 125656
rect 387208 125644 387214 125656
rect 387702 125644 387708 125656
rect 387208 125616 387708 125644
rect 387208 125604 387214 125616
rect 387702 125604 387708 125616
rect 387760 125604 387766 125656
rect 389910 125604 389916 125656
rect 389968 125644 389974 125656
rect 390462 125644 390468 125656
rect 389968 125616 390468 125644
rect 389968 125604 389974 125616
rect 390462 125604 390468 125616
rect 390520 125604 390526 125656
rect 390830 125604 390836 125656
rect 390888 125644 390894 125656
rect 392578 125644 392584 125656
rect 390888 125616 392584 125644
rect 390888 125604 390894 125616
rect 392578 125604 392584 125616
rect 392636 125604 392642 125656
rect 392670 125604 392676 125656
rect 392728 125644 392734 125656
rect 393222 125644 393228 125656
rect 392728 125616 393228 125644
rect 392728 125604 392734 125616
rect 393222 125604 393228 125616
rect 393280 125604 393286 125656
rect 395338 125604 395344 125656
rect 395396 125644 395402 125656
rect 395982 125644 395988 125656
rect 395396 125616 395988 125644
rect 395396 125604 395402 125616
rect 395982 125604 395988 125616
rect 396040 125604 396046 125656
rect 396258 125604 396264 125656
rect 396316 125644 396322 125656
rect 397270 125644 397276 125656
rect 396316 125616 397276 125644
rect 396316 125604 396322 125616
rect 397270 125604 397276 125616
rect 397328 125604 397334 125656
rect 398098 125604 398104 125656
rect 398156 125644 398162 125656
rect 398742 125644 398748 125656
rect 398156 125616 398748 125644
rect 398156 125604 398162 125616
rect 398742 125604 398748 125616
rect 398800 125604 398806 125656
rect 400766 125604 400772 125656
rect 400824 125644 400830 125656
rect 401502 125644 401508 125656
rect 400824 125616 401508 125644
rect 400824 125604 400830 125616
rect 401502 125604 401508 125616
rect 401560 125604 401566 125656
rect 403526 125604 403532 125656
rect 403584 125644 403590 125656
rect 404262 125644 404268 125656
rect 403584 125616 404268 125644
rect 403584 125604 403590 125616
rect 404262 125604 404268 125616
rect 404320 125604 404326 125656
rect 406194 125604 406200 125656
rect 406252 125644 406258 125656
rect 407022 125644 407028 125656
rect 406252 125616 407028 125644
rect 406252 125604 406258 125616
rect 407022 125604 407028 125616
rect 407080 125604 407086 125656
rect 408954 125604 408960 125656
rect 409012 125644 409018 125656
rect 409782 125644 409788 125656
rect 409012 125616 409788 125644
rect 409012 125604 409018 125616
rect 409782 125604 409788 125616
rect 409840 125604 409846 125656
rect 411714 125604 411720 125656
rect 411772 125644 411778 125656
rect 412542 125644 412548 125656
rect 411772 125616 412548 125644
rect 411772 125604 411778 125616
rect 412542 125604 412548 125616
rect 412600 125604 412606 125656
rect 413462 125604 413468 125656
rect 413520 125644 413526 125656
rect 413922 125644 413928 125656
rect 413520 125616 413928 125644
rect 413520 125604 413526 125616
rect 413922 125604 413928 125616
rect 413980 125604 413986 125656
rect 414382 125604 414388 125656
rect 414440 125644 414446 125656
rect 415302 125644 415308 125656
rect 414440 125616 415308 125644
rect 414440 125604 414446 125616
rect 415302 125604 415308 125616
rect 415360 125604 415366 125656
rect 416222 125604 416228 125656
rect 416280 125644 416286 125656
rect 416682 125644 416688 125656
rect 416280 125616 416688 125644
rect 416280 125604 416286 125616
rect 416682 125604 416688 125616
rect 416740 125604 416746 125656
rect 417142 125604 417148 125656
rect 417200 125644 417206 125656
rect 418062 125644 418068 125656
rect 417200 125616 418068 125644
rect 417200 125604 417206 125616
rect 418062 125604 418068 125616
rect 418120 125604 418126 125656
rect 418890 125604 418896 125656
rect 418948 125644 418954 125656
rect 419442 125644 419448 125656
rect 418948 125616 419448 125644
rect 418948 125604 418954 125616
rect 419442 125604 419448 125616
rect 419500 125604 419506 125656
rect 421650 125604 421656 125656
rect 421708 125644 421714 125656
rect 422202 125644 422208 125656
rect 421708 125616 422208 125644
rect 421708 125604 421714 125616
rect 422202 125604 422208 125616
rect 422260 125604 422266 125656
rect 422570 125604 422576 125656
rect 422628 125644 422634 125656
rect 423582 125644 423588 125656
rect 422628 125616 423588 125644
rect 422628 125604 422634 125616
rect 423582 125604 423588 125616
rect 423640 125604 423646 125656
rect 424410 125604 424416 125656
rect 424468 125644 424474 125656
rect 424962 125644 424968 125656
rect 424468 125616 424968 125644
rect 424468 125604 424474 125616
rect 424962 125604 424968 125616
rect 425020 125604 425026 125656
rect 425238 125604 425244 125656
rect 425296 125644 425302 125656
rect 426342 125644 426348 125656
rect 425296 125616 426348 125644
rect 425296 125604 425302 125616
rect 426342 125604 426348 125616
rect 426400 125604 426406 125656
rect 427078 125604 427084 125656
rect 427136 125644 427142 125656
rect 427722 125644 427728 125656
rect 427136 125616 427728 125644
rect 427136 125604 427142 125616
rect 427722 125604 427728 125616
rect 427780 125604 427786 125656
rect 427998 125604 428004 125656
rect 428056 125644 428062 125656
rect 429102 125644 429108 125656
rect 428056 125616 429108 125644
rect 428056 125604 428062 125616
rect 429102 125604 429108 125616
rect 429160 125604 429166 125656
rect 429838 125604 429844 125656
rect 429896 125644 429902 125656
rect 430482 125644 430488 125656
rect 429896 125616 430488 125644
rect 429896 125604 429902 125616
rect 430482 125604 430488 125616
rect 430540 125604 430546 125656
rect 430758 125604 430764 125656
rect 430816 125644 430822 125656
rect 431862 125644 431868 125656
rect 430816 125616 431868 125644
rect 430816 125604 430822 125616
rect 431862 125604 431868 125616
rect 431920 125604 431926 125656
rect 432506 125604 432512 125656
rect 432564 125644 432570 125656
rect 433242 125644 433248 125656
rect 432564 125616 433248 125644
rect 432564 125604 432570 125616
rect 433242 125604 433248 125616
rect 433300 125604 433306 125656
rect 433426 125604 433432 125656
rect 433484 125644 433490 125656
rect 434622 125644 434628 125656
rect 433484 125616 434628 125644
rect 433484 125604 433490 125616
rect 434622 125604 434628 125616
rect 434680 125604 434686 125656
rect 435266 125604 435272 125656
rect 435324 125644 435330 125656
rect 436002 125644 436008 125656
rect 435324 125616 436008 125644
rect 435324 125604 435330 125616
rect 436002 125604 436008 125616
rect 436060 125604 436066 125656
rect 436186 125604 436192 125656
rect 436244 125644 436250 125656
rect 437382 125644 437388 125656
rect 436244 125616 437388 125644
rect 436244 125604 436250 125616
rect 437382 125604 437388 125616
rect 437440 125604 437446 125656
rect 438026 125604 438032 125656
rect 438084 125644 438090 125656
rect 439498 125644 439504 125656
rect 438084 125616 439504 125644
rect 438084 125604 438090 125616
rect 439498 125604 439504 125616
rect 439556 125604 439562 125656
rect 443454 125604 443460 125656
rect 443512 125644 443518 125656
rect 444190 125644 444196 125656
rect 443512 125616 444196 125644
rect 443512 125604 443518 125616
rect 444190 125604 444196 125616
rect 444248 125604 444254 125656
rect 446122 125604 446128 125656
rect 446180 125644 446186 125656
rect 446950 125644 446956 125656
rect 446180 125616 446956 125644
rect 446180 125604 446186 125616
rect 446950 125604 446956 125616
rect 447008 125604 447014 125656
rect 447962 125604 447968 125656
rect 448020 125644 448026 125656
rect 448422 125644 448428 125656
rect 448020 125616 448428 125644
rect 448020 125604 448026 125616
rect 448422 125604 448428 125616
rect 448480 125604 448486 125656
rect 450722 125604 450728 125656
rect 450780 125644 450786 125656
rect 451182 125644 451188 125656
rect 450780 125616 451188 125644
rect 450780 125604 450786 125616
rect 451182 125604 451188 125616
rect 451240 125604 451246 125656
rect 453390 125604 453396 125656
rect 453448 125644 453454 125656
rect 453942 125644 453948 125656
rect 453448 125616 453948 125644
rect 453448 125604 453454 125616
rect 453942 125604 453948 125616
rect 454000 125604 454006 125656
rect 454310 125604 454316 125656
rect 454368 125644 454374 125656
rect 455230 125644 455236 125656
rect 454368 125616 455236 125644
rect 454368 125604 454374 125616
rect 455230 125604 455236 125616
rect 455288 125604 455294 125656
rect 458818 125604 458824 125656
rect 458876 125644 458882 125656
rect 459462 125644 459468 125656
rect 458876 125616 459468 125644
rect 458876 125604 458882 125616
rect 459462 125604 459468 125616
rect 459520 125604 459526 125656
rect 461578 125604 461584 125656
rect 461636 125644 461642 125656
rect 462222 125644 462228 125656
rect 461636 125616 462228 125644
rect 461636 125604 461642 125616
rect 462222 125604 462228 125616
rect 462280 125604 462286 125656
rect 464246 125604 464252 125656
rect 464304 125644 464310 125656
rect 464982 125644 464988 125656
rect 464304 125616 464988 125644
rect 464304 125604 464310 125616
rect 464982 125604 464988 125616
rect 465040 125604 465046 125656
rect 465166 125604 465172 125656
rect 465224 125644 465230 125656
rect 466362 125644 466368 125656
rect 465224 125616 466368 125644
rect 465224 125604 465230 125616
rect 466362 125604 466368 125616
rect 466420 125604 466426 125656
rect 467006 125604 467012 125656
rect 467064 125644 467070 125656
rect 467742 125644 467748 125656
rect 467064 125616 467748 125644
rect 467064 125604 467070 125616
rect 467742 125604 467748 125616
rect 467800 125604 467806 125656
rect 467926 125604 467932 125656
rect 467984 125644 467990 125656
rect 469030 125644 469036 125656
rect 467984 125616 469036 125644
rect 467984 125604 467990 125616
rect 469030 125604 469036 125616
rect 469088 125604 469094 125656
rect 479702 125604 479708 125656
rect 479760 125644 479766 125656
rect 480162 125644 480168 125656
rect 479760 125616 480168 125644
rect 479760 125604 479766 125616
rect 480162 125604 480168 125616
rect 480220 125604 480226 125656
rect 480622 125604 480628 125656
rect 480680 125644 480686 125656
rect 480680 125616 485084 125644
rect 480680 125604 480686 125616
rect 66220 125344 115934 125372
rect 485056 125372 485084 125616
rect 485130 125604 485136 125656
rect 485188 125644 485194 125656
rect 485682 125644 485688 125656
rect 485188 125616 485688 125644
rect 485188 125604 485194 125616
rect 485682 125604 485688 125616
rect 485740 125604 485746 125656
rect 487890 125604 487896 125656
rect 487948 125644 487954 125656
rect 488442 125644 488448 125656
rect 487948 125616 488448 125644
rect 487948 125604 487954 125616
rect 488442 125604 488448 125616
rect 488500 125604 488506 125656
rect 490558 125604 490564 125656
rect 490616 125644 490622 125656
rect 491202 125644 491208 125656
rect 490616 125616 491208 125644
rect 490616 125604 490622 125616
rect 491202 125604 491208 125616
rect 491260 125604 491266 125656
rect 493318 125604 493324 125656
rect 493376 125644 493382 125656
rect 493962 125644 493968 125656
rect 493376 125616 493968 125644
rect 493376 125604 493382 125616
rect 493962 125604 493968 125616
rect 494020 125604 494026 125656
rect 496078 125604 496084 125656
rect 496136 125644 496142 125656
rect 496722 125644 496728 125656
rect 496136 125616 496728 125644
rect 496136 125604 496142 125616
rect 496722 125604 496728 125616
rect 496780 125604 496786 125656
rect 498746 125604 498752 125656
rect 498804 125644 498810 125656
rect 499482 125644 499488 125656
rect 498804 125616 499488 125644
rect 498804 125604 498810 125616
rect 499482 125604 499488 125616
rect 499540 125604 499546 125656
rect 501506 125604 501512 125656
rect 501564 125644 501570 125656
rect 502242 125644 502248 125656
rect 501564 125616 502248 125644
rect 501564 125604 501570 125616
rect 502242 125604 502248 125616
rect 502300 125604 502306 125656
rect 504174 125604 504180 125656
rect 504232 125644 504238 125656
rect 505002 125644 505008 125656
rect 504232 125616 505008 125644
rect 504232 125604 504238 125616
rect 505002 125604 505008 125616
rect 505060 125604 505066 125656
rect 506934 125604 506940 125656
rect 506992 125644 506998 125656
rect 507762 125644 507768 125656
rect 506992 125616 507768 125644
rect 506992 125604 506998 125616
rect 507762 125604 507768 125616
rect 507820 125604 507826 125656
rect 509602 125604 509608 125656
rect 509660 125644 509666 125656
rect 510522 125644 510528 125656
rect 509660 125616 510528 125644
rect 509660 125604 509666 125616
rect 510522 125604 510528 125616
rect 510580 125604 510586 125656
rect 511442 125604 511448 125656
rect 511500 125644 511506 125656
rect 511902 125644 511908 125656
rect 511500 125616 511908 125644
rect 511500 125604 511506 125616
rect 511902 125604 511908 125616
rect 511960 125604 511966 125656
rect 512362 125604 512368 125656
rect 512420 125644 512426 125656
rect 513282 125644 513288 125656
rect 512420 125616 513288 125644
rect 512420 125604 512426 125616
rect 513282 125604 513288 125616
rect 513340 125604 513346 125656
rect 514202 125604 514208 125656
rect 514260 125644 514266 125656
rect 514662 125644 514668 125656
rect 514260 125616 514668 125644
rect 514260 125604 514266 125616
rect 514662 125604 514668 125616
rect 514720 125604 514726 125656
rect 515398 125604 515404 125656
rect 515456 125644 515462 125656
rect 516042 125644 516048 125656
rect 515456 125616 516048 125644
rect 515456 125604 515462 125616
rect 516042 125604 516048 125616
rect 516100 125604 516106 125656
rect 507854 125400 507860 125452
rect 507912 125440 507918 125452
rect 550634 125440 550640 125452
rect 507912 125412 550640 125440
rect 507912 125400 507918 125412
rect 550634 125400 550640 125412
rect 550692 125400 550698 125452
rect 536834 125372 536840 125384
rect 485056 125344 536840 125372
rect 66220 125332 66226 125344
rect 536834 125332 536840 125344
rect 536892 125332 536898 125384
rect 33778 125264 33784 125316
rect 33836 125304 33842 125316
rect 85022 125304 85028 125316
rect 33836 125276 85028 125304
rect 33836 125264 33842 125276
rect 85022 125264 85028 125276
rect 85080 125264 85086 125316
rect 475194 125264 475200 125316
rect 475252 125304 475258 125316
rect 529934 125304 529940 125316
rect 475252 125276 529940 125304
rect 475252 125264 475258 125276
rect 529934 125264 529940 125276
rect 529992 125264 529998 125316
rect 18598 125196 18604 125248
rect 18656 125236 18662 125248
rect 69566 125236 69572 125248
rect 18656 125208 69572 125236
rect 18656 125196 18662 125208
rect 69566 125196 69572 125208
rect 69624 125196 69630 125248
rect 481634 125196 481640 125248
rect 481692 125236 481698 125248
rect 538214 125236 538220 125248
rect 481692 125208 538220 125236
rect 481692 125196 481698 125208
rect 538214 125196 538220 125208
rect 538272 125196 538278 125248
rect 62022 125128 62028 125180
rect 62080 125168 62086 125180
rect 115842 125168 115848 125180
rect 62080 125140 115848 125168
rect 62080 125128 62086 125140
rect 115842 125128 115848 125140
rect 115900 125128 115906 125180
rect 488810 125128 488816 125180
rect 488868 125168 488874 125180
rect 547874 125168 547880 125180
rect 488868 125140 547880 125168
rect 488868 125128 488874 125140
rect 547874 125128 547880 125140
rect 547932 125128 547938 125180
rect 55122 125060 55128 125112
rect 55180 125100 55186 125112
rect 110414 125100 110420 125112
rect 55180 125072 110420 125100
rect 55180 125060 55186 125072
rect 110414 125060 110420 125072
rect 110472 125060 110478 125112
rect 494238 125060 494244 125112
rect 494296 125100 494302 125112
rect 554774 125100 554780 125112
rect 494296 125072 554780 125100
rect 494296 125060 494302 125072
rect 554774 125060 554780 125072
rect 554832 125060 554838 125112
rect 52362 124992 52368 125044
rect 52420 125032 52426 125044
rect 107654 125032 107660 125044
rect 52420 125004 107660 125032
rect 52420 124992 52426 125004
rect 107654 124992 107660 125004
rect 107712 124992 107718 125044
rect 496906 124992 496912 125044
rect 496964 125032 496970 125044
rect 557534 125032 557540 125044
rect 496964 125004 557540 125032
rect 496964 124992 496970 125004
rect 557534 124992 557540 125004
rect 557592 124992 557598 125044
rect 48222 124924 48228 124976
rect 48280 124964 48286 124976
rect 104986 124964 104992 124976
rect 48280 124936 104992 124964
rect 48280 124924 48286 124936
rect 104986 124924 104992 124936
rect 105044 124924 105050 124976
rect 499666 124924 499672 124976
rect 499724 124964 499730 124976
rect 561674 124964 561680 124976
rect 499724 124936 561680 124964
rect 499724 124924 499730 124936
rect 561674 124924 561680 124936
rect 561732 124924 561738 124976
rect 4798 124856 4804 124908
rect 4856 124896 4862 124908
rect 70486 124896 70492 124908
rect 4856 124868 70492 124896
rect 4856 124856 4862 124868
rect 70486 124856 70492 124868
rect 70544 124856 70550 124908
rect 111610 124856 111616 124908
rect 111668 124896 111674 124908
rect 152550 124896 152556 124908
rect 111668 124868 152556 124896
rect 111668 124856 111674 124868
rect 152550 124856 152556 124868
rect 152608 124856 152614 124908
rect 502426 124856 502432 124908
rect 502484 124896 502490 124908
rect 564526 124896 564532 124908
rect 502484 124868 564532 124896
rect 502484 124856 502490 124868
rect 564526 124856 564532 124868
rect 564584 124856 564590 124908
rect 41322 123564 41328 123616
rect 41380 123604 41386 123616
rect 88242 123604 88248 123616
rect 41380 123576 88248 123604
rect 41380 123564 41386 123576
rect 88242 123564 88248 123576
rect 88300 123564 88306 123616
rect 37182 123496 37188 123548
rect 37240 123536 37246 123548
rect 88978 123536 88984 123548
rect 37240 123508 88984 123536
rect 37240 123496 37246 123508
rect 88978 123496 88984 123508
rect 89036 123496 89042 123548
rect 35158 123428 35164 123480
rect 35216 123468 35222 123480
rect 94130 123468 94136 123480
rect 35216 123440 94136 123468
rect 35216 123428 35222 123440
rect 94130 123428 94136 123440
rect 94188 123428 94194 123480
rect 507670 123428 507676 123480
rect 507728 123468 507734 123480
rect 572806 123468 572812 123480
rect 507728 123440 572812 123468
rect 507728 123428 507734 123440
rect 572806 123428 572812 123440
rect 572864 123428 572870 123480
rect 455230 90312 455236 90364
rect 455288 90352 455294 90364
rect 502334 90352 502340 90364
rect 455288 90324 502340 90352
rect 455288 90312 455294 90324
rect 502334 90312 502340 90324
rect 502392 90312 502398 90364
rect 3510 88952 3516 89004
rect 3568 88992 3574 89004
rect 67634 88992 67640 89004
rect 3568 88964 67640 88992
rect 3568 88952 3574 88964
rect 67634 88952 67640 88964
rect 67692 88952 67698 89004
rect 447778 88952 447784 89004
rect 447836 88992 447842 89004
rect 490006 88992 490012 89004
rect 447836 88964 490012 88992
rect 447836 88952 447842 88964
rect 490006 88952 490012 88964
rect 490064 88952 490070 89004
rect 533430 50328 533436 50380
rect 533488 50368 533494 50380
rect 575474 50368 575480 50380
rect 533488 50340 575480 50368
rect 533488 50328 533494 50340
rect 575474 50328 575480 50340
rect 575532 50328 575538 50380
rect 84102 48968 84108 49020
rect 84160 49008 84166 49020
rect 128998 49008 129004 49020
rect 84160 48980 129004 49008
rect 84160 48968 84166 48980
rect 128998 48968 129004 48980
rect 129056 48968 129062 49020
rect 102042 26868 102048 26920
rect 102100 26908 102106 26920
rect 126238 26908 126244 26920
rect 102100 26880 126244 26908
rect 102100 26868 102106 26880
rect 126238 26868 126244 26880
rect 126296 26868 126302 26920
rect 126882 26868 126888 26920
rect 126940 26908 126946 26920
rect 164234 26908 164240 26920
rect 126940 26880 164240 26908
rect 126940 26868 126946 26880
rect 164234 26868 164240 26880
rect 164292 26868 164298 26920
rect 459462 26868 459468 26920
rect 459520 26908 459526 26920
rect 507854 26908 507860 26920
rect 459520 26880 507860 26908
rect 459520 26868 459526 26880
rect 507854 26868 507860 26880
rect 507912 26868 507918 26920
rect 91002 18572 91008 18624
rect 91060 18612 91066 18624
rect 133138 18612 133144 18624
rect 91060 18584 133144 18612
rect 91060 18572 91066 18584
rect 133138 18572 133144 18584
rect 133196 18572 133202 18624
rect 133782 15920 133788 15972
rect 133840 15960 133846 15972
rect 169754 15960 169760 15972
rect 133840 15932 169760 15960
rect 133840 15920 133846 15932
rect 169754 15920 169760 15932
rect 169812 15920 169818 15972
rect 86862 15852 86868 15904
rect 86920 15892 86926 15904
rect 134150 15892 134156 15904
rect 86920 15864 134156 15892
rect 86920 15852 86926 15864
rect 134150 15852 134156 15864
rect 134208 15852 134214 15904
rect 439498 15852 439504 15904
rect 439556 15892 439562 15904
rect 481726 15892 481732 15904
rect 439556 15864 481732 15892
rect 439556 15852 439562 15864
rect 481726 15852 481732 15864
rect 481784 15852 481790 15904
rect 115842 11704 115848 11756
rect 115900 11744 115906 11756
rect 155954 11744 155960 11756
rect 115900 11716 155960 11744
rect 115900 11704 115906 11716
rect 155954 11704 155960 11716
rect 156012 11704 156018 11756
rect 386230 11704 386236 11756
rect 386288 11744 386294 11756
rect 412634 11744 412640 11756
rect 386288 11716 412640 11744
rect 386288 11704 386294 11716
rect 412634 11704 412640 11716
rect 412692 11704 412698 11756
rect 450538 11704 450544 11756
rect 450596 11744 450602 11756
rect 484762 11744 484768 11756
rect 450596 11716 484768 11744
rect 450596 11704 450602 11716
rect 484762 11704 484768 11716
rect 484820 11704 484826 11756
rect 77110 10276 77116 10328
rect 77168 10316 77174 10328
rect 125686 10316 125692 10328
rect 77168 10288 125692 10316
rect 77168 10276 77174 10288
rect 125686 10276 125692 10288
rect 125744 10276 125750 10328
rect 426250 10276 426256 10328
rect 426308 10316 426314 10328
rect 465810 10316 465816 10328
rect 426308 10288 465816 10316
rect 426308 10276 426314 10288
rect 465810 10276 465816 10288
rect 465868 10276 465874 10328
rect 469030 10276 469036 10328
rect 469088 10316 469094 10328
rect 520274 10316 520280 10328
rect 469088 10288 520280 10316
rect 469088 10276 469094 10288
rect 520274 10276 520280 10288
rect 520332 10276 520338 10328
rect 519538 9596 519544 9648
rect 519596 9636 519602 9648
rect 526622 9636 526628 9648
rect 519596 9608 526628 9636
rect 519596 9596 519602 9608
rect 526622 9596 526628 9608
rect 526680 9596 526686 9648
rect 444190 8984 444196 9036
rect 444248 9024 444254 9036
rect 488810 9024 488816 9036
rect 444248 8996 488816 9024
rect 444248 8984 444254 8996
rect 488810 8984 488816 8996
rect 488868 8984 488874 9036
rect 130562 8916 130568 8968
rect 130620 8956 130626 8968
rect 144178 8956 144184 8968
rect 130620 8928 144184 8956
rect 130620 8916 130626 8928
rect 144178 8916 144184 8928
rect 144236 8916 144242 8968
rect 178126 8956 178132 8968
rect 151786 8928 178132 8956
rect 143534 8848 143540 8900
rect 143592 8888 143598 8900
rect 151786 8888 151814 8928
rect 178126 8916 178132 8928
rect 178184 8916 178190 8968
rect 467742 8916 467748 8968
rect 467800 8956 467806 8968
rect 519538 8956 519544 8968
rect 467800 8928 519544 8956
rect 467800 8916 467806 8928
rect 519538 8916 519544 8928
rect 519596 8916 519602 8968
rect 526438 8916 526444 8968
rect 526496 8956 526502 8968
rect 544378 8956 544384 8968
rect 526496 8928 544384 8956
rect 526496 8916 526502 8928
rect 544378 8916 544384 8928
rect 544436 8916 544442 8968
rect 143592 8860 151814 8888
rect 143592 8848 143598 8860
rect 79686 7624 79692 7676
rect 79744 7664 79750 7676
rect 128446 7664 128452 7676
rect 79744 7636 128452 7664
rect 79744 7624 79750 7636
rect 128446 7624 128452 7636
rect 128504 7624 128510 7676
rect 464338 7624 464344 7676
rect 464396 7664 464402 7676
rect 506474 7664 506480 7676
rect 464396 7636 506480 7664
rect 464396 7624 464402 7636
rect 506474 7624 506480 7636
rect 506532 7624 506538 7676
rect 44266 7556 44272 7608
rect 44324 7596 44330 7608
rect 58618 7596 58624 7608
rect 44324 7568 58624 7596
rect 44324 7556 44330 7568
rect 58618 7556 58624 7568
rect 58676 7556 58682 7608
rect 112530 7596 112536 7608
rect 64846 7568 112536 7596
rect 58434 7488 58440 7540
rect 58492 7528 58498 7540
rect 64846 7528 64874 7568
rect 112530 7556 112536 7568
rect 112588 7556 112594 7608
rect 129366 7556 129372 7608
rect 129424 7596 129430 7608
rect 151078 7596 151084 7608
rect 129424 7568 151084 7596
rect 129424 7556 129430 7568
rect 151078 7556 151084 7568
rect 151136 7556 151142 7608
rect 372522 7556 372528 7608
rect 372580 7596 372586 7608
rect 395338 7596 395344 7608
rect 372580 7568 395344 7596
rect 372580 7556 372586 7568
rect 395338 7556 395344 7568
rect 395396 7556 395402 7608
rect 432598 7556 432604 7608
rect 432656 7596 432662 7608
rect 459186 7596 459192 7608
rect 432656 7568 459192 7596
rect 432656 7556 432662 7568
rect 459186 7556 459192 7568
rect 459244 7556 459250 7608
rect 489730 7556 489736 7608
rect 489788 7596 489794 7608
rect 549070 7596 549076 7608
rect 489788 7568 549076 7596
rect 489788 7556 489794 7568
rect 549070 7556 549076 7568
rect 549128 7556 549134 7608
rect 58492 7500 64874 7528
rect 58492 7488 58498 7500
rect 466362 6196 466368 6248
rect 466420 6236 466426 6248
rect 517146 6236 517152 6248
rect 466420 6208 517152 6236
rect 466420 6196 466426 6208
rect 517146 6196 517152 6208
rect 517204 6196 517210 6248
rect 473262 6128 473268 6180
rect 473320 6168 473326 6180
rect 527818 6168 527824 6180
rect 473320 6140 527824 6168
rect 473320 6128 473326 6140
rect 527818 6128 527824 6140
rect 527876 6128 527882 6180
rect 476758 5448 476764 5500
rect 476816 5488 476822 5500
rect 505370 5488 505376 5500
rect 476816 5460 505376 5488
rect 476816 5448 476822 5460
rect 505370 5448 505376 5460
rect 505428 5448 505434 5500
rect 471238 5380 471244 5432
rect 471296 5420 471302 5432
rect 510062 5420 510068 5432
rect 471296 5392 510068 5420
rect 471296 5380 471302 5392
rect 510062 5380 510068 5392
rect 510120 5380 510126 5432
rect 440142 5312 440148 5364
rect 440200 5352 440206 5364
rect 483014 5352 483020 5364
rect 440200 5324 483020 5352
rect 440200 5312 440206 5324
rect 483014 5312 483020 5324
rect 483072 5312 483078 5364
rect 483658 5312 483664 5364
rect 483716 5352 483722 5364
rect 499390 5352 499396 5364
rect 483716 5324 499396 5352
rect 483716 5312 483722 5324
rect 499390 5312 499396 5324
rect 499448 5312 499454 5364
rect 136450 5244 136456 5296
rect 136508 5284 136514 5296
rect 148318 5284 148324 5296
rect 136508 5256 148324 5284
rect 136508 5244 136514 5256
rect 148318 5244 148324 5256
rect 148376 5244 148382 5296
rect 446950 5244 446956 5296
rect 447008 5284 447014 5296
rect 485041 5287 485099 5293
rect 485041 5284 485053 5287
rect 447008 5256 485053 5284
rect 447008 5244 447014 5256
rect 485041 5253 485053 5256
rect 485087 5253 485099 5287
rect 485041 5247 485099 5253
rect 134150 5176 134156 5228
rect 134208 5216 134214 5228
rect 164878 5216 164884 5228
rect 134208 5188 164884 5216
rect 134208 5176 134214 5188
rect 164878 5176 164884 5188
rect 164936 5176 164942 5228
rect 407758 5176 407764 5228
rect 407816 5216 407822 5228
rect 416682 5216 416688 5228
rect 407816 5188 416688 5216
rect 407816 5176 407822 5188
rect 416682 5176 416688 5188
rect 416740 5176 416746 5228
rect 418798 5176 418804 5228
rect 418856 5216 418862 5228
rect 430850 5216 430856 5228
rect 418856 5188 430856 5216
rect 418856 5176 418862 5188
rect 430850 5176 430856 5188
rect 430908 5176 430914 5228
rect 448422 5176 448428 5228
rect 448480 5216 448486 5228
rect 494698 5216 494704 5228
rect 448480 5188 494704 5216
rect 448480 5176 448486 5188
rect 494698 5176 494704 5188
rect 494756 5176 494762 5228
rect 59630 5108 59636 5160
rect 59688 5148 59694 5160
rect 68278 5148 68284 5160
rect 59688 5120 68284 5148
rect 59688 5108 59694 5120
rect 68278 5108 68284 5120
rect 68336 5108 68342 5160
rect 69106 5108 69112 5160
rect 69164 5148 69170 5160
rect 112438 5148 112444 5160
rect 69164 5120 112444 5148
rect 69164 5108 69170 5120
rect 112438 5108 112444 5120
rect 112496 5108 112502 5160
rect 135346 5108 135352 5160
rect 135404 5148 135410 5160
rect 170398 5148 170404 5160
rect 135404 5120 170404 5148
rect 135404 5108 135410 5120
rect 170398 5108 170404 5120
rect 170456 5108 170462 5160
rect 392578 5108 392584 5160
rect 392636 5148 392642 5160
rect 420178 5148 420184 5160
rect 392636 5120 420184 5148
rect 392636 5108 392642 5120
rect 420178 5108 420184 5120
rect 420236 5108 420242 5160
rect 429838 5108 429844 5160
rect 429896 5148 429902 5160
rect 445018 5148 445024 5160
rect 429896 5120 445024 5148
rect 429896 5108 429902 5120
rect 445018 5108 445024 5120
rect 445076 5108 445082 5160
rect 453942 5108 453948 5160
rect 454000 5148 454006 5160
rect 501782 5148 501788 5160
rect 454000 5120 501788 5148
rect 454000 5108 454006 5120
rect 501782 5108 501788 5120
rect 501840 5108 501846 5160
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 53098 5080 53104 5092
rect 12400 5052 53104 5080
rect 12400 5040 12406 5052
rect 53098 5040 53104 5052
rect 53156 5040 53162 5092
rect 107838 5080 107844 5092
rect 53208 5052 107844 5080
rect 30098 4972 30104 5024
rect 30156 5012 30162 5024
rect 50338 5012 50344 5024
rect 30156 4984 50344 5012
rect 30156 4972 30162 4984
rect 50338 4972 50344 4984
rect 50396 4972 50402 5024
rect 52546 4972 52552 5024
rect 52604 5012 52610 5024
rect 53208 5012 53236 5052
rect 107838 5040 107844 5052
rect 107896 5040 107902 5092
rect 131758 5040 131764 5092
rect 131816 5080 131822 5092
rect 168650 5080 168656 5092
rect 131816 5052 168656 5080
rect 131816 5040 131822 5052
rect 168650 5040 168656 5052
rect 168708 5040 168714 5092
rect 403618 5040 403624 5092
rect 403676 5080 403682 5092
rect 434438 5080 434444 5092
rect 403676 5052 434444 5080
rect 403676 5040 403682 5052
rect 434438 5040 434444 5052
rect 434496 5040 434502 5092
rect 451182 5040 451188 5092
rect 451240 5080 451246 5092
rect 498194 5080 498200 5092
rect 451240 5052 498200 5080
rect 451240 5040 451246 5052
rect 498194 5040 498200 5052
rect 498252 5040 498258 5092
rect 504358 5040 504364 5092
rect 504416 5080 504422 5092
rect 513558 5080 513564 5092
rect 504416 5052 513564 5080
rect 504416 5040 504422 5052
rect 513558 5040 513564 5052
rect 513616 5040 513622 5092
rect 52604 4984 53236 5012
rect 53285 5015 53343 5021
rect 52604 4972 52610 4984
rect 53285 4981 53297 5015
rect 53331 5012 53343 5015
rect 104894 5012 104900 5024
rect 53331 4984 104900 5012
rect 53331 4981 53343 4984
rect 53285 4975 53343 4981
rect 104894 4972 104900 4984
rect 104952 4972 104958 5024
rect 108114 4972 108120 5024
rect 108172 5012 108178 5024
rect 150526 5012 150532 5024
rect 108172 4984 150532 5012
rect 108172 4972 108178 4984
rect 150526 4972 150532 4984
rect 150584 4972 150590 5024
rect 389818 4972 389824 5024
rect 389876 5012 389882 5024
rect 402514 5012 402520 5024
rect 389876 4984 402520 5012
rect 389876 4972 389882 4984
rect 402514 4972 402520 4984
rect 402572 4972 402578 5024
rect 406930 4972 406936 5024
rect 406988 5012 406994 5024
rect 441430 5012 441436 5024
rect 406988 4984 441436 5012
rect 406988 4972 406994 4984
rect 441430 4972 441436 4984
rect 441488 4972 441494 5024
rect 442258 4972 442264 5024
rect 442316 5012 442322 5024
rect 452102 5012 452108 5024
rect 442316 4984 452108 5012
rect 442316 4972 442322 4984
rect 452102 4972 452108 4984
rect 452160 4972 452166 5024
rect 475378 4972 475384 5024
rect 475436 5012 475442 5024
rect 524230 5012 524236 5024
rect 475436 4984 524236 5012
rect 475436 4972 475442 4984
rect 524230 4972 524236 4984
rect 524288 4972 524294 5024
rect 26510 4904 26516 4956
rect 26568 4944 26574 4956
rect 88426 4944 88432 4956
rect 26568 4916 88432 4944
rect 26568 4904 26574 4916
rect 88426 4904 88432 4916
rect 88484 4904 88490 4956
rect 93946 4904 93952 4956
rect 94004 4944 94010 4956
rect 139670 4944 139676 4956
rect 94004 4916 139676 4944
rect 94004 4904 94010 4916
rect 139670 4904 139676 4916
rect 139728 4904 139734 4956
rect 140038 4904 140044 4956
rect 140096 4944 140102 4956
rect 175274 4944 175280 4956
rect 140096 4916 175280 4944
rect 140096 4904 140102 4916
rect 175274 4904 175280 4916
rect 175332 4904 175338 4956
rect 375190 4904 375196 4956
rect 375248 4944 375254 4956
rect 398926 4944 398932 4956
rect 375248 4916 398932 4944
rect 375248 4904 375254 4916
rect 398926 4904 398932 4916
rect 398984 4904 398990 4956
rect 400858 4904 400864 4956
rect 400916 4944 400922 4956
rect 406010 4944 406016 4956
rect 400916 4916 406016 4944
rect 400916 4904 400922 4916
rect 406010 4904 406016 4916
rect 406068 4904 406074 4956
rect 412450 4904 412456 4956
rect 412508 4944 412514 4956
rect 448606 4944 448612 4956
rect 412508 4916 448612 4944
rect 412508 4904 412514 4916
rect 448606 4904 448612 4916
rect 448664 4904 448670 4956
rect 464982 4904 464988 4956
rect 465040 4944 465046 4956
rect 515950 4944 515956 4956
rect 465040 4916 515956 4944
rect 465040 4904 465046 4916
rect 515950 4904 515956 4916
rect 516008 4904 516014 4956
rect 522298 4904 522304 4956
rect 522356 4944 522362 4956
rect 533706 4944 533712 4956
rect 522356 4916 533712 4944
rect 522356 4904 522362 4916
rect 533706 4904 533712 4916
rect 533764 4904 533770 4956
rect 7650 4836 7656 4888
rect 7708 4876 7714 4888
rect 72418 4876 72424 4888
rect 7708 4848 72424 4876
rect 7708 4836 7714 4848
rect 72418 4836 72424 4848
rect 72476 4836 72482 4888
rect 97442 4836 97448 4888
rect 97500 4876 97506 4888
rect 142338 4876 142344 4888
rect 97500 4848 142344 4876
rect 97500 4836 97506 4848
rect 142338 4836 142344 4848
rect 142396 4836 142402 4888
rect 161290 4836 161296 4888
rect 161348 4876 161354 4888
rect 178678 4876 178684 4888
rect 161348 4848 178684 4876
rect 161348 4836 161354 4848
rect 178678 4836 178684 4848
rect 178736 4836 178742 4888
rect 383470 4836 383476 4888
rect 383528 4876 383534 4888
rect 409598 4876 409604 4888
rect 383528 4848 409604 4876
rect 383528 4836 383534 4848
rect 409598 4836 409604 4848
rect 409656 4836 409662 4888
rect 417970 4836 417976 4888
rect 418028 4876 418034 4888
rect 455690 4876 455696 4888
rect 418028 4848 455696 4876
rect 418028 4836 418034 4848
rect 455690 4836 455696 4848
rect 455748 4836 455754 4888
rect 462222 4836 462228 4888
rect 462280 4876 462286 4888
rect 512454 4876 512460 4888
rect 462280 4848 512460 4876
rect 462280 4836 462286 4848
rect 512454 4836 512460 4848
rect 512512 4836 512518 4888
rect 529198 4836 529204 4888
rect 529256 4876 529262 4888
rect 540790 4876 540796 4888
rect 529256 4848 540796 4876
rect 529256 4836 529262 4848
rect 540790 4836 540796 4848
rect 540848 4836 540854 4888
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 70394 4808 70400 4820
rect 4120 4780 70400 4808
rect 4120 4768 4126 4780
rect 70394 4768 70400 4780
rect 70452 4768 70458 4820
rect 72602 4768 72608 4820
rect 72660 4808 72666 4820
rect 122098 4808 122104 4820
rect 72660 4780 122104 4808
rect 72660 4768 72666 4780
rect 122098 4768 122104 4780
rect 122156 4768 122162 4820
rect 128170 4768 128176 4820
rect 128228 4808 128234 4820
rect 165706 4808 165712 4820
rect 128228 4780 165712 4808
rect 128228 4768 128234 4780
rect 165706 4768 165712 4780
rect 165764 4768 165770 4820
rect 371878 4768 371884 4820
rect 371936 4808 371942 4820
rect 391750 4808 391756 4820
rect 371936 4780 391756 4808
rect 371936 4768 371942 4780
rect 391750 4768 391756 4780
rect 391808 4768 391814 4820
rect 397270 4768 397276 4820
rect 397328 4808 397334 4820
rect 427262 4808 427268 4820
rect 397328 4780 427268 4808
rect 397328 4768 397334 4780
rect 427262 4768 427268 4780
rect 427320 4768 427326 4820
rect 431770 4768 431776 4820
rect 431828 4808 431834 4820
rect 473446 4808 473452 4820
rect 431828 4780 473452 4808
rect 431828 4768 431834 4780
rect 473446 4768 473452 4780
rect 473504 4768 473510 4820
rect 475930 4768 475936 4820
rect 475988 4808 475994 4820
rect 531314 4808 531320 4820
rect 475988 4780 531320 4808
rect 475988 4768 475994 4780
rect 531314 4768 531320 4780
rect 531372 4768 531378 4820
rect 536098 4768 536104 4820
rect 536156 4808 536162 4820
rect 541986 4808 541992 4820
rect 536156 4780 541992 4808
rect 536156 4768 536162 4780
rect 541986 4768 541992 4780
rect 542044 4768 542050 4820
rect 547138 4768 547144 4820
rect 547196 4808 547202 4820
rect 552658 4808 552664 4820
rect 547196 4780 552664 4808
rect 547196 4768 547202 4780
rect 552658 4768 552664 4780
rect 552716 4768 552722 4820
rect 50890 4700 50896 4752
rect 50948 4740 50954 4752
rect 53285 4743 53343 4749
rect 53285 4740 53297 4743
rect 50948 4712 53297 4740
rect 50948 4700 50954 4712
rect 53285 4709 53297 4712
rect 53331 4709 53343 4743
rect 53285 4703 53343 4709
rect 479518 4700 479524 4752
rect 479576 4740 479582 4752
rect 495894 4740 495900 4752
rect 479576 4712 495900 4740
rect 479576 4700 479582 4712
rect 495894 4700 495900 4712
rect 495952 4700 495958 4752
rect 471330 4632 471336 4684
rect 471388 4672 471394 4684
rect 480530 4672 480536 4684
rect 471388 4644 480536 4672
rect 471388 4632 471394 4644
rect 480530 4632 480536 4644
rect 480588 4632 480594 4684
rect 485041 4607 485099 4613
rect 485041 4573 485053 4607
rect 485087 4604 485099 4607
rect 492306 4604 492312 4616
rect 485087 4576 492312 4604
rect 485087 4573 485099 4576
rect 485041 4567 485099 4573
rect 492306 4564 492312 4576
rect 492364 4564 492370 4616
rect 421558 4428 421564 4480
rect 421616 4468 421622 4480
rect 423766 4468 423772 4480
rect 421616 4440 423772 4468
rect 421616 4428 421622 4440
rect 423766 4428 423772 4440
rect 423824 4428 423830 4480
rect 483014 4224 483020 4276
rect 483072 4264 483078 4276
rect 484026 4264 484032 4276
rect 483072 4236 484032 4264
rect 483072 4224 483078 4236
rect 484026 4224 484032 4236
rect 484084 4224 484090 4276
rect 126974 4156 126980 4208
rect 127032 4196 127038 4208
rect 130378 4196 130384 4208
rect 127032 4168 130384 4196
rect 127032 4156 127038 4168
rect 130378 4156 130384 4168
rect 130436 4156 130442 4208
rect 436738 4156 436744 4208
rect 436796 4196 436802 4208
rect 437934 4196 437940 4208
rect 436796 4168 437940 4196
rect 436796 4156 436802 4168
rect 437934 4156 437940 4168
rect 437992 4156 437998 4208
rect 461578 4156 461584 4208
rect 461636 4196 461642 4208
rect 462774 4196 462780 4208
rect 461636 4168 462780 4196
rect 461636 4156 461642 4168
rect 462774 4156 462780 4168
rect 462832 4156 462838 4208
rect 467098 4156 467104 4208
rect 467156 4196 467162 4208
rect 469858 4196 469864 4208
rect 467156 4168 469864 4196
rect 467156 4156 467162 4168
rect 469858 4156 469864 4168
rect 469916 4156 469922 4208
rect 472618 4156 472624 4208
rect 472676 4196 472682 4208
rect 476942 4196 476948 4208
rect 472676 4168 476948 4196
rect 472676 4156 472682 4168
rect 476942 4156 476948 4168
rect 477000 4156 477006 4208
rect 482278 4156 482284 4208
rect 482336 4196 482342 4208
rect 487614 4196 487620 4208
rect 482336 4168 487620 4196
rect 482336 4156 482342 4168
rect 487614 4156 487620 4168
rect 487672 4156 487678 4208
rect 520918 4156 520924 4208
rect 520976 4196 520982 4208
rect 523034 4196 523040 4208
rect 520976 4168 523040 4196
rect 520976 4156 520982 4168
rect 523034 4156 523040 4168
rect 523092 4156 523098 4208
rect 533338 4156 533344 4208
rect 533396 4196 533402 4208
rect 534902 4196 534908 4208
rect 533396 4168 534908 4196
rect 533396 4156 533402 4168
rect 534902 4156 534908 4168
rect 534960 4156 534966 4208
rect 542998 4156 543004 4208
rect 543056 4196 543062 4208
rect 545482 4196 545488 4208
rect 543056 4168 545488 4196
rect 543056 4156 543062 4168
rect 545482 4156 545488 4168
rect 545540 4156 545546 4208
rect 34790 4088 34796 4140
rect 34848 4128 34854 4140
rect 88981 4131 89039 4137
rect 88981 4128 88993 4131
rect 34848 4100 88993 4128
rect 34848 4088 34854 4100
rect 88981 4097 88993 4100
rect 89027 4097 89039 4131
rect 88981 4091 89039 4097
rect 89073 4131 89131 4137
rect 89073 4097 89085 4131
rect 89119 4128 89131 4131
rect 91649 4131 91707 4137
rect 91649 4128 91661 4131
rect 89119 4100 91661 4128
rect 89119 4097 89131 4100
rect 89073 4091 89131 4097
rect 91649 4097 91661 4100
rect 91695 4097 91707 4131
rect 91649 4091 91707 4097
rect 95421 4131 95479 4137
rect 95421 4097 95433 4131
rect 95467 4128 95479 4131
rect 99742 4128 99748 4140
rect 95467 4100 99748 4128
rect 95467 4097 95479 4100
rect 95421 4091 95479 4097
rect 99742 4088 99748 4100
rect 99800 4088 99806 4140
rect 102226 4088 102232 4140
rect 102284 4128 102290 4140
rect 146386 4128 146392 4140
rect 102284 4100 146392 4128
rect 102284 4088 102290 4100
rect 146386 4088 146392 4100
rect 146444 4088 146450 4140
rect 163682 4088 163688 4140
rect 163740 4128 163746 4140
rect 193214 4128 193220 4140
rect 163740 4100 193220 4128
rect 163740 4088 163746 4100
rect 193214 4088 193220 4100
rect 193272 4088 193278 4140
rect 219250 4088 219256 4140
rect 219308 4128 219314 4140
rect 220078 4128 220084 4140
rect 219308 4100 220084 4128
rect 219308 4088 219314 4100
rect 220078 4088 220084 4100
rect 220136 4088 220142 4140
rect 286594 4088 286600 4140
rect 286652 4128 286658 4140
rect 287146 4128 287152 4140
rect 286652 4100 287152 4128
rect 286652 4088 286658 4100
rect 287146 4088 287152 4100
rect 287204 4088 287210 4140
rect 296622 4088 296628 4140
rect 296680 4128 296686 4140
rect 297266 4128 297272 4140
rect 296680 4100 297272 4128
rect 296680 4088 296686 4100
rect 297266 4088 297272 4100
rect 297324 4088 297330 4140
rect 304902 4088 304908 4140
rect 304960 4128 304966 4140
rect 307938 4128 307944 4140
rect 304960 4100 307944 4128
rect 304960 4088 304966 4100
rect 307938 4088 307944 4100
rect 307996 4088 308002 4140
rect 331858 4088 331864 4140
rect 331916 4128 331922 4140
rect 336274 4128 336280 4140
rect 331916 4100 336280 4128
rect 331916 4088 331922 4100
rect 336274 4088 336280 4100
rect 336332 4088 336338 4140
rect 336642 4088 336648 4140
rect 336700 4128 336706 4140
rect 349246 4128 349252 4140
rect 336700 4100 349252 4128
rect 336700 4088 336706 4100
rect 349246 4088 349252 4100
rect 349304 4088 349310 4140
rect 356698 4088 356704 4140
rect 356756 4128 356762 4140
rect 374086 4128 374092 4140
rect 356756 4100 374092 4128
rect 356756 4088 356762 4100
rect 374086 4088 374092 4100
rect 374144 4088 374150 4140
rect 375282 4088 375288 4140
rect 375340 4128 375346 4140
rect 400030 4128 400036 4140
rect 375340 4100 400036 4128
rect 375340 4088 375346 4100
rect 400030 4088 400036 4100
rect 400088 4088 400094 4140
rect 400122 4088 400128 4140
rect 400180 4128 400186 4140
rect 432046 4128 432052 4140
rect 400180 4100 432052 4128
rect 400180 4088 400186 4100
rect 432046 4088 432052 4100
rect 432104 4088 432110 4140
rect 437293 4131 437351 4137
rect 437293 4128 437305 4131
rect 432984 4100 437305 4128
rect 38378 4020 38384 4072
rect 38436 4060 38442 4072
rect 96706 4060 96712 4072
rect 38436 4032 96712 4060
rect 38436 4020 38442 4032
rect 96706 4020 96712 4032
rect 96764 4020 96770 4072
rect 103330 4020 103336 4072
rect 103388 4060 103394 4072
rect 146294 4060 146300 4072
rect 103388 4032 146300 4060
rect 103388 4020 103394 4032
rect 146294 4020 146300 4032
rect 146352 4020 146358 4072
rect 164878 4020 164884 4072
rect 164936 4060 164942 4072
rect 194686 4060 194692 4072
rect 164936 4032 194692 4060
rect 164936 4020 164942 4032
rect 194686 4020 194692 4032
rect 194744 4020 194750 4072
rect 242894 4020 242900 4072
rect 242952 4060 242958 4072
rect 249150 4060 249156 4072
rect 242952 4032 249156 4060
rect 242952 4020 242958 4032
rect 249150 4020 249156 4032
rect 249208 4020 249214 4072
rect 253474 4020 253480 4072
rect 253532 4060 253538 4072
rect 260098 4060 260104 4072
rect 253532 4032 260104 4060
rect 253532 4020 253538 4032
rect 260098 4020 260104 4032
rect 260156 4020 260162 4072
rect 273622 4020 273628 4072
rect 273680 4060 273686 4072
rect 277486 4060 277492 4072
rect 273680 4032 277492 4060
rect 273680 4020 273686 4032
rect 277486 4020 277492 4032
rect 277544 4020 277550 4072
rect 325510 4020 325516 4072
rect 325568 4060 325574 4072
rect 333882 4060 333888 4072
rect 325568 4032 333888 4060
rect 325568 4020 325574 4032
rect 333882 4020 333888 4032
rect 333940 4020 333946 4072
rect 339402 4020 339408 4072
rect 339460 4060 339466 4072
rect 352834 4060 352840 4072
rect 339460 4032 352840 4060
rect 339460 4020 339466 4032
rect 352834 4020 352840 4032
rect 352892 4020 352898 4072
rect 354582 4020 354588 4072
rect 354640 4060 354646 4072
rect 371694 4060 371700 4072
rect 354640 4032 371700 4060
rect 354640 4020 354646 4032
rect 371694 4020 371700 4032
rect 371752 4020 371758 4072
rect 373810 4020 373816 4072
rect 373868 4060 373874 4072
rect 397730 4060 397736 4072
rect 373868 4032 397736 4060
rect 373868 4020 373874 4032
rect 397730 4020 397736 4032
rect 397788 4020 397794 4072
rect 402882 4020 402888 4072
rect 402940 4060 402946 4072
rect 432877 4063 432935 4069
rect 432877 4060 432889 4063
rect 402940 4032 432889 4060
rect 402940 4020 402946 4032
rect 432877 4029 432889 4032
rect 432923 4029 432935 4063
rect 432877 4023 432935 4029
rect 21818 3952 21824 4004
rect 21876 3992 21882 4004
rect 33778 3992 33784 4004
rect 21876 3964 33784 3992
rect 21876 3952 21882 3964
rect 33778 3952 33784 3964
rect 33836 3952 33842 4004
rect 39574 3952 39580 4004
rect 39632 3992 39638 4004
rect 97994 3992 98000 4004
rect 39632 3964 98000 3992
rect 39632 3952 39638 3964
rect 97994 3952 98000 3964
rect 98052 3952 98058 4004
rect 102410 3992 102416 4004
rect 98104 3964 102416 3992
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 32398 3924 32404 3936
rect 17092 3896 32404 3924
rect 17092 3884 17098 3896
rect 32398 3884 32404 3896
rect 32456 3884 32462 3936
rect 35986 3884 35992 3936
rect 36044 3924 36050 3936
rect 88889 3927 88947 3933
rect 88889 3924 88901 3927
rect 36044 3896 88901 3924
rect 36044 3884 36050 3896
rect 88889 3893 88901 3896
rect 88935 3893 88947 3927
rect 88889 3887 88947 3893
rect 88981 3927 89039 3933
rect 88981 3893 88993 3927
rect 89027 3924 89039 3927
rect 93854 3924 93860 3936
rect 89027 3896 93860 3924
rect 89027 3893 89039 3896
rect 88981 3887 89039 3893
rect 93854 3884 93860 3896
rect 93912 3884 93918 3936
rect 95513 3927 95571 3933
rect 95513 3893 95525 3927
rect 95559 3924 95571 3927
rect 98104 3924 98132 3964
rect 102410 3952 102416 3964
rect 102468 3952 102474 4004
rect 105722 3952 105728 4004
rect 105780 3992 105786 4004
rect 149146 3992 149152 4004
rect 105780 3964 149152 3992
rect 105780 3952 105786 3964
rect 149146 3952 149152 3964
rect 149204 3952 149210 4004
rect 155402 3952 155408 4004
rect 155460 3992 155466 4004
rect 186406 3992 186412 4004
rect 155460 3964 186412 3992
rect 155460 3952 155466 3964
rect 186406 3952 186412 3964
rect 186464 3952 186470 4004
rect 324222 3952 324228 4004
rect 324280 3992 324286 4004
rect 332686 3992 332692 4004
rect 324280 3964 332692 3992
rect 324280 3952 324286 3964
rect 332686 3952 332692 3964
rect 332744 3952 332750 4004
rect 342070 3952 342076 4004
rect 342128 3992 342134 4004
rect 355226 3992 355232 4004
rect 342128 3964 355232 3992
rect 342128 3952 342134 3964
rect 355226 3952 355232 3964
rect 355284 3952 355290 4004
rect 361482 3952 361488 4004
rect 361540 3992 361546 4004
rect 381170 3992 381176 4004
rect 361540 3964 381176 3992
rect 361540 3952 361546 3964
rect 381170 3952 381176 3964
rect 381228 3952 381234 4004
rect 382182 3952 382188 4004
rect 382240 3992 382246 4004
rect 382240 3964 405596 3992
rect 382240 3952 382246 3964
rect 95559 3896 98132 3924
rect 95559 3893 95571 3896
rect 95513 3887 95571 3893
rect 99834 3884 99840 3936
rect 99892 3924 99898 3936
rect 144914 3924 144920 3936
rect 99892 3896 144920 3924
rect 99892 3884 99898 3896
rect 144914 3884 144920 3896
rect 144972 3884 144978 3936
rect 151814 3884 151820 3936
rect 151872 3924 151878 3936
rect 183646 3924 183652 3936
rect 151872 3896 183652 3924
rect 151872 3884 151878 3896
rect 183646 3884 183652 3896
rect 183704 3884 183710 3936
rect 200298 3884 200304 3936
rect 200356 3924 200362 3936
rect 220906 3924 220912 3936
rect 200356 3896 220912 3924
rect 200356 3884 200362 3896
rect 220906 3884 220912 3896
rect 220964 3884 220970 3936
rect 328362 3884 328368 3936
rect 328420 3924 328426 3936
rect 337470 3924 337476 3936
rect 328420 3896 337476 3924
rect 328420 3884 328426 3896
rect 337470 3884 337476 3896
rect 337528 3884 337534 3936
rect 345658 3884 345664 3936
rect 345716 3924 345722 3936
rect 359918 3924 359924 3936
rect 345716 3896 359924 3924
rect 345716 3884 345722 3896
rect 359918 3884 359924 3896
rect 359976 3884 359982 3936
rect 360102 3884 360108 3936
rect 360160 3924 360166 3936
rect 378870 3924 378876 3936
rect 360160 3896 378876 3924
rect 360160 3884 360166 3896
rect 378870 3884 378876 3896
rect 378928 3884 378934 3936
rect 379422 3884 379428 3936
rect 379480 3924 379486 3936
rect 404814 3924 404820 3936
rect 379480 3896 404820 3924
rect 379480 3884 379486 3896
rect 404814 3884 404820 3896
rect 404872 3884 404878 3936
rect 5258 3816 5264 3868
rect 5316 3856 5322 3868
rect 7558 3856 7564 3868
rect 5316 3828 7564 3856
rect 5316 3816 5322 3828
rect 7558 3816 7564 3828
rect 7616 3816 7622 3868
rect 31294 3816 31300 3868
rect 31352 3856 31358 3868
rect 91278 3856 91284 3868
rect 31352 3828 91284 3856
rect 31352 3816 31358 3828
rect 91278 3816 91284 3828
rect 91336 3816 91342 3868
rect 91554 3816 91560 3868
rect 91612 3856 91618 3868
rect 138014 3856 138020 3868
rect 91612 3828 138020 3856
rect 91612 3816 91618 3828
rect 138014 3816 138020 3828
rect 138072 3816 138078 3868
rect 156598 3816 156604 3868
rect 156656 3856 156662 3868
rect 187694 3856 187700 3868
rect 156656 3828 187700 3856
rect 156656 3816 156662 3828
rect 187694 3816 187700 3828
rect 187752 3816 187758 3868
rect 193214 3816 193220 3868
rect 193272 3856 193278 3868
rect 215386 3856 215392 3868
rect 193272 3828 215392 3856
rect 193272 3816 193278 3828
rect 215386 3816 215392 3828
rect 215444 3816 215450 3868
rect 332502 3816 332508 3868
rect 332560 3856 332566 3868
rect 343358 3856 343364 3868
rect 332560 3828 343364 3856
rect 332560 3816 332566 3828
rect 343358 3816 343364 3828
rect 343416 3816 343422 3868
rect 343542 3816 343548 3868
rect 343600 3856 343606 3868
rect 357526 3856 357532 3868
rect 343600 3828 357532 3856
rect 343600 3816 343606 3828
rect 357526 3816 357532 3828
rect 357584 3816 357590 3868
rect 358722 3816 358728 3868
rect 358780 3856 358786 3868
rect 377674 3856 377680 3868
rect 358780 3828 377680 3856
rect 358780 3816 358786 3828
rect 377674 3816 377680 3828
rect 377732 3816 377738 3868
rect 378042 3816 378048 3868
rect 378100 3856 378106 3868
rect 403618 3856 403624 3868
rect 378100 3828 403624 3856
rect 378100 3816 378106 3828
rect 403618 3816 403624 3828
rect 403676 3816 403682 3868
rect 405568 3856 405596 3964
rect 407022 3952 407028 4004
rect 407080 3992 407086 4004
rect 432984 3992 433012 4100
rect 437293 4097 437305 4100
rect 437339 4097 437351 4131
rect 437293 4091 437351 4097
rect 437382 4088 437388 4140
rect 437440 4128 437446 4140
rect 479334 4128 479340 4140
rect 437440 4100 479340 4128
rect 437440 4088 437446 4100
rect 479334 4088 479340 4100
rect 479392 4088 479398 4140
rect 498010 4088 498016 4140
rect 498068 4128 498074 4140
rect 559742 4128 559748 4140
rect 498068 4100 559748 4128
rect 498068 4088 498074 4100
rect 559742 4088 559748 4100
rect 559800 4088 559806 4140
rect 433061 4063 433119 4069
rect 433061 4029 433073 4063
rect 433107 4060 433119 4063
rect 435542 4060 435548 4072
rect 433107 4032 435548 4060
rect 433107 4029 433119 4032
rect 433061 4023 433119 4029
rect 435542 4020 435548 4032
rect 435600 4020 435606 4072
rect 436002 4020 436008 4072
rect 436060 4060 436066 4072
rect 478138 4060 478144 4072
rect 436060 4032 478144 4060
rect 436060 4020 436066 4032
rect 478138 4020 478144 4032
rect 478196 4020 478202 4072
rect 495250 4020 495256 4072
rect 495308 4060 495314 4072
rect 556154 4060 556160 4072
rect 495308 4032 556160 4060
rect 495308 4020 495314 4032
rect 556154 4020 556160 4032
rect 556212 4020 556218 4072
rect 407080 3964 433012 3992
rect 407080 3952 407086 3964
rect 433150 3952 433156 4004
rect 433208 3992 433214 4004
rect 436925 3995 436983 4001
rect 436925 3992 436937 3995
rect 433208 3964 436937 3992
rect 433208 3952 433214 3964
rect 436925 3961 436937 3964
rect 436971 3961 436983 3995
rect 436925 3955 436983 3961
rect 437293 3995 437351 4001
rect 437293 3961 437305 3995
rect 437339 3992 437351 3995
rect 440326 3992 440332 4004
rect 437339 3964 440332 3992
rect 437339 3961 437351 3964
rect 437293 3955 437351 3961
rect 440326 3952 440332 3964
rect 440384 3952 440390 4004
rect 441522 3952 441528 4004
rect 441580 3992 441586 4004
rect 486418 3992 486424 4004
rect 441580 3964 486424 3992
rect 441580 3952 441586 3964
rect 486418 3952 486424 3964
rect 486476 3952 486482 4004
rect 502242 3952 502248 4004
rect 502300 3992 502306 4004
rect 564434 3992 564440 4004
rect 502300 3964 564440 3992
rect 502300 3952 502306 3964
rect 564434 3952 564440 3964
rect 564492 3952 564498 4004
rect 405642 3884 405648 3936
rect 405700 3924 405706 3936
rect 439130 3924 439136 3936
rect 405700 3896 439136 3924
rect 405700 3884 405706 3896
rect 439130 3884 439136 3896
rect 439188 3884 439194 3936
rect 444282 3884 444288 3936
rect 444340 3924 444346 3936
rect 489914 3924 489920 3936
rect 444340 3896 489920 3924
rect 444340 3884 444346 3896
rect 489914 3884 489920 3896
rect 489972 3884 489978 3936
rect 505002 3884 505008 3936
rect 505060 3924 505066 3936
rect 568022 3924 568028 3936
rect 505060 3896 568028 3924
rect 505060 3884 505066 3896
rect 568022 3884 568028 3896
rect 568080 3884 568086 3936
rect 408218 3856 408224 3868
rect 405568 3828 408224 3856
rect 408218 3816 408224 3828
rect 408276 3816 408282 3868
rect 408310 3816 408316 3868
rect 408368 3856 408374 3868
rect 442626 3856 442632 3868
rect 408368 3828 442632 3856
rect 408368 3816 408374 3828
rect 442626 3816 442632 3828
rect 442684 3816 442690 3868
rect 447042 3816 447048 3868
rect 447100 3856 447106 3868
rect 493502 3856 493508 3868
rect 447100 3828 493508 3856
rect 447100 3816 447106 3828
rect 493502 3816 493508 3828
rect 493560 3816 493566 3868
rect 500770 3816 500776 3868
rect 500828 3856 500834 3868
rect 563238 3856 563244 3868
rect 500828 3828 563244 3856
rect 500828 3816 500834 3828
rect 563238 3816 563244 3828
rect 563296 3816 563302 3868
rect 14734 3748 14740 3800
rect 14792 3788 14798 3800
rect 17218 3788 17224 3800
rect 14792 3760 17224 3788
rect 14792 3748 14798 3760
rect 17218 3748 17224 3760
rect 17276 3748 17282 3800
rect 32398 3748 32404 3800
rect 32456 3788 32462 3800
rect 92474 3788 92480 3800
rect 32456 3760 92480 3788
rect 32456 3748 32462 3760
rect 92474 3748 92480 3760
rect 92532 3748 92538 3800
rect 92750 3748 92756 3800
rect 92808 3788 92814 3800
rect 93762 3788 93768 3800
rect 92808 3760 93768 3788
rect 92808 3748 92814 3760
rect 93762 3748 93768 3760
rect 93820 3748 93826 3800
rect 95142 3748 95148 3800
rect 95200 3788 95206 3800
rect 140774 3788 140780 3800
rect 95200 3760 140780 3788
rect 95200 3748 95206 3760
rect 140774 3748 140780 3760
rect 140832 3748 140838 3800
rect 149514 3748 149520 3800
rect 149572 3788 149578 3800
rect 172977 3791 173035 3797
rect 172977 3788 172989 3791
rect 149572 3760 172989 3788
rect 149572 3748 149578 3760
rect 172977 3757 172989 3760
rect 173023 3757 173035 3791
rect 172977 3751 173035 3757
rect 173069 3791 173127 3797
rect 173069 3757 173081 3791
rect 173115 3788 173127 3791
rect 176838 3788 176844 3800
rect 173115 3760 176844 3788
rect 173115 3757 173127 3760
rect 173069 3751 173127 3757
rect 176838 3748 176844 3760
rect 176896 3748 176902 3800
rect 180242 3748 180248 3800
rect 180300 3788 180306 3800
rect 180702 3788 180708 3800
rect 180300 3760 180708 3788
rect 180300 3748 180306 3760
rect 180702 3748 180708 3760
rect 180760 3748 180766 3800
rect 196802 3748 196808 3800
rect 196860 3788 196866 3800
rect 218146 3788 218152 3800
rect 196860 3760 218152 3788
rect 196860 3748 196866 3760
rect 218146 3748 218152 3760
rect 218204 3748 218210 3800
rect 322842 3748 322848 3800
rect 322900 3788 322906 3800
rect 330386 3788 330392 3800
rect 322900 3760 330392 3788
rect 322900 3748 322906 3760
rect 330386 3748 330392 3760
rect 330444 3748 330450 3800
rect 331122 3748 331128 3800
rect 331180 3788 331186 3800
rect 340966 3788 340972 3800
rect 331180 3760 340972 3788
rect 331180 3748 331186 3760
rect 340966 3748 340972 3760
rect 341024 3748 341030 3800
rect 342162 3748 342168 3800
rect 342220 3788 342226 3800
rect 356330 3788 356336 3800
rect 342220 3760 356336 3788
rect 342220 3748 342226 3760
rect 356330 3748 356336 3760
rect 356388 3748 356394 3800
rect 362862 3748 362868 3800
rect 362920 3788 362926 3800
rect 382366 3788 382372 3800
rect 362920 3760 382372 3788
rect 362920 3748 362926 3760
rect 382366 3748 382372 3760
rect 382424 3748 382430 3800
rect 383562 3748 383568 3800
rect 383620 3788 383626 3800
rect 410794 3788 410800 3800
rect 383620 3760 410800 3788
rect 383620 3748 383626 3760
rect 410794 3748 410800 3760
rect 410852 3748 410858 3800
rect 411162 3748 411168 3800
rect 411220 3788 411226 3800
rect 446214 3788 446220 3800
rect 411220 3760 446220 3788
rect 411220 3748 411226 3760
rect 446214 3748 446220 3760
rect 446272 3748 446278 3800
rect 449710 3748 449716 3800
rect 449768 3788 449774 3800
rect 497090 3788 497096 3800
rect 449768 3760 497096 3788
rect 449768 3748 449774 3760
rect 497090 3748 497096 3760
rect 497148 3748 497154 3800
rect 503530 3748 503536 3800
rect 503588 3788 503594 3800
rect 566826 3788 566832 3800
rect 503588 3760 566832 3788
rect 503588 3748 503594 3760
rect 566826 3748 566832 3760
rect 566884 3748 566890 3800
rect 25314 3680 25320 3732
rect 25372 3720 25378 3732
rect 25372 3692 83136 3720
rect 25372 3680 25378 3692
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 19484 3624 26234 3652
rect 19484 3612 19490 3624
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 14458 3584 14464 3596
rect 6512 3556 14464 3584
rect 6512 3544 6518 3556
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 18598 3584 18604 3596
rect 16546 3556 18604 3584
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4798 3516 4804 3528
rect 2924 3488 4804 3516
rect 2924 3476 2930 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 16546 3516 16574 3556
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 23014 3544 23020 3596
rect 23072 3584 23078 3596
rect 26206 3584 26234 3624
rect 27706 3612 27712 3664
rect 27764 3652 27770 3664
rect 29638 3652 29644 3664
rect 27764 3624 29644 3652
rect 27764 3612 27770 3624
rect 29638 3612 29644 3624
rect 29696 3612 29702 3664
rect 33594 3612 33600 3664
rect 33652 3652 33658 3664
rect 35158 3652 35164 3664
rect 33652 3624 35164 3652
rect 33652 3612 33658 3624
rect 35158 3612 35164 3624
rect 35216 3612 35222 3664
rect 35253 3655 35311 3661
rect 35253 3621 35265 3655
rect 35299 3652 35311 3655
rect 83001 3655 83059 3661
rect 83001 3652 83013 3655
rect 35299 3624 83013 3652
rect 35299 3621 35311 3624
rect 35253 3615 35311 3621
rect 83001 3621 83013 3624
rect 83047 3621 83059 3655
rect 83001 3615 83059 3621
rect 74813 3587 74871 3593
rect 74813 3584 74825 3587
rect 23072 3556 25636 3584
rect 26206 3556 74825 3584
rect 23072 3544 23078 3556
rect 6886 3488 16574 3516
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 6886 3448 6914 3488
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 21358 3516 21364 3528
rect 18288 3488 21364 3516
rect 18288 3476 18294 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 25498 3516 25504 3528
rect 24268 3488 25504 3516
rect 24268 3476 24274 3488
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 25608 3516 25636 3556
rect 74813 3553 74825 3556
rect 74859 3553 74871 3587
rect 74813 3547 74871 3553
rect 74905 3587 74963 3593
rect 74905 3553 74917 3587
rect 74951 3584 74963 3587
rect 76098 3584 76104 3596
rect 74951 3556 76104 3584
rect 74951 3553 74963 3556
rect 74905 3547 74963 3553
rect 76098 3544 76104 3556
rect 76156 3544 76162 3596
rect 76193 3587 76251 3593
rect 76193 3553 76205 3587
rect 76239 3584 76251 3587
rect 82906 3584 82912 3596
rect 76239 3556 82912 3584
rect 76239 3553 76251 3556
rect 76193 3547 76251 3553
rect 82906 3544 82912 3556
rect 82964 3544 82970 3596
rect 83108 3584 83136 3692
rect 84470 3680 84476 3732
rect 84528 3720 84534 3732
rect 91557 3723 91615 3729
rect 91557 3720 91569 3723
rect 84528 3692 91569 3720
rect 84528 3680 84534 3692
rect 91557 3689 91569 3692
rect 91603 3689 91615 3723
rect 91557 3683 91615 3689
rect 91649 3723 91707 3729
rect 91649 3689 91661 3723
rect 91695 3720 91707 3723
rect 123294 3720 123300 3732
rect 91695 3692 123300 3720
rect 91695 3689 91707 3692
rect 91649 3683 91707 3689
rect 123294 3680 123300 3692
rect 123352 3680 123358 3732
rect 123389 3723 123447 3729
rect 123389 3689 123401 3723
rect 123435 3720 123447 3723
rect 132586 3720 132592 3732
rect 123435 3692 132592 3720
rect 123435 3689 123447 3692
rect 123389 3683 123447 3689
rect 132586 3680 132592 3692
rect 132644 3680 132650 3732
rect 132865 3723 132923 3729
rect 132865 3689 132877 3723
rect 132911 3720 132923 3723
rect 136726 3720 136732 3732
rect 132911 3692 136732 3720
rect 132911 3689 132923 3692
rect 132865 3683 132923 3689
rect 136726 3680 136732 3692
rect 136784 3680 136790 3732
rect 142341 3723 142399 3729
rect 142341 3689 142353 3723
rect 142387 3720 142399 3723
rect 149054 3720 149060 3732
rect 142387 3692 149060 3720
rect 142387 3689 142399 3692
rect 142341 3683 142399 3689
rect 149054 3680 149060 3692
rect 149112 3680 149118 3732
rect 150618 3680 150624 3732
rect 150676 3720 150682 3732
rect 183554 3720 183560 3732
rect 150676 3692 183560 3720
rect 150676 3680 150682 3692
rect 183554 3680 183560 3692
rect 183612 3680 183618 3732
rect 189718 3680 189724 3732
rect 189776 3720 189782 3732
rect 212626 3720 212632 3732
rect 189776 3692 212632 3720
rect 189776 3680 189782 3692
rect 212626 3680 212632 3692
rect 212684 3680 212690 3732
rect 317322 3680 317328 3732
rect 317380 3720 317386 3732
rect 324406 3720 324412 3732
rect 317380 3692 324412 3720
rect 317380 3680 317386 3692
rect 324406 3680 324412 3692
rect 324464 3680 324470 3732
rect 329742 3680 329748 3732
rect 329800 3720 329806 3732
rect 339862 3720 339868 3732
rect 329800 3692 339868 3720
rect 329800 3680 329806 3692
rect 339862 3680 339868 3692
rect 339920 3680 339926 3732
rect 340782 3680 340788 3732
rect 340840 3720 340846 3732
rect 354030 3720 354036 3732
rect 340840 3692 354036 3720
rect 340840 3680 340846 3692
rect 354030 3680 354036 3692
rect 354088 3680 354094 3732
rect 354490 3680 354496 3732
rect 354548 3720 354554 3732
rect 372890 3720 372896 3732
rect 354548 3692 372896 3720
rect 354548 3680 354554 3692
rect 372890 3680 372896 3692
rect 372948 3680 372954 3732
rect 380802 3680 380808 3732
rect 380860 3720 380866 3732
rect 407206 3720 407212 3732
rect 380860 3692 407212 3720
rect 380860 3680 380866 3692
rect 407206 3680 407212 3692
rect 407264 3680 407270 3732
rect 407301 3723 407359 3729
rect 407301 3689 407313 3723
rect 407347 3720 407359 3723
rect 412085 3723 412143 3729
rect 412085 3720 412097 3723
rect 407347 3692 412097 3720
rect 407347 3689 407359 3692
rect 407301 3683 407359 3689
rect 412085 3689 412097 3692
rect 412131 3689 412143 3723
rect 412085 3683 412143 3689
rect 413922 3680 413928 3732
rect 413980 3720 413986 3732
rect 417973 3723 418031 3729
rect 417973 3720 417985 3723
rect 413980 3692 417985 3720
rect 413980 3680 413986 3692
rect 417973 3689 417985 3692
rect 418019 3689 418031 3723
rect 417973 3683 418031 3689
rect 418062 3680 418068 3732
rect 418120 3720 418126 3732
rect 421653 3723 421711 3729
rect 418120 3692 421604 3720
rect 418120 3680 418126 3692
rect 83185 3655 83243 3661
rect 83185 3621 83197 3655
rect 83231 3652 83243 3655
rect 88889 3655 88947 3661
rect 83231 3624 87184 3652
rect 83231 3621 83243 3624
rect 83185 3615 83243 3621
rect 87046 3584 87052 3596
rect 83108 3556 87052 3584
rect 87046 3544 87052 3556
rect 87104 3544 87110 3596
rect 85758 3516 85764 3528
rect 25608 3488 85764 3516
rect 85758 3476 85764 3488
rect 85816 3476 85822 3528
rect 87156 3516 87184 3624
rect 88889 3621 88901 3655
rect 88935 3652 88947 3655
rect 95234 3652 95240 3664
rect 88935 3624 95240 3652
rect 88935 3621 88947 3624
rect 88889 3615 88947 3621
rect 95234 3612 95240 3624
rect 95292 3612 95298 3664
rect 98638 3612 98644 3664
rect 98696 3652 98702 3664
rect 99282 3652 99288 3664
rect 98696 3624 99288 3652
rect 98696 3612 98702 3624
rect 99282 3612 99288 3624
rect 99340 3612 99346 3664
rect 101030 3612 101036 3664
rect 101088 3652 101094 3664
rect 102042 3652 102048 3664
rect 101088 3624 102048 3652
rect 101088 3612 101094 3624
rect 102042 3612 102048 3624
rect 102100 3612 102106 3664
rect 102137 3655 102195 3661
rect 102137 3621 102149 3655
rect 102183 3652 102195 3655
rect 142154 3652 142160 3664
rect 102183 3624 142160 3652
rect 102183 3621 102195 3624
rect 102137 3615 102195 3621
rect 142154 3612 142160 3624
rect 142212 3612 142218 3664
rect 147122 3612 147128 3664
rect 147180 3652 147186 3664
rect 147180 3624 173848 3652
rect 147180 3612 147186 3624
rect 87966 3544 87972 3596
rect 88024 3584 88030 3596
rect 135254 3584 135260 3596
rect 88024 3556 135260 3584
rect 88024 3544 88030 3556
rect 135254 3544 135260 3556
rect 135312 3544 135318 3596
rect 145926 3544 145932 3596
rect 145984 3584 145990 3596
rect 173713 3587 173771 3593
rect 173713 3584 173725 3587
rect 145984 3556 173725 3584
rect 145984 3544 145990 3556
rect 173713 3553 173725 3556
rect 173759 3553 173771 3587
rect 173820 3584 173848 3624
rect 174262 3612 174268 3664
rect 174320 3652 174326 3664
rect 181438 3652 181444 3664
rect 174320 3624 181444 3652
rect 174320 3612 174326 3624
rect 181438 3612 181444 3624
rect 181496 3612 181502 3664
rect 182542 3612 182548 3664
rect 182600 3652 182606 3664
rect 187053 3655 187111 3661
rect 187053 3652 187065 3655
rect 182600 3624 187065 3652
rect 182600 3612 182606 3624
rect 187053 3621 187065 3624
rect 187099 3621 187111 3655
rect 187053 3615 187111 3621
rect 188522 3612 188528 3664
rect 188580 3652 188586 3664
rect 188982 3652 188988 3664
rect 188580 3624 188988 3652
rect 188580 3612 188586 3624
rect 188982 3612 188988 3624
rect 189040 3612 189046 3664
rect 208486 3652 208492 3664
rect 201328 3624 208492 3652
rect 180978 3584 180984 3596
rect 173820 3556 180984 3584
rect 173713 3547 173771 3553
rect 180978 3544 180984 3556
rect 181036 3544 181042 3596
rect 186130 3544 186136 3596
rect 186188 3584 186194 3596
rect 200117 3587 200175 3593
rect 200117 3584 200129 3587
rect 186188 3556 200129 3584
rect 186188 3544 186194 3556
rect 200117 3553 200129 3556
rect 200163 3553 200175 3587
rect 200117 3547 200175 3553
rect 89714 3516 89720 3528
rect 87156 3488 89720 3516
rect 89714 3476 89720 3488
rect 89772 3476 89778 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 132865 3519 132923 3525
rect 132865 3516 132877 3519
rect 91480 3488 132877 3516
rect 1728 3420 6914 3448
rect 1728 3408 1734 3420
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 74905 3451 74963 3457
rect 74905 3448 74917 3451
rect 11204 3420 74917 3448
rect 11204 3408 11210 3420
rect 74905 3417 74917 3420
rect 74951 3417 74963 3451
rect 74905 3411 74963 3417
rect 74994 3408 75000 3460
rect 75052 3448 75058 3460
rect 75822 3448 75828 3460
rect 75052 3420 75828 3448
rect 75052 3408 75058 3420
rect 75822 3408 75828 3420
rect 75880 3408 75886 3460
rect 76190 3408 76196 3460
rect 76248 3448 76254 3460
rect 77110 3448 77116 3460
rect 76248 3420 77116 3448
rect 76248 3408 76254 3420
rect 77110 3408 77116 3420
rect 77168 3408 77174 3460
rect 77386 3408 77392 3460
rect 77444 3448 77450 3460
rect 78490 3448 78496 3460
rect 77444 3420 78496 3448
rect 77444 3408 77450 3420
rect 78490 3408 78496 3420
rect 78548 3408 78554 3460
rect 83274 3408 83280 3460
rect 83332 3448 83338 3460
rect 84102 3448 84108 3460
rect 83332 3420 84108 3448
rect 83332 3408 83338 3420
rect 84102 3408 84108 3420
rect 84160 3408 84166 3460
rect 85666 3408 85672 3460
rect 85724 3448 85730 3460
rect 89073 3451 89131 3457
rect 89073 3448 89085 3451
rect 85724 3420 89085 3448
rect 85724 3408 85730 3420
rect 89073 3417 89085 3420
rect 89119 3417 89131 3451
rect 89073 3411 89131 3417
rect 89162 3408 89168 3460
rect 89220 3448 89226 3460
rect 91480 3448 91508 3488
rect 132865 3485 132877 3488
rect 132911 3485 132923 3519
rect 132865 3479 132923 3485
rect 132954 3476 132960 3528
rect 133012 3516 133018 3528
rect 133782 3516 133788 3528
rect 133012 3488 133788 3516
rect 133012 3476 133018 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
rect 141234 3476 141240 3528
rect 141292 3516 141298 3528
rect 142062 3516 142068 3528
rect 141292 3488 142068 3516
rect 141292 3476 141298 3488
rect 142062 3476 142068 3488
rect 142120 3476 142126 3528
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 149057 3519 149115 3525
rect 149057 3485 149069 3519
rect 149103 3516 149115 3519
rect 173069 3519 173127 3525
rect 173069 3516 173081 3519
rect 149103 3488 173081 3516
rect 149103 3485 149115 3488
rect 149057 3479 149115 3485
rect 173069 3485 173081 3488
rect 173115 3485 173127 3519
rect 173069 3479 173127 3485
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173802 3516 173808 3528
rect 173216 3488 173808 3516
rect 173216 3476 173222 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 173897 3519 173955 3525
rect 173897 3485 173909 3519
rect 173943 3516 173955 3519
rect 173943 3488 174216 3516
rect 173943 3485 173955 3488
rect 173897 3479 173955 3485
rect 89220 3420 91508 3448
rect 91557 3451 91615 3457
rect 89220 3408 89226 3420
rect 91557 3417 91569 3451
rect 91603 3448 91615 3451
rect 123389 3451 123447 3457
rect 123389 3448 123401 3451
rect 91603 3420 123401 3448
rect 91603 3417 91615 3420
rect 91557 3411 91615 3417
rect 123389 3417 123401 3420
rect 123435 3417 123447 3451
rect 123389 3411 123447 3417
rect 123478 3408 123484 3460
rect 123536 3448 123542 3460
rect 124122 3448 124128 3460
rect 123536 3420 124128 3448
rect 123536 3408 123542 3420
rect 124122 3408 124128 3420
rect 124180 3408 124186 3460
rect 124674 3408 124680 3460
rect 124732 3448 124738 3460
rect 125318 3448 125324 3460
rect 124732 3420 125324 3448
rect 124732 3408 124738 3420
rect 125318 3408 125324 3420
rect 125376 3408 125382 3460
rect 125870 3408 125876 3460
rect 125928 3448 125934 3460
rect 126882 3448 126888 3460
rect 125928 3420 126888 3448
rect 125928 3408 125934 3420
rect 126882 3408 126888 3420
rect 126940 3408 126946 3460
rect 127066 3408 127072 3460
rect 127124 3448 127130 3460
rect 133874 3448 133880 3460
rect 127124 3420 133880 3448
rect 127124 3408 127130 3420
rect 133874 3408 133880 3420
rect 133932 3408 133938 3460
rect 138842 3408 138848 3460
rect 138900 3448 138906 3460
rect 174078 3448 174084 3460
rect 138900 3420 174084 3448
rect 138900 3408 138906 3420
rect 174078 3408 174084 3420
rect 174136 3408 174142 3460
rect 174188 3448 174216 3488
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177942 3516 177948 3528
rect 176712 3488 177948 3516
rect 176712 3476 176718 3488
rect 177942 3476 177948 3488
rect 178000 3476 178006 3528
rect 179506 3516 179512 3528
rect 178052 3488 179512 3516
rect 178052 3448 178080 3488
rect 179506 3476 179512 3488
rect 179564 3476 179570 3528
rect 183738 3476 183744 3528
rect 183796 3516 183802 3528
rect 184842 3516 184848 3528
rect 183796 3488 184848 3516
rect 183796 3476 183802 3488
rect 184842 3476 184848 3488
rect 184900 3476 184906 3528
rect 184934 3476 184940 3528
rect 184992 3516 184998 3528
rect 186958 3516 186964 3528
rect 184992 3488 186964 3516
rect 184992 3476 184998 3488
rect 186958 3476 186964 3488
rect 187016 3476 187022 3528
rect 187053 3519 187111 3525
rect 187053 3485 187065 3519
rect 187099 3516 187111 3519
rect 201328 3516 201356 3624
rect 208486 3612 208492 3624
rect 208544 3612 208550 3664
rect 277118 3612 277124 3664
rect 277176 3652 277182 3664
rect 280338 3652 280344 3664
rect 277176 3624 280344 3652
rect 277176 3612 277182 3624
rect 280338 3612 280344 3624
rect 280396 3612 280402 3664
rect 321462 3612 321468 3664
rect 321520 3652 321526 3664
rect 329190 3652 329196 3664
rect 321520 3624 329196 3652
rect 321520 3612 321526 3624
rect 329190 3612 329196 3624
rect 329248 3612 329254 3664
rect 331030 3612 331036 3664
rect 331088 3652 331094 3664
rect 342162 3652 342168 3664
rect 331088 3624 342168 3652
rect 331088 3612 331094 3624
rect 342162 3612 342168 3624
rect 342220 3612 342226 3664
rect 346302 3612 346308 3664
rect 346360 3652 346366 3664
rect 361114 3652 361120 3664
rect 346360 3624 361120 3652
rect 346360 3612 346366 3624
rect 361114 3612 361120 3624
rect 361172 3612 361178 3664
rect 362770 3612 362776 3664
rect 362828 3652 362834 3664
rect 383562 3652 383568 3664
rect 362828 3624 383568 3652
rect 362828 3612 362834 3624
rect 383562 3612 383568 3624
rect 383620 3612 383626 3664
rect 387702 3612 387708 3664
rect 387760 3652 387766 3664
rect 415486 3652 415492 3664
rect 387760 3624 415492 3652
rect 387760 3612 387766 3624
rect 415486 3612 415492 3624
rect 415544 3612 415550 3664
rect 416590 3612 416596 3664
rect 416648 3652 416654 3664
rect 417513 3655 417571 3661
rect 417513 3652 417525 3655
rect 416648 3624 417525 3652
rect 416648 3612 416654 3624
rect 417513 3621 417525 3624
rect 417559 3621 417571 3655
rect 417513 3615 417571 3621
rect 417605 3655 417663 3661
rect 417605 3621 417617 3655
rect 417651 3652 417663 3655
rect 419077 3655 419135 3661
rect 419077 3652 419089 3655
rect 417651 3624 419089 3652
rect 417651 3621 417663 3624
rect 417605 3615 417663 3621
rect 419077 3621 419089 3624
rect 419123 3621 419135 3655
rect 419077 3615 419135 3621
rect 419442 3612 419448 3664
rect 419500 3652 419506 3664
rect 421576 3652 421604 3692
rect 421653 3689 421665 3723
rect 421699 3720 421711 3723
rect 449802 3720 449808 3732
rect 421699 3692 449808 3720
rect 421699 3689 421711 3692
rect 421653 3683 421711 3689
rect 449802 3680 449808 3692
rect 449860 3680 449866 3732
rect 452562 3680 452568 3732
rect 452620 3720 452626 3732
rect 500586 3720 500592 3732
rect 452620 3692 500592 3720
rect 452620 3680 452626 3692
rect 500586 3680 500592 3692
rect 500644 3680 500650 3732
rect 507762 3680 507768 3732
rect 507820 3720 507826 3732
rect 571518 3720 571524 3732
rect 507820 3692 571524 3720
rect 507820 3680 507826 3692
rect 571518 3680 571524 3692
rect 571576 3680 571582 3732
rect 454494 3652 454500 3664
rect 419500 3624 421512 3652
rect 421576 3624 454500 3652
rect 419500 3612 419506 3624
rect 211154 3584 211160 3596
rect 205836 3556 211160 3584
rect 187099 3488 201356 3516
rect 187099 3485 187111 3488
rect 187053 3479 187111 3485
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 202782 3516 202788 3528
rect 201552 3488 202788 3516
rect 201552 3476 201558 3488
rect 202782 3476 202788 3488
rect 202840 3476 202846 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 205542 3516 205548 3528
rect 205140 3488 205548 3516
rect 205140 3476 205146 3488
rect 205542 3476 205548 3488
rect 205600 3476 205606 3528
rect 174188 3420 178080 3448
rect 179046 3408 179052 3460
rect 179104 3448 179110 3460
rect 205726 3448 205732 3460
rect 179104 3420 205732 3448
rect 179104 3408 179110 3420
rect 205726 3408 205732 3420
rect 205784 3408 205790 3460
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 39298 3380 39304 3392
rect 8812 3352 39304 3380
rect 8812 3340 8818 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 51350 3340 51356 3392
rect 51408 3380 51414 3392
rect 52362 3380 52368 3392
rect 51408 3352 52368 3380
rect 51408 3340 51414 3352
rect 52362 3340 52368 3352
rect 52420 3340 52426 3392
rect 52457 3383 52515 3389
rect 52457 3349 52469 3383
rect 52503 3380 52515 3383
rect 103606 3380 103612 3392
rect 52503 3352 103612 3380
rect 52503 3349 52515 3352
rect 52457 3343 52515 3349
rect 103606 3340 103612 3352
rect 103664 3340 103670 3392
rect 110506 3340 110512 3392
rect 110564 3380 110570 3392
rect 111702 3380 111708 3392
rect 110564 3352 111708 3380
rect 110564 3340 110570 3352
rect 111702 3340 111708 3352
rect 111760 3340 111766 3392
rect 112806 3340 112812 3392
rect 112864 3380 112870 3392
rect 154574 3380 154580 3392
rect 112864 3352 154580 3380
rect 112864 3340 112870 3352
rect 154574 3340 154580 3352
rect 154632 3340 154638 3392
rect 157794 3340 157800 3392
rect 157852 3380 157858 3392
rect 158622 3380 158628 3392
rect 157852 3352 158628 3380
rect 157852 3340 157858 3352
rect 158622 3340 158628 3352
rect 158680 3340 158686 3392
rect 158898 3340 158904 3392
rect 158956 3380 158962 3392
rect 160002 3380 160008 3392
rect 158956 3352 160008 3380
rect 158956 3340 158962 3352
rect 160002 3340 160008 3352
rect 160060 3340 160066 3392
rect 160094 3340 160100 3392
rect 160152 3380 160158 3392
rect 190546 3380 190552 3392
rect 160152 3352 190552 3380
rect 160152 3340 160158 3352
rect 190546 3340 190552 3352
rect 190604 3340 190610 3392
rect 190822 3340 190828 3392
rect 190880 3380 190886 3392
rect 191742 3380 191748 3392
rect 190880 3352 191748 3380
rect 190880 3340 190886 3352
rect 191742 3340 191748 3352
rect 191800 3340 191806 3392
rect 192018 3340 192024 3392
rect 192076 3380 192082 3392
rect 193122 3380 193128 3392
rect 192076 3352 193128 3380
rect 192076 3340 192082 3352
rect 193122 3340 193128 3352
rect 193180 3340 193186 3392
rect 194410 3340 194416 3392
rect 194468 3380 194474 3392
rect 195238 3380 195244 3392
rect 194468 3352 195244 3380
rect 194468 3340 194474 3352
rect 195238 3340 195244 3352
rect 195296 3340 195302 3392
rect 197906 3340 197912 3392
rect 197964 3380 197970 3392
rect 198642 3380 198648 3392
rect 197964 3352 198648 3380
rect 197964 3340 197970 3352
rect 198642 3340 198648 3352
rect 198700 3340 198706 3392
rect 199102 3340 199108 3392
rect 199160 3380 199166 3392
rect 200022 3380 200028 3392
rect 199160 3352 200028 3380
rect 199160 3340 199166 3352
rect 200022 3340 200028 3352
rect 200080 3340 200086 3392
rect 200117 3383 200175 3389
rect 200117 3349 200129 3383
rect 200163 3380 200175 3383
rect 205836 3380 205864 3556
rect 211154 3544 211160 3556
rect 211212 3544 211218 3596
rect 242158 3584 242164 3596
rect 238726 3556 242164 3584
rect 206186 3476 206192 3528
rect 206244 3516 206250 3528
rect 206922 3516 206928 3528
rect 206244 3488 206928 3516
rect 206244 3476 206250 3488
rect 206922 3476 206928 3488
rect 206980 3476 206986 3528
rect 208578 3476 208584 3528
rect 208636 3516 208642 3528
rect 209682 3516 209688 3528
rect 208636 3488 209688 3516
rect 208636 3476 208642 3488
rect 209682 3476 209688 3488
rect 209740 3476 209746 3528
rect 213362 3476 213368 3528
rect 213420 3516 213426 3528
rect 213822 3516 213828 3528
rect 213420 3488 213828 3516
rect 213420 3476 213426 3488
rect 213822 3476 213828 3488
rect 213880 3476 213886 3528
rect 214466 3476 214472 3528
rect 214524 3516 214530 3528
rect 215202 3516 215208 3528
rect 214524 3488 215208 3516
rect 214524 3476 214530 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 216582 3516 216588 3528
rect 215720 3488 216588 3516
rect 215720 3476 215726 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 219342 3516 219348 3528
rect 218112 3488 219348 3516
rect 218112 3476 218118 3488
rect 219342 3476 219348 3488
rect 219400 3476 219406 3528
rect 222746 3476 222752 3528
rect 222804 3516 222810 3528
rect 223482 3516 223488 3528
rect 222804 3488 223488 3516
rect 222804 3476 222810 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 224862 3516 224868 3528
rect 224000 3488 224868 3516
rect 224000 3476 224006 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 227622 3516 227628 3528
rect 226392 3488 227628 3516
rect 226392 3476 226398 3488
rect 227622 3476 227628 3488
rect 227680 3476 227686 3528
rect 231026 3476 231032 3528
rect 231084 3516 231090 3528
rect 231762 3516 231768 3528
rect 231084 3488 231768 3516
rect 231084 3476 231090 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 234614 3476 234620 3528
rect 234672 3516 234678 3528
rect 238726 3516 238754 3556
rect 242158 3544 242164 3556
rect 242216 3544 242222 3596
rect 247586 3544 247592 3596
rect 247644 3584 247650 3596
rect 249058 3584 249064 3596
rect 247644 3556 249064 3584
rect 247644 3544 247650 3556
rect 249058 3544 249064 3556
rect 249116 3544 249122 3596
rect 262950 3584 262956 3596
rect 258046 3556 262956 3584
rect 234672 3488 238754 3516
rect 234672 3476 234678 3488
rect 241698 3476 241704 3528
rect 241756 3516 241762 3528
rect 242802 3516 242808 3528
rect 241756 3488 242808 3516
rect 241756 3476 241762 3488
rect 242802 3476 242808 3488
rect 242860 3476 242866 3528
rect 244090 3476 244096 3528
rect 244148 3516 244154 3528
rect 244918 3516 244924 3528
rect 244148 3488 244924 3516
rect 244148 3476 244154 3488
rect 244918 3476 244924 3488
rect 244976 3476 244982 3528
rect 246390 3476 246396 3528
rect 246448 3516 246454 3528
rect 246942 3516 246948 3528
rect 246448 3488 246948 3516
rect 246448 3476 246454 3488
rect 246942 3476 246948 3488
rect 247000 3476 247006 3528
rect 248782 3476 248788 3528
rect 248840 3516 248846 3528
rect 250438 3516 250444 3528
rect 248840 3488 250444 3516
rect 248840 3476 248846 3488
rect 250438 3476 250444 3488
rect 250496 3476 250502 3528
rect 252370 3476 252376 3528
rect 252428 3516 252434 3528
rect 253198 3516 253204 3528
rect 252428 3488 253204 3516
rect 252428 3476 252434 3488
rect 253198 3476 253204 3488
rect 253256 3476 253262 3528
rect 254670 3476 254676 3528
rect 254728 3516 254734 3528
rect 255222 3516 255228 3528
rect 254728 3488 255228 3516
rect 254728 3476 254734 3488
rect 255222 3476 255228 3488
rect 255280 3476 255286 3528
rect 255866 3476 255872 3528
rect 255924 3516 255930 3528
rect 256602 3516 256608 3528
rect 255924 3488 256608 3516
rect 255924 3476 255930 3488
rect 256602 3476 256608 3488
rect 256660 3476 256666 3528
rect 257062 3476 257068 3528
rect 257120 3516 257126 3528
rect 258046 3516 258074 3556
rect 262950 3544 262956 3556
rect 263008 3544 263014 3596
rect 292574 3544 292580 3596
rect 292632 3584 292638 3596
rect 293678 3584 293684 3596
rect 292632 3556 293684 3584
rect 292632 3544 292638 3556
rect 293678 3544 293684 3556
rect 293736 3544 293742 3596
rect 314470 3544 314476 3596
rect 314528 3584 314534 3596
rect 319714 3584 319720 3596
rect 314528 3556 319720 3584
rect 314528 3544 314534 3556
rect 319714 3544 319720 3556
rect 319772 3544 319778 3596
rect 328270 3544 328276 3596
rect 328328 3584 328334 3596
rect 338666 3584 338672 3596
rect 328328 3556 338672 3584
rect 328328 3544 328334 3556
rect 338666 3544 338672 3556
rect 338724 3544 338730 3596
rect 343450 3544 343456 3596
rect 343508 3584 343514 3596
rect 358722 3584 358728 3596
rect 343508 3556 358728 3584
rect 343508 3544 343514 3556
rect 358722 3544 358728 3556
rect 358780 3544 358786 3596
rect 360010 3544 360016 3596
rect 360068 3584 360074 3596
rect 379974 3584 379980 3596
rect 360068 3556 379980 3584
rect 360068 3544 360074 3556
rect 379974 3544 379980 3556
rect 380032 3544 380038 3596
rect 386322 3544 386328 3596
rect 386380 3584 386386 3596
rect 414290 3584 414296 3596
rect 386380 3556 414296 3584
rect 386380 3544 386386 3556
rect 414290 3544 414296 3556
rect 414348 3544 414354 3596
rect 415302 3544 415308 3596
rect 415360 3584 415366 3596
rect 417145 3587 417203 3593
rect 417145 3584 417157 3587
rect 415360 3556 417157 3584
rect 415360 3544 415366 3556
rect 417145 3553 417157 3556
rect 417191 3553 417203 3587
rect 417145 3547 417203 3553
rect 417237 3587 417295 3593
rect 417237 3553 417249 3587
rect 417283 3584 417295 3587
rect 421374 3584 421380 3596
rect 417283 3556 421380 3584
rect 417283 3553 417295 3556
rect 417237 3547 417295 3553
rect 421374 3544 421380 3556
rect 421432 3544 421438 3596
rect 421484 3584 421512 3624
rect 454494 3612 454500 3624
rect 454552 3612 454558 3664
rect 458082 3612 458088 3664
rect 458140 3652 458146 3664
rect 507670 3652 507676 3664
rect 458140 3624 507676 3652
rect 458140 3612 458146 3624
rect 507670 3612 507676 3624
rect 507728 3612 507734 3664
rect 509142 3612 509148 3664
rect 509200 3652 509206 3664
rect 573910 3652 573916 3664
rect 509200 3624 573916 3652
rect 509200 3612 509206 3624
rect 573910 3612 573916 3624
rect 573968 3612 573974 3664
rect 427173 3587 427231 3593
rect 421484 3556 427124 3584
rect 257120 3488 258074 3516
rect 257120 3476 257126 3488
rect 261754 3476 261760 3528
rect 261812 3516 261818 3528
rect 262858 3516 262864 3528
rect 261812 3488 262864 3516
rect 261812 3476 261818 3488
rect 262858 3476 262864 3488
rect 262916 3476 262922 3528
rect 266538 3476 266544 3528
rect 266596 3516 266602 3528
rect 267642 3516 267648 3528
rect 266596 3488 267648 3516
rect 266596 3476 266602 3488
rect 267642 3476 267648 3488
rect 267700 3476 267706 3528
rect 267734 3476 267740 3528
rect 267792 3516 267798 3528
rect 269022 3516 269028 3528
rect 267792 3488 269028 3516
rect 267792 3476 267798 3488
rect 269022 3476 269028 3488
rect 269080 3476 269086 3528
rect 271230 3476 271236 3528
rect 271288 3516 271294 3528
rect 271782 3516 271788 3528
rect 271288 3488 271788 3516
rect 271288 3476 271294 3488
rect 271782 3476 271788 3488
rect 271840 3476 271846 3528
rect 276014 3476 276020 3528
rect 276072 3516 276078 3528
rect 277302 3516 277308 3528
rect 276072 3488 277308 3516
rect 276072 3476 276078 3488
rect 277302 3476 277308 3488
rect 277360 3476 277366 3528
rect 281902 3476 281908 3528
rect 281960 3516 281966 3528
rect 282822 3516 282828 3528
rect 281960 3488 282828 3516
rect 281960 3476 281966 3488
rect 282822 3476 282828 3488
rect 282880 3476 282886 3528
rect 283098 3476 283104 3528
rect 283156 3516 283162 3528
rect 284478 3516 284484 3528
rect 283156 3488 284484 3516
rect 283156 3476 283162 3488
rect 284478 3476 284484 3488
rect 284536 3476 284542 3528
rect 288986 3476 288992 3528
rect 289044 3516 289050 3528
rect 289722 3516 289728 3528
rect 289044 3488 289728 3516
rect 289044 3476 289050 3488
rect 289722 3476 289728 3488
rect 289780 3476 289786 3528
rect 293954 3476 293960 3528
rect 294012 3516 294018 3528
rect 294874 3516 294880 3528
rect 294012 3488 294880 3516
rect 294012 3476 294018 3488
rect 294874 3476 294880 3488
rect 294932 3476 294938 3528
rect 295334 3476 295340 3528
rect 295392 3516 295398 3528
rect 296070 3516 296076 3528
rect 295392 3488 296076 3516
rect 295392 3476 295398 3488
rect 296070 3476 296076 3488
rect 296128 3476 296134 3528
rect 300762 3476 300768 3528
rect 300820 3516 300826 3528
rect 301958 3516 301964 3528
rect 300820 3488 301964 3516
rect 300820 3476 300826 3488
rect 301958 3476 301964 3488
rect 302016 3476 302022 3528
rect 318150 3476 318156 3528
rect 318208 3516 318214 3528
rect 322106 3516 322112 3528
rect 318208 3488 322112 3516
rect 318208 3476 318214 3488
rect 322106 3476 322112 3488
rect 322164 3476 322170 3528
rect 325602 3476 325608 3528
rect 325660 3516 325666 3528
rect 335078 3516 335084 3528
rect 325660 3488 335084 3516
rect 325660 3476 325666 3488
rect 335078 3476 335084 3488
rect 335136 3476 335142 3528
rect 345750 3516 345756 3528
rect 335326 3488 345756 3516
rect 229830 3408 229836 3460
rect 229888 3448 229894 3460
rect 231118 3448 231124 3460
rect 229888 3420 231124 3448
rect 229888 3408 229894 3420
rect 231118 3408 231124 3420
rect 231176 3408 231182 3460
rect 238110 3408 238116 3460
rect 238168 3448 238174 3460
rect 238662 3448 238668 3460
rect 238168 3420 238668 3448
rect 238168 3408 238174 3420
rect 238662 3408 238668 3420
rect 238720 3408 238726 3460
rect 251174 3408 251180 3460
rect 251232 3448 251238 3460
rect 252462 3448 252468 3460
rect 251232 3420 252468 3448
rect 251232 3408 251238 3420
rect 252462 3408 252468 3420
rect 252520 3408 252526 3460
rect 259454 3408 259460 3460
rect 259512 3448 259518 3460
rect 264238 3448 264244 3460
rect 259512 3420 264244 3448
rect 259512 3408 259518 3420
rect 264238 3408 264244 3420
rect 264296 3408 264302 3460
rect 265342 3408 265348 3460
rect 265400 3448 265406 3460
rect 266998 3448 267004 3460
rect 265400 3420 267004 3448
rect 265400 3408 265406 3420
rect 266998 3408 267004 3420
rect 267056 3408 267062 3460
rect 306282 3408 306288 3460
rect 306340 3448 306346 3460
rect 309042 3448 309048 3460
rect 306340 3420 309048 3448
rect 306340 3408 306346 3420
rect 309042 3408 309048 3420
rect 309100 3408 309106 3460
rect 314562 3408 314568 3460
rect 314620 3448 314626 3460
rect 320910 3448 320916 3460
rect 314620 3420 320916 3448
rect 314620 3408 314626 3420
rect 320910 3408 320916 3420
rect 320968 3408 320974 3460
rect 322750 3408 322756 3460
rect 322808 3448 322814 3460
rect 331582 3448 331588 3460
rect 322808 3420 331588 3448
rect 322808 3408 322814 3420
rect 331582 3408 331588 3420
rect 331640 3408 331646 3460
rect 334618 3408 334624 3460
rect 334676 3448 334682 3460
rect 335326 3448 335354 3488
rect 345750 3476 345756 3488
rect 345808 3476 345814 3528
rect 346210 3476 346216 3528
rect 346268 3516 346274 3528
rect 362310 3516 362316 3528
rect 346268 3488 362316 3516
rect 346268 3476 346274 3488
rect 362310 3476 362316 3488
rect 362368 3476 362374 3528
rect 365530 3476 365536 3528
rect 365588 3516 365594 3528
rect 387150 3516 387156 3528
rect 365588 3488 387156 3516
rect 365588 3476 365594 3488
rect 387150 3476 387156 3488
rect 387208 3476 387214 3528
rect 389082 3476 389088 3528
rect 389140 3516 389146 3528
rect 417878 3516 417884 3528
rect 389140 3488 417884 3516
rect 389140 3476 389146 3488
rect 417878 3476 417884 3488
rect 417936 3476 417942 3528
rect 417973 3519 418031 3525
rect 417973 3485 417985 3519
rect 418019 3516 418031 3519
rect 421653 3519 421711 3525
rect 421653 3516 421665 3519
rect 418019 3488 421665 3516
rect 418019 3485 418031 3488
rect 417973 3479 418031 3485
rect 421653 3485 421665 3488
rect 421699 3485 421711 3519
rect 421653 3479 421711 3485
rect 422202 3476 422208 3528
rect 422260 3516 422266 3528
rect 427096 3516 427124 3556
rect 427173 3553 427185 3587
rect 427219 3584 427231 3587
rect 453298 3584 453304 3596
rect 427219 3556 453304 3584
rect 427219 3553 427231 3556
rect 427173 3547 427231 3553
rect 453298 3544 453304 3556
rect 453356 3544 453362 3596
rect 455322 3544 455328 3596
rect 455380 3584 455386 3596
rect 504174 3584 504180 3596
rect 455380 3556 504180 3584
rect 455380 3544 455386 3556
rect 504174 3544 504180 3556
rect 504232 3544 504238 3596
rect 506382 3544 506388 3596
rect 506440 3584 506446 3596
rect 570322 3584 570328 3596
rect 506440 3556 570328 3584
rect 506440 3544 506446 3556
rect 570322 3544 570328 3556
rect 570380 3544 570386 3596
rect 456886 3516 456892 3528
rect 422260 3488 427032 3516
rect 427096 3488 456892 3516
rect 422260 3476 422266 3488
rect 334676 3420 335354 3448
rect 334676 3408 334682 3420
rect 336550 3408 336556 3460
rect 336608 3448 336614 3460
rect 348050 3448 348056 3460
rect 336608 3420 348056 3448
rect 336608 3408 336614 3420
rect 348050 3408 348056 3420
rect 348108 3408 348114 3460
rect 349062 3408 349068 3460
rect 349120 3448 349126 3460
rect 365806 3448 365812 3460
rect 349120 3420 365812 3448
rect 349120 3408 349126 3420
rect 365806 3408 365812 3420
rect 365864 3408 365870 3460
rect 368290 3408 368296 3460
rect 368348 3448 368354 3460
rect 390646 3448 390652 3460
rect 368348 3420 390652 3448
rect 368348 3408 368354 3420
rect 390646 3408 390652 3420
rect 390704 3408 390710 3460
rect 391842 3408 391848 3460
rect 391900 3448 391906 3460
rect 417237 3451 417295 3457
rect 417237 3448 417249 3451
rect 391900 3420 417249 3448
rect 391900 3408 391906 3420
rect 417237 3417 417249 3420
rect 417283 3417 417295 3451
rect 417237 3411 417295 3417
rect 417329 3451 417387 3457
rect 417329 3417 417341 3451
rect 417375 3448 417387 3451
rect 424962 3448 424968 3460
rect 417375 3420 424968 3448
rect 417375 3417 417387 3420
rect 417329 3411 417387 3417
rect 424962 3408 424968 3420
rect 425020 3408 425026 3460
rect 425057 3451 425115 3457
rect 425057 3417 425069 3451
rect 425103 3448 425115 3451
rect 426253 3451 426311 3457
rect 426253 3448 426265 3451
rect 425103 3420 426265 3448
rect 425103 3417 425115 3420
rect 425057 3411 425115 3417
rect 426253 3417 426265 3420
rect 426299 3417 426311 3451
rect 427004 3448 427032 3488
rect 456886 3476 456892 3488
rect 456944 3476 456950 3528
rect 460842 3476 460848 3528
rect 460900 3516 460906 3528
rect 511258 3516 511264 3528
rect 460900 3488 511264 3516
rect 460900 3476 460906 3488
rect 511258 3476 511264 3488
rect 511316 3476 511322 3528
rect 511902 3476 511908 3528
rect 511960 3516 511966 3528
rect 577406 3516 577412 3528
rect 511960 3488 577412 3516
rect 511960 3476 511966 3488
rect 577406 3476 577412 3488
rect 577464 3476 577470 3528
rect 460382 3448 460388 3460
rect 427004 3420 460388 3448
rect 426253 3411 426311 3417
rect 460382 3408 460388 3420
rect 460440 3408 460446 3460
rect 463602 3408 463608 3460
rect 463660 3448 463666 3460
rect 514754 3448 514760 3460
rect 463660 3420 514760 3448
rect 463660 3408 463666 3420
rect 514754 3408 514760 3420
rect 514812 3408 514818 3460
rect 516042 3408 516048 3460
rect 516100 3448 516106 3460
rect 583386 3448 583392 3460
rect 516100 3420 583392 3448
rect 516100 3408 516106 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 200163 3352 205864 3380
rect 200163 3349 200175 3352
rect 200117 3343 200175 3349
rect 227530 3340 227536 3392
rect 227588 3380 227594 3392
rect 238018 3380 238024 3392
rect 227588 3352 238024 3380
rect 227588 3340 227594 3352
rect 238018 3340 238024 3352
rect 238076 3340 238082 3392
rect 279510 3340 279516 3392
rect 279568 3380 279574 3392
rect 280798 3380 280804 3392
rect 279568 3352 280804 3380
rect 279568 3340 279574 3352
rect 280798 3340 280804 3352
rect 280856 3340 280862 3392
rect 311802 3340 311808 3392
rect 311860 3380 311866 3392
rect 317322 3380 317328 3392
rect 311860 3352 317328 3380
rect 311860 3340 311866 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 318702 3340 318708 3392
rect 318760 3380 318766 3392
rect 325602 3380 325608 3392
rect 318760 3352 325608 3380
rect 318760 3340 318766 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 339310 3340 339316 3392
rect 339368 3380 339374 3392
rect 351638 3380 351644 3392
rect 339368 3352 351644 3380
rect 339368 3340 339374 3352
rect 351638 3340 351644 3352
rect 351696 3340 351702 3392
rect 353202 3340 353208 3392
rect 353260 3380 353266 3392
rect 370590 3380 370596 3392
rect 353260 3352 370596 3380
rect 353260 3340 353266 3352
rect 370590 3340 370596 3352
rect 370648 3340 370654 3392
rect 371050 3340 371056 3392
rect 371108 3380 371114 3392
rect 394234 3380 394240 3392
rect 371108 3352 394240 3380
rect 371108 3340 371114 3352
rect 394234 3340 394240 3352
rect 394292 3340 394298 3392
rect 397362 3340 397368 3392
rect 397420 3380 397426 3392
rect 428458 3380 428464 3392
rect 397420 3352 428464 3380
rect 397420 3340 397426 3352
rect 428458 3340 428464 3352
rect 428516 3340 428522 3392
rect 428553 3383 428611 3389
rect 428553 3349 428565 3383
rect 428599 3380 428611 3383
rect 436833 3383 436891 3389
rect 436833 3380 436845 3383
rect 428599 3352 436845 3380
rect 428599 3349 428611 3352
rect 428553 3343 428611 3349
rect 436833 3349 436845 3352
rect 436879 3349 436891 3383
rect 436833 3343 436891 3349
rect 436925 3383 436983 3389
rect 436925 3349 436937 3383
rect 436971 3380 436983 3383
rect 474550 3380 474556 3392
rect 436971 3352 474556 3380
rect 436971 3349 436983 3352
rect 436925 3343 436983 3349
rect 474550 3340 474556 3352
rect 474608 3340 474614 3392
rect 499482 3340 499488 3392
rect 499540 3380 499546 3392
rect 560846 3380 560852 3392
rect 499540 3352 560852 3380
rect 499540 3340 499546 3352
rect 560846 3340 560852 3352
rect 560904 3340 560910 3392
rect 28902 3272 28908 3324
rect 28960 3312 28966 3324
rect 35253 3315 35311 3321
rect 35253 3312 35265 3315
rect 28960 3284 35265 3312
rect 28960 3272 28966 3284
rect 35253 3281 35265 3284
rect 35299 3281 35311 3315
rect 35253 3275 35311 3281
rect 43070 3272 43076 3324
rect 43128 3312 43134 3324
rect 43128 3284 95648 3312
rect 43128 3272 43134 3284
rect 41874 3204 41880 3256
rect 41932 3244 41938 3256
rect 95421 3247 95479 3253
rect 95421 3244 95433 3247
rect 41932 3216 95433 3244
rect 41932 3204 41938 3216
rect 95421 3213 95433 3216
rect 95467 3213 95479 3247
rect 95421 3207 95479 3213
rect 566 3136 572 3188
rect 624 3176 630 3188
rect 3418 3176 3424 3188
rect 624 3148 3424 3176
rect 624 3136 630 3148
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 45462 3136 45468 3188
rect 45520 3176 45526 3188
rect 95513 3179 95571 3185
rect 95513 3176 95525 3179
rect 45520 3148 95525 3176
rect 45520 3136 45526 3148
rect 95513 3145 95525 3148
rect 95559 3145 95571 3179
rect 95620 3176 95648 3284
rect 96246 3272 96252 3324
rect 96304 3312 96310 3324
rect 102137 3315 102195 3321
rect 102137 3312 102149 3315
rect 96304 3284 102149 3312
rect 96304 3272 96310 3284
rect 102137 3281 102149 3284
rect 102183 3281 102195 3315
rect 102137 3275 102195 3281
rect 106918 3272 106924 3324
rect 106976 3312 106982 3324
rect 142341 3315 142399 3321
rect 142341 3312 142353 3315
rect 106976 3284 142353 3312
rect 106976 3272 106982 3284
rect 142341 3281 142353 3284
rect 142387 3281 142399 3315
rect 142341 3275 142399 3281
rect 142430 3272 142436 3324
rect 142488 3312 142494 3324
rect 149057 3315 149115 3321
rect 149057 3312 149069 3315
rect 142488 3284 149069 3312
rect 142488 3272 142494 3284
rect 149057 3281 149069 3284
rect 149103 3281 149115 3315
rect 149057 3275 149115 3281
rect 166074 3272 166080 3324
rect 166132 3312 166138 3324
rect 166902 3312 166908 3324
rect 166132 3284 166908 3312
rect 166132 3272 166138 3284
rect 166902 3272 166908 3284
rect 166960 3272 166966 3324
rect 171962 3272 171968 3324
rect 172020 3312 172026 3324
rect 200206 3312 200212 3324
rect 172020 3284 200212 3312
rect 172020 3272 172026 3284
rect 200206 3272 200212 3284
rect 200264 3272 200270 3324
rect 209774 3272 209780 3324
rect 209832 3312 209838 3324
rect 213178 3312 213184 3324
rect 209832 3284 213184 3312
rect 209832 3272 209838 3284
rect 213178 3272 213184 3284
rect 213236 3272 213242 3324
rect 262950 3272 262956 3324
rect 263008 3312 263014 3324
rect 269390 3312 269396 3324
rect 263008 3284 269396 3312
rect 263008 3272 263014 3284
rect 269390 3272 269396 3284
rect 269448 3272 269454 3324
rect 287790 3272 287796 3324
rect 287848 3312 287854 3324
rect 288342 3312 288348 3324
rect 287848 3284 288348 3312
rect 287848 3272 287854 3284
rect 288342 3272 288348 3284
rect 288400 3272 288406 3324
rect 310422 3272 310428 3324
rect 310480 3312 310486 3324
rect 315022 3312 315028 3324
rect 310480 3284 315028 3312
rect 310480 3272 310486 3284
rect 315022 3272 315028 3284
rect 315080 3272 315086 3324
rect 320818 3272 320824 3324
rect 320876 3312 320882 3324
rect 327994 3312 328000 3324
rect 320876 3284 328000 3312
rect 320876 3272 320882 3284
rect 327994 3272 328000 3284
rect 328052 3272 328058 3324
rect 335262 3272 335268 3324
rect 335320 3312 335326 3324
rect 346946 3312 346952 3324
rect 335320 3284 346952 3312
rect 335320 3272 335326 3284
rect 346946 3272 346952 3284
rect 347004 3272 347010 3324
rect 357342 3272 357348 3324
rect 357400 3312 357406 3324
rect 375282 3312 375288 3324
rect 357400 3284 375288 3312
rect 357400 3272 357406 3284
rect 375282 3272 375288 3284
rect 375340 3272 375346 3324
rect 376662 3272 376668 3324
rect 376720 3312 376726 3324
rect 401318 3312 401324 3324
rect 376720 3284 401324 3312
rect 376720 3272 376726 3284
rect 401318 3272 401324 3284
rect 401376 3272 401382 3324
rect 401502 3272 401508 3324
rect 401560 3312 401566 3324
rect 433242 3312 433248 3324
rect 401560 3284 433248 3312
rect 401560 3272 401566 3284
rect 433242 3272 433248 3284
rect 433300 3272 433306 3324
rect 434622 3272 434628 3324
rect 434680 3312 434686 3324
rect 436741 3315 436799 3321
rect 434680 3284 436600 3312
rect 434680 3272 434686 3284
rect 109310 3204 109316 3256
rect 109368 3244 109374 3256
rect 151998 3244 152004 3256
rect 109368 3216 152004 3244
rect 109368 3204 109374 3216
rect 151998 3204 152004 3216
rect 152056 3204 152062 3256
rect 154666 3244 154672 3256
rect 153212 3216 154672 3244
rect 100846 3176 100852 3188
rect 95620 3148 100852 3176
rect 95513 3139 95571 3145
rect 100846 3136 100852 3148
rect 100904 3136 100910 3188
rect 115198 3136 115204 3188
rect 115256 3176 115262 3188
rect 115842 3176 115848 3188
rect 115256 3148 115848 3176
rect 115256 3136 115262 3148
rect 115842 3136 115848 3148
rect 115900 3136 115906 3188
rect 116394 3136 116400 3188
rect 116452 3176 116458 3188
rect 117222 3176 117228 3188
rect 116452 3148 117228 3176
rect 116452 3136 116458 3148
rect 117222 3136 117228 3148
rect 117280 3136 117286 3188
rect 153212 3176 153240 3216
rect 154666 3204 154672 3216
rect 154724 3204 154730 3256
rect 168374 3204 168380 3256
rect 168432 3244 168438 3256
rect 197446 3244 197452 3256
rect 168432 3216 197452 3244
rect 168432 3204 168438 3216
rect 197446 3204 197452 3216
rect 197504 3204 197510 3256
rect 216858 3204 216864 3256
rect 216916 3244 216922 3256
rect 217962 3244 217968 3256
rect 216916 3216 217968 3244
rect 216916 3204 216922 3216
rect 217962 3204 217968 3216
rect 218020 3204 218026 3256
rect 258258 3204 258264 3256
rect 258316 3244 258322 3256
rect 259362 3244 259368 3256
rect 258316 3216 259368 3244
rect 258316 3204 258322 3216
rect 259362 3204 259368 3216
rect 259420 3204 259426 3256
rect 307662 3204 307668 3256
rect 307720 3244 307726 3256
rect 311434 3244 311440 3256
rect 307720 3216 311440 3244
rect 307720 3204 307726 3216
rect 311434 3204 311440 3216
rect 311492 3204 311498 3256
rect 317230 3204 317236 3256
rect 317288 3244 317294 3256
rect 323302 3244 323308 3256
rect 317288 3216 323308 3244
rect 317288 3204 317294 3216
rect 323302 3204 323308 3216
rect 323360 3204 323366 3256
rect 340138 3204 340144 3256
rect 340196 3244 340202 3256
rect 350442 3244 350448 3256
rect 340196 3216 350448 3244
rect 340196 3204 340202 3216
rect 350442 3204 350448 3216
rect 350500 3204 350506 3256
rect 351822 3204 351828 3256
rect 351880 3244 351886 3256
rect 369394 3244 369400 3256
rect 351880 3216 369400 3244
rect 351880 3204 351886 3216
rect 369394 3204 369400 3216
rect 369452 3204 369458 3256
rect 373902 3204 373908 3256
rect 373960 3244 373966 3256
rect 396534 3244 396540 3256
rect 373960 3216 396540 3244
rect 373960 3204 373966 3216
rect 396534 3204 396540 3216
rect 396592 3204 396598 3256
rect 404262 3204 404268 3256
rect 404320 3244 404326 3256
rect 407301 3247 407359 3253
rect 407301 3244 407313 3247
rect 404320 3216 407313 3244
rect 404320 3204 404326 3216
rect 407301 3213 407313 3216
rect 407347 3213 407359 3247
rect 407301 3207 407359 3213
rect 409782 3204 409788 3256
rect 409840 3244 409846 3256
rect 411993 3247 412051 3253
rect 411993 3244 412005 3247
rect 409840 3216 412005 3244
rect 409840 3204 409846 3216
rect 411993 3213 412005 3216
rect 412039 3213 412051 3247
rect 411993 3207 412051 3213
rect 412085 3247 412143 3253
rect 412085 3213 412097 3247
rect 412131 3244 412143 3247
rect 436462 3244 436468 3256
rect 412131 3216 436468 3244
rect 412131 3213 412143 3216
rect 412085 3207 412143 3213
rect 436462 3204 436468 3216
rect 436520 3204 436526 3256
rect 436572 3244 436600 3284
rect 436741 3281 436753 3315
rect 436787 3312 436799 3315
rect 471054 3312 471060 3324
rect 436787 3284 471060 3312
rect 436787 3281 436799 3284
rect 436741 3275 436799 3281
rect 471054 3272 471060 3284
rect 471112 3272 471118 3324
rect 496722 3272 496728 3324
rect 496780 3312 496786 3324
rect 557350 3312 557356 3324
rect 496780 3284 557356 3312
rect 496780 3272 496786 3284
rect 557350 3272 557356 3284
rect 557408 3272 557414 3324
rect 475746 3244 475752 3256
rect 436572 3216 475752 3244
rect 475746 3204 475752 3216
rect 475804 3204 475810 3256
rect 493962 3204 493968 3256
rect 494020 3244 494026 3256
rect 553762 3244 553768 3256
rect 494020 3216 553768 3244
rect 494020 3204 494026 3216
rect 553762 3204 553768 3216
rect 553820 3204 553826 3256
rect 117332 3148 153240 3176
rect 50154 3068 50160 3120
rect 50212 3108 50218 3120
rect 106274 3108 106280 3120
rect 50212 3080 106280 3108
rect 50212 3068 50218 3080
rect 106274 3068 106280 3080
rect 106332 3068 106338 3120
rect 114002 3068 114008 3120
rect 114060 3108 114066 3120
rect 117332 3108 117360 3148
rect 154206 3136 154212 3188
rect 154264 3176 154270 3188
rect 173066 3176 173072 3188
rect 154264 3148 173072 3176
rect 154264 3136 154270 3148
rect 173066 3136 173072 3148
rect 173124 3136 173130 3188
rect 175458 3136 175464 3188
rect 175516 3176 175522 3188
rect 202966 3176 202972 3188
rect 175516 3148 202972 3176
rect 175516 3136 175522 3148
rect 202966 3136 202972 3148
rect 203024 3136 203030 3188
rect 207382 3136 207388 3188
rect 207440 3176 207446 3188
rect 208302 3176 208308 3188
rect 207440 3148 208308 3176
rect 207440 3136 207446 3148
rect 208302 3136 208308 3148
rect 208360 3136 208366 3188
rect 239306 3136 239312 3188
rect 239364 3176 239370 3188
rect 246298 3176 246304 3188
rect 239364 3148 246304 3176
rect 239364 3136 239370 3148
rect 246298 3136 246304 3148
rect 246356 3136 246362 3188
rect 280706 3136 280712 3188
rect 280764 3176 280770 3188
rect 282178 3176 282184 3188
rect 280764 3148 282184 3176
rect 280764 3136 280770 3148
rect 282178 3136 282184 3148
rect 282236 3136 282242 3188
rect 311710 3136 311716 3188
rect 311768 3176 311774 3188
rect 316218 3176 316224 3188
rect 311768 3148 316224 3176
rect 311768 3136 311774 3148
rect 316218 3136 316224 3148
rect 316276 3136 316282 3188
rect 347682 3136 347688 3188
rect 347740 3176 347746 3188
rect 363506 3176 363512 3188
rect 347740 3148 363512 3176
rect 347740 3136 347746 3148
rect 363506 3136 363512 3148
rect 363564 3136 363570 3188
rect 371142 3136 371148 3188
rect 371200 3176 371206 3188
rect 393038 3176 393044 3188
rect 371200 3148 393044 3176
rect 371200 3136 371206 3148
rect 393038 3136 393044 3148
rect 393096 3136 393102 3188
rect 394602 3136 394608 3188
rect 394660 3176 394666 3188
rect 417329 3179 417387 3185
rect 417329 3176 417341 3179
rect 394660 3148 417341 3176
rect 394660 3136 394666 3148
rect 417329 3145 417341 3148
rect 417375 3145 417387 3179
rect 417329 3139 417387 3145
rect 417421 3179 417479 3185
rect 417421 3145 417433 3179
rect 417467 3176 417479 3179
rect 422570 3176 422576 3188
rect 417467 3148 422576 3176
rect 417467 3145 417479 3148
rect 417421 3139 417479 3145
rect 422570 3136 422576 3148
rect 422628 3136 422634 3188
rect 423582 3136 423588 3188
rect 423640 3176 423646 3188
rect 424781 3179 424839 3185
rect 424781 3176 424793 3179
rect 423640 3148 424793 3176
rect 423640 3136 423646 3148
rect 424781 3145 424793 3148
rect 424827 3145 424839 3179
rect 424781 3139 424839 3145
rect 424870 3136 424876 3188
rect 424928 3176 424934 3188
rect 427081 3179 427139 3185
rect 427081 3176 427093 3179
rect 424928 3148 427093 3176
rect 424928 3136 424934 3148
rect 427081 3145 427093 3148
rect 427127 3145 427139 3179
rect 427081 3139 427139 3145
rect 427722 3136 427728 3188
rect 427780 3176 427786 3188
rect 428553 3179 428611 3185
rect 428553 3176 428565 3179
rect 427780 3148 428565 3176
rect 427780 3136 427786 3148
rect 428553 3145 428565 3148
rect 428599 3145 428611 3179
rect 428553 3139 428611 3145
rect 428645 3179 428703 3185
rect 428645 3145 428657 3179
rect 428691 3176 428703 3179
rect 463970 3176 463976 3188
rect 428691 3148 463976 3176
rect 428691 3145 428703 3148
rect 428645 3139 428703 3145
rect 463970 3136 463976 3148
rect 464028 3136 464034 3188
rect 491202 3136 491208 3188
rect 491260 3176 491266 3188
rect 550266 3176 550272 3188
rect 491260 3148 550272 3176
rect 491260 3136 491266 3148
rect 550266 3136 550272 3148
rect 550324 3136 550330 3188
rect 114060 3080 117360 3108
rect 114060 3068 114066 3080
rect 117590 3068 117596 3120
rect 117648 3108 117654 3120
rect 125965 3111 126023 3117
rect 125965 3108 125977 3111
rect 117648 3080 125977 3108
rect 117648 3068 117654 3080
rect 125965 3077 125977 3080
rect 126011 3077 126023 3111
rect 125965 3071 126023 3077
rect 126054 3068 126060 3120
rect 126112 3108 126118 3120
rect 160186 3108 160192 3120
rect 126112 3080 160192 3108
rect 126112 3068 126118 3080
rect 160186 3068 160192 3080
rect 160244 3068 160250 3120
rect 167178 3068 167184 3120
rect 167236 3108 167242 3120
rect 180058 3108 180064 3120
rect 167236 3080 180064 3108
rect 167236 3068 167242 3080
rect 180058 3068 180064 3080
rect 180116 3068 180122 3120
rect 181438 3068 181444 3120
rect 181496 3108 181502 3120
rect 206278 3108 206284 3120
rect 181496 3080 206284 3108
rect 181496 3068 181502 3080
rect 206278 3068 206284 3080
rect 206336 3068 206342 3120
rect 221550 3068 221556 3120
rect 221608 3108 221614 3120
rect 222102 3108 222108 3120
rect 221608 3080 222108 3108
rect 221608 3068 221614 3080
rect 222102 3068 222108 3080
rect 222160 3068 222166 3120
rect 350350 3068 350356 3120
rect 350408 3108 350414 3120
rect 367002 3108 367008 3120
rect 350408 3080 367008 3108
rect 350408 3068 350414 3080
rect 367002 3068 367008 3080
rect 367060 3068 367066 3120
rect 368382 3068 368388 3120
rect 368440 3108 368446 3120
rect 389450 3108 389456 3120
rect 368440 3080 389456 3108
rect 368440 3068 368446 3080
rect 389450 3068 389456 3080
rect 389508 3068 389514 3120
rect 398742 3068 398748 3120
rect 398800 3108 398806 3120
rect 429654 3108 429660 3120
rect 398800 3080 429660 3108
rect 398800 3068 398806 3080
rect 429654 3068 429660 3080
rect 429712 3068 429718 3120
rect 430482 3068 430488 3120
rect 430540 3108 430546 3120
rect 436649 3111 436707 3117
rect 436649 3108 436661 3111
rect 430540 3080 436661 3108
rect 430540 3068 430546 3080
rect 436649 3077 436661 3080
rect 436695 3077 436707 3111
rect 468662 3108 468668 3120
rect 436649 3071 436707 3077
rect 436756 3080 468668 3108
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 11698 3040 11704 3052
rect 10008 3012 11704 3040
rect 10008 3000 10014 3012
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 22738 3040 22744 3052
rect 20680 3012 22744 3040
rect 20680 3000 20686 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 46658 3000 46664 3052
rect 46716 3040 46722 3052
rect 52457 3043 52515 3049
rect 52457 3040 52469 3043
rect 46716 3012 52469 3040
rect 46716 3000 46722 3012
rect 52457 3009 52469 3012
rect 52503 3009 52515 3043
rect 52457 3003 52515 3009
rect 53742 3000 53748 3052
rect 53800 3040 53806 3052
rect 109034 3040 109040 3052
rect 53800 3012 109040 3040
rect 53800 3000 53806 3012
rect 109034 3000 109040 3012
rect 109092 3000 109098 3052
rect 120258 3040 120264 3052
rect 114848 3012 120264 3040
rect 56042 2932 56048 2984
rect 56100 2972 56106 2984
rect 56502 2972 56508 2984
rect 56100 2944 56508 2972
rect 56100 2932 56106 2944
rect 56502 2932 56508 2944
rect 56560 2932 56566 2984
rect 57238 2932 57244 2984
rect 57296 2972 57302 2984
rect 57882 2972 57888 2984
rect 57296 2944 57888 2972
rect 57296 2932 57302 2944
rect 57882 2932 57888 2944
rect 57940 2932 57946 2984
rect 64322 2932 64328 2984
rect 64380 2972 64386 2984
rect 64782 2972 64788 2984
rect 64380 2944 64788 2972
rect 64380 2932 64386 2944
rect 64782 2932 64788 2944
rect 64840 2932 64846 2984
rect 65518 2932 65524 2984
rect 65576 2972 65582 2984
rect 66162 2972 66168 2984
rect 65576 2944 66168 2972
rect 65576 2932 65582 2944
rect 66162 2932 66168 2944
rect 66220 2932 66226 2984
rect 114738 2972 114744 2984
rect 68388 2944 114744 2972
rect 60826 2864 60832 2916
rect 60884 2904 60890 2916
rect 68388 2904 68416 2944
rect 114738 2932 114744 2944
rect 114796 2932 114802 2984
rect 114848 2904 114876 3012
rect 120258 3000 120264 3012
rect 120316 3000 120322 3052
rect 122282 3000 122288 3052
rect 122340 3040 122346 3052
rect 161566 3040 161572 3052
rect 122340 3012 161572 3040
rect 122340 3000 122346 3012
rect 161566 3000 161572 3012
rect 161624 3000 161630 3052
rect 177850 3000 177856 3052
rect 177908 3040 177914 3052
rect 184198 3040 184204 3052
rect 177908 3012 184204 3040
rect 177908 3000 177914 3012
rect 184198 3000 184204 3012
rect 184256 3000 184262 3052
rect 225138 3000 225144 3052
rect 225196 3040 225202 3052
rect 226978 3040 226984 3052
rect 225196 3012 226984 3040
rect 225196 3000 225202 3012
rect 226978 3000 226984 3012
rect 227036 3000 227042 3052
rect 240502 3000 240508 3052
rect 240560 3040 240566 3052
rect 241422 3040 241428 3052
rect 240560 3012 241428 3040
rect 240560 3000 240566 3012
rect 241422 3000 241428 3012
rect 241480 3000 241486 3052
rect 249978 3000 249984 3052
rect 250036 3040 250042 3052
rect 251818 3040 251824 3052
rect 250036 3012 251824 3040
rect 250036 3000 250042 3012
rect 251818 3000 251824 3012
rect 251876 3000 251882 3052
rect 272426 3000 272432 3052
rect 272484 3040 272490 3052
rect 273990 3040 273996 3052
rect 272484 3012 273996 3040
rect 272484 3000 272490 3012
rect 273990 3000 273996 3012
rect 274048 3000 274054 3052
rect 274818 3000 274824 3052
rect 274876 3040 274882 3052
rect 276658 3040 276664 3052
rect 274876 3012 276664 3040
rect 274876 3000 274882 3012
rect 276658 3000 276664 3012
rect 276716 3000 276722 3052
rect 322198 3000 322204 3052
rect 322256 3040 322262 3052
rect 326798 3040 326804 3052
rect 322256 3012 326804 3040
rect 322256 3000 322262 3012
rect 326798 3000 326804 3012
rect 326856 3000 326862 3052
rect 353938 3000 353944 3052
rect 353996 3040 354002 3052
rect 364610 3040 364616 3052
rect 353996 3012 364616 3040
rect 353996 3000 354002 3012
rect 364610 3000 364616 3012
rect 364668 3000 364674 3052
rect 366910 3000 366916 3052
rect 366968 3040 366974 3052
rect 388254 3040 388260 3052
rect 366968 3012 388260 3040
rect 366968 3000 366974 3012
rect 388254 3000 388260 3012
rect 388312 3000 388318 3052
rect 393222 3000 393228 3052
rect 393280 3040 393286 3052
rect 417421 3043 417479 3049
rect 417421 3040 417433 3043
rect 393280 3012 417433 3040
rect 393280 3000 393286 3012
rect 417421 3009 417433 3012
rect 417467 3009 417479 3043
rect 417421 3003 417479 3009
rect 417513 3043 417571 3049
rect 417513 3009 417525 3043
rect 417559 3040 417571 3043
rect 427173 3043 427231 3049
rect 427173 3040 427185 3043
rect 417559 3012 427185 3040
rect 417559 3009 417571 3012
rect 417513 3003 417571 3009
rect 427173 3009 427185 3012
rect 427219 3009 427231 3043
rect 427173 3003 427231 3009
rect 427265 3043 427323 3049
rect 427265 3009 427277 3043
rect 427311 3040 427323 3043
rect 428645 3043 428703 3049
rect 428645 3040 428657 3043
rect 427311 3012 428657 3040
rect 427311 3009 427323 3012
rect 427265 3003 427323 3009
rect 428645 3009 428657 3012
rect 428691 3009 428703 3043
rect 428645 3003 428703 3009
rect 429102 3000 429108 3052
rect 429160 3040 429166 3052
rect 436756 3040 436784 3080
rect 468662 3068 468668 3080
rect 468720 3068 468726 3120
rect 488442 3068 488448 3120
rect 488500 3108 488506 3120
rect 546678 3108 546684 3120
rect 488500 3080 546684 3108
rect 488500 3068 488506 3080
rect 546678 3068 546684 3080
rect 546736 3068 546742 3120
rect 429160 3012 436784 3040
rect 436833 3043 436891 3049
rect 429160 3000 429166 3012
rect 436833 3009 436845 3043
rect 436879 3040 436891 3043
rect 467466 3040 467472 3052
rect 436879 3012 467472 3040
rect 436879 3009 436891 3012
rect 436833 3003 436891 3009
rect 467466 3000 467472 3012
rect 467524 3000 467530 3052
rect 485682 3000 485688 3052
rect 485740 3040 485746 3052
rect 543182 3040 543188 3052
rect 485740 3012 543188 3040
rect 485740 3000 485746 3012
rect 543182 3000 543188 3012
rect 543240 3000 543246 3052
rect 119890 2932 119896 2984
rect 119948 2972 119954 2984
rect 126054 2972 126060 2984
rect 119948 2944 126060 2972
rect 119948 2932 119954 2944
rect 126054 2932 126060 2944
rect 126112 2932 126118 2984
rect 126149 2975 126207 2981
rect 126149 2941 126161 2975
rect 126195 2972 126207 2975
rect 157426 2972 157432 2984
rect 126195 2944 157432 2972
rect 126195 2941 126207 2944
rect 126149 2935 126207 2941
rect 157426 2932 157432 2944
rect 157484 2932 157490 2984
rect 172977 2975 173035 2981
rect 172977 2941 172989 2975
rect 173023 2972 173035 2975
rect 182266 2972 182272 2984
rect 173023 2944 182272 2972
rect 173023 2941 173035 2944
rect 172977 2935 173035 2941
rect 182266 2932 182272 2944
rect 182324 2932 182330 2984
rect 264146 2932 264152 2984
rect 264204 2972 264210 2984
rect 268378 2972 268384 2984
rect 264204 2944 268384 2972
rect 264204 2932 264210 2944
rect 268378 2932 268384 2944
rect 268436 2932 268442 2984
rect 365622 2932 365628 2984
rect 365680 2972 365686 2984
rect 385954 2972 385960 2984
rect 365680 2944 385960 2972
rect 365680 2932 365686 2944
rect 385954 2932 385960 2944
rect 386012 2932 386018 2984
rect 395982 2932 395988 2984
rect 396040 2972 396046 2984
rect 426158 2972 426164 2984
rect 396040 2944 426164 2972
rect 396040 2932 396046 2944
rect 426158 2932 426164 2944
rect 426216 2932 426222 2984
rect 426253 2975 426311 2981
rect 426253 2941 426265 2975
rect 426299 2972 426311 2975
rect 461578 2972 461584 2984
rect 426299 2944 461584 2972
rect 426299 2941 426311 2944
rect 426253 2935 426311 2941
rect 461578 2932 461584 2944
rect 461636 2932 461642 2984
rect 480162 2932 480168 2984
rect 480220 2972 480226 2984
rect 536098 2972 536104 2984
rect 480220 2944 536104 2972
rect 480220 2932 480226 2944
rect 536098 2932 536104 2944
rect 536156 2932 536162 2984
rect 118970 2904 118976 2916
rect 60884 2876 68416 2904
rect 68480 2876 114876 2904
rect 115860 2876 118976 2904
rect 60884 2864 60890 2876
rect 48958 2796 48964 2848
rect 49016 2836 49022 2848
rect 50890 2836 50896 2848
rect 49016 2808 50896 2836
rect 49016 2796 49022 2808
rect 50890 2796 50896 2808
rect 50948 2796 50954 2848
rect 66714 2796 66720 2848
rect 66772 2836 66778 2848
rect 66772 2808 67864 2836
rect 66772 2796 66778 2808
rect 67836 2768 67864 2808
rect 67910 2796 67916 2848
rect 67968 2836 67974 2848
rect 68480 2836 68508 2876
rect 115860 2836 115888 2876
rect 118970 2864 118976 2876
rect 119028 2864 119034 2916
rect 121086 2864 121092 2916
rect 121144 2904 121150 2916
rect 160462 2904 160468 2916
rect 121144 2876 160468 2904
rect 121144 2864 121150 2876
rect 160462 2864 160468 2876
rect 160520 2864 160526 2916
rect 268838 2864 268844 2916
rect 268896 2904 268902 2916
rect 273898 2904 273904 2916
rect 268896 2876 273904 2904
rect 268896 2864 268902 2876
rect 273898 2864 273904 2876
rect 273956 2864 273962 2916
rect 284294 2864 284300 2916
rect 284352 2904 284358 2916
rect 285674 2904 285680 2916
rect 284352 2876 285680 2904
rect 284352 2864 284358 2876
rect 285674 2864 285680 2876
rect 285732 2864 285738 2916
rect 335998 2864 336004 2916
rect 336056 2904 336062 2916
rect 344554 2904 344560 2916
rect 336056 2876 344560 2904
rect 336056 2864 336062 2876
rect 344554 2864 344560 2876
rect 344612 2864 344618 2916
rect 364242 2864 364248 2916
rect 364300 2904 364306 2916
rect 384758 2904 384764 2916
rect 364300 2876 384764 2904
rect 364300 2864 364306 2876
rect 384758 2864 384764 2876
rect 384816 2864 384822 2916
rect 390462 2864 390468 2916
rect 390520 2904 390526 2916
rect 418982 2904 418988 2916
rect 390520 2876 418988 2904
rect 390520 2864 390526 2876
rect 418982 2864 418988 2876
rect 419040 2864 419046 2916
rect 419077 2907 419135 2913
rect 419077 2873 419089 2907
rect 419123 2904 419135 2907
rect 450906 2904 450912 2916
rect 419123 2876 450912 2904
rect 419123 2873 419135 2876
rect 419077 2867 419135 2873
rect 450906 2864 450912 2876
rect 450964 2864 450970 2916
rect 474642 2864 474648 2916
rect 474700 2904 474706 2916
rect 529014 2904 529020 2916
rect 474700 2876 529020 2904
rect 474700 2864 474706 2876
rect 529014 2864 529020 2876
rect 529072 2864 529078 2916
rect 67968 2808 68508 2836
rect 68572 2808 115888 2836
rect 67968 2796 67974 2808
rect 68572 2768 68600 2808
rect 118786 2796 118792 2848
rect 118844 2836 118850 2848
rect 158806 2836 158812 2848
rect 118844 2808 158812 2836
rect 118844 2796 118850 2808
rect 158806 2796 158812 2808
rect 158864 2796 158870 2848
rect 359458 2796 359464 2848
rect 359516 2836 359522 2848
rect 368198 2836 368204 2848
rect 359516 2808 368204 2836
rect 359516 2796 359522 2808
rect 368198 2796 368204 2808
rect 368256 2796 368262 2848
rect 384942 2796 384948 2848
rect 385000 2836 385006 2848
rect 411898 2836 411904 2848
rect 385000 2808 411904 2836
rect 385000 2796 385006 2808
rect 411898 2796 411904 2808
rect 411956 2796 411962 2848
rect 411993 2839 412051 2845
rect 411993 2805 412005 2839
rect 412039 2836 412051 2839
rect 443822 2836 443828 2848
rect 412039 2808 443828 2836
rect 412039 2805 412051 2808
rect 411993 2799 412051 2805
rect 443822 2796 443828 2808
rect 443880 2796 443886 2848
rect 469122 2796 469128 2848
rect 469180 2836 469186 2848
rect 521838 2836 521844 2848
rect 469180 2808 521844 2836
rect 469180 2796 469186 2808
rect 521838 2796 521844 2808
rect 521896 2796 521902 2848
rect 67836 2740 68600 2768
<< via1 >>
rect 154120 700952 154172 701004
rect 324320 700952 324372 701004
rect 137836 700884 137888 700936
rect 320180 700884 320232 700936
rect 263508 700816 263560 700868
rect 462320 700816 462372 700868
rect 267648 700748 267700 700800
rect 478512 700748 478564 700800
rect 89168 700680 89220 700732
rect 336740 700680 336792 700732
rect 72976 700612 73028 700664
rect 332600 700612 332652 700664
rect 251088 700544 251140 700596
rect 527180 700544 527232 700596
rect 255228 700476 255280 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 340880 700408 340932 700460
rect 24308 700340 24360 700392
rect 347780 700340 347832 700392
rect 8116 700272 8168 700324
rect 343640 700272 343692 700324
rect 278688 700204 278740 700256
rect 413652 700204 413704 700256
rect 274548 700136 274600 700188
rect 397460 700136 397512 700188
rect 202788 700068 202840 700120
rect 309140 700068 309192 700120
rect 218980 700000 219032 700052
rect 313280 700000 313332 700052
rect 291108 699932 291160 699984
rect 348792 699932 348844 699984
rect 286968 699864 287020 699916
rect 332508 699864 332560 699916
rect 267556 699796 267608 699848
rect 296720 699796 296772 699848
rect 283840 699728 283892 699780
rect 300860 699728 300912 699780
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 240048 696940 240100 696992
rect 580172 696940 580224 696992
rect 244188 683204 244240 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 351920 683136 351972 683188
rect 235816 670760 235868 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 360200 670692 360252 670744
rect 3424 656888 3476 656940
rect 356060 656888 356112 656940
rect 227628 643084 227680 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 364432 632068 364484 632120
rect 231768 630640 231820 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 371240 618264 371292 618316
rect 223488 616836 223540 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 367100 605820 367152 605872
rect 216588 590656 216640 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 375840 579640 375892 579692
rect 4804 578280 4856 578332
rect 430856 578280 430908 578332
rect 14464 578212 14516 578264
rect 442632 578212 442684 578264
rect 215760 578144 215812 578196
rect 216588 578144 216640 578196
rect 235356 578144 235408 578196
rect 235816 578144 235868 578196
rect 239312 578144 239364 578196
rect 240048 578144 240100 578196
rect 243268 578144 243320 578196
rect 244188 578144 244240 578196
rect 262864 578144 262916 578196
rect 263508 578144 263560 578196
rect 266820 578144 266872 578196
rect 267648 578144 267700 578196
rect 282460 578144 282512 578196
rect 235908 578076 235960 578128
rect 286416 578008 286468 578060
rect 286968 578008 287020 578060
rect 290280 578144 290332 578196
rect 291108 578144 291160 578196
rect 293868 578144 293920 578196
rect 299480 578144 299532 578196
rect 305368 578076 305420 578128
rect 364340 578008 364392 578060
rect 171048 577940 171100 577992
rect 317420 577940 317472 577992
rect 270408 577872 270460 577924
rect 429200 577872 429252 577924
rect 106188 577804 106240 577856
rect 328920 577804 328972 577856
rect 258908 577736 258960 577788
rect 494060 577736 494112 577788
rect 246948 577668 247000 577720
rect 558920 577668 558972 577720
rect 53104 577600 53156 577652
rect 407396 577600 407448 577652
rect 184388 577532 184440 577584
rect 538864 577532 538916 577584
rect 219348 577464 219400 577516
rect 580172 577464 580224 577516
rect 172428 577396 172480 577448
rect 537484 577396 537536 577448
rect 160836 577328 160888 577380
rect 536104 577328 536156 577380
rect 168748 577260 168800 577312
rect 551284 577260 551336 577312
rect 148968 577192 149020 577244
rect 533344 577192 533396 577244
rect 137284 577124 137336 577176
rect 530584 577124 530636 577176
rect 125324 577056 125376 577108
rect 529204 577056 529256 577108
rect 121368 576988 121420 577040
rect 543004 576988 543056 577040
rect 17224 576920 17276 576972
rect 454408 576920 454460 576972
rect 18604 576852 18656 576904
rect 466460 576852 466512 576904
rect 211896 576716 211948 576768
rect 519544 576716 519596 576768
rect 199936 576648 199988 576700
rect 518164 576648 518216 576700
rect 188344 576580 188396 576632
rect 516784 576580 516836 576632
rect 66904 576512 66956 576564
rect 423036 576512 423088 576564
rect 36544 576444 36596 576496
rect 399484 576444 399536 576496
rect 57244 576376 57296 576428
rect 426992 576376 427044 576428
rect 153016 576308 153068 576360
rect 525064 576308 525116 576360
rect 61384 576240 61436 576292
rect 434812 576240 434864 576292
rect 11704 576172 11756 576224
rect 387800 576172 387852 576224
rect 39304 576104 39356 576156
rect 419080 576104 419132 576156
rect 65524 576036 65576 576088
rect 446588 576036 446640 576088
rect 141240 575968 141292 576020
rect 522304 575968 522356 576020
rect 25504 575900 25556 575952
rect 411260 575900 411312 575952
rect 156972 575832 157024 575884
rect 548524 575832 548576 575884
rect 129464 575764 129516 575816
rect 520924 575764 520976 575816
rect 47584 575696 47636 575748
rect 458686 575696 458738 575748
rect 133420 575628 133472 575680
rect 544384 575628 544436 575680
rect 51724 575560 51776 575612
rect 470140 575560 470192 575612
rect 50344 575492 50396 575544
rect 474004 575492 474056 575544
rect 54484 575288 54536 575340
rect 395620 575288 395672 575340
rect 207940 575220 207992 575272
rect 580816 575220 580868 575272
rect 3884 575152 3936 575204
rect 379888 575152 379940 575204
rect 203984 575084 204036 575136
rect 580908 575084 580960 575136
rect 3976 575016 4028 575068
rect 383844 575016 383896 575068
rect 391848 575059 391900 575068
rect 391848 575025 391857 575059
rect 391857 575025 391891 575059
rect 391891 575025 391900 575059
rect 391848 575016 391900 575025
rect 403440 575059 403492 575068
rect 403440 575025 403449 575059
rect 403449 575025 403483 575059
rect 403483 575025 403492 575059
rect 403440 575016 403492 575025
rect 415400 575059 415452 575068
rect 415400 575025 415409 575059
rect 415409 575025 415443 575059
rect 415443 575025 415452 575059
rect 415400 575016 415452 575025
rect 438860 575059 438912 575068
rect 438860 575025 438869 575059
rect 438869 575025 438903 575059
rect 438903 575025 438912 575059
rect 438860 575016 438912 575025
rect 450544 575059 450596 575068
rect 450544 575025 450553 575059
rect 450553 575025 450587 575059
rect 450587 575025 450596 575059
rect 450544 575016 450596 575025
rect 462320 575059 462372 575068
rect 462320 575025 462329 575059
rect 462329 575025 462363 575059
rect 462363 575025 462372 575059
rect 462320 575016 462372 575025
rect 195980 574948 196032 575000
rect 580632 574948 580684 575000
rect 109868 574923 109920 574932
rect 109868 574889 109877 574923
rect 109877 574889 109911 574923
rect 109911 574889 109920 574923
rect 109868 574880 109920 574889
rect 117688 574923 117740 574932
rect 117688 574889 117697 574923
rect 117697 574889 117731 574923
rect 117731 574889 117740 574923
rect 117688 574880 117740 574889
rect 145012 574923 145064 574932
rect 145012 574889 145021 574923
rect 145021 574889 145055 574923
rect 145055 574889 145064 574923
rect 145012 574880 145064 574889
rect 164792 574923 164844 574932
rect 164792 574889 164801 574923
rect 164801 574889 164835 574923
rect 164835 574889 164844 574923
rect 164792 574880 164844 574889
rect 176568 574923 176620 574932
rect 176568 574889 176577 574923
rect 176577 574889 176611 574923
rect 176611 574889 176620 574923
rect 176568 574880 176620 574889
rect 180432 574923 180484 574932
rect 180432 574889 180441 574923
rect 180441 574889 180475 574923
rect 180475 574889 180484 574923
rect 180432 574880 180484 574889
rect 192208 574880 192260 574932
rect 580724 574880 580776 574932
rect 3792 574812 3844 574864
rect 58624 574744 58676 574796
rect 3700 574676 3752 574728
rect 580540 574608 580592 574660
rect 547144 574540 547196 574592
rect 580448 574472 580500 574524
rect 3608 574404 3660 574456
rect 580356 574336 580408 574388
rect 540244 574268 540296 574320
rect 3516 574200 3568 574252
rect 3424 574132 3476 574184
rect 580264 574064 580316 574116
rect 519544 564340 519596 564392
rect 580172 564340 580224 564392
rect 3240 528504 3292 528556
rect 11704 528504 11756 528556
rect 3332 516060 3384 516112
rect 54484 516060 54536 516112
rect 518164 511912 518216 511964
rect 580172 511912 580224 511964
rect 3332 476008 3384 476060
rect 36544 476008 36596 476060
rect 3332 463632 3384 463684
rect 53104 463632 53156 463684
rect 516784 458124 516836 458176
rect 580172 458124 580224 458176
rect 3332 423580 3384 423632
rect 25504 423580 25556 423632
rect 538864 419432 538916 419484
rect 579712 419432 579764 419484
rect 3332 411204 3384 411256
rect 39304 411204 39356 411256
rect 551284 379448 551336 379500
rect 580172 379448 580224 379500
rect 3332 372512 3384 372564
rect 66904 372512 66956 372564
rect 537484 365644 537536 365696
rect 579988 365644 580040 365696
rect 2780 358436 2832 358488
rect 4804 358436 4856 358488
rect 3332 346332 3384 346384
rect 57244 346332 57296 346384
rect 548524 325592 548576 325644
rect 579896 325592 579948 325644
rect 3332 320084 3384 320136
rect 61384 320084 61436 320136
rect 536104 313216 536156 313268
rect 580172 313216 580224 313268
rect 3332 306280 3384 306332
rect 14464 306280 14516 306332
rect 525064 299412 525116 299464
rect 579620 299412 579672 299464
rect 547144 273164 547196 273216
rect 579896 273164 579948 273216
rect 3516 267656 3568 267708
rect 65524 267656 65576 267708
rect 533344 259360 533396 259412
rect 579804 259360 579856 259412
rect 3148 255212 3200 255264
rect 17224 255212 17276 255264
rect 522304 245556 522356 245608
rect 580172 245556 580224 245608
rect 3516 241408 3568 241460
rect 58624 241408 58676 241460
rect 544384 233180 544436 233232
rect 580172 233180 580224 233232
rect 530584 219376 530636 219428
rect 579896 219376 579948 219428
rect 3332 215228 3384 215280
rect 47584 215228 47636 215280
rect 520924 206932 520976 206984
rect 580172 206932 580224 206984
rect 3056 202784 3108 202836
rect 18604 202784 18656 202836
rect 543004 193128 543056 193180
rect 580172 193128 580224 193180
rect 529204 179324 529256 179376
rect 579988 179324 580040 179376
rect 3240 164160 3292 164212
rect 51724 164160 51776 164212
rect 540244 153144 540296 153196
rect 580172 153144 580224 153196
rect 3424 150356 3476 150408
rect 21364 150356 21416 150408
rect 526444 139340 526496 139392
rect 580172 139340 580224 139392
rect 3240 137912 3292 137964
rect 50344 137912 50396 137964
rect 93860 128188 93912 128240
rect 95010 128188 95062 128240
rect 125692 128188 125744 128240
rect 126842 128188 126894 128240
rect 146300 128188 146352 128240
rect 147634 128188 147686 128240
rect 149060 128188 149112 128240
rect 150394 128188 150446 128240
rect 157432 128188 157484 128240
rect 158582 128188 158634 128240
rect 186412 128188 186464 128240
rect 187562 128188 187614 128240
rect 212632 128188 212684 128240
rect 213874 128188 213926 128240
rect 215392 128188 215444 128240
rect 216634 128188 216686 128240
rect 218152 128188 218204 128240
rect 219302 128188 219354 128240
rect 220912 128188 220964 128240
rect 222062 128188 222114 128240
rect 287152 128188 287204 128240
rect 288302 128188 288354 128240
rect 64788 126896 64840 126948
rect 117688 126896 117740 126948
rect 122104 126896 122156 126948
rect 124036 126896 124088 126948
rect 125508 126896 125560 126948
rect 163964 126896 164016 126948
rect 170404 126896 170456 126948
rect 172152 126896 172204 126948
rect 199292 126896 199344 126948
rect 200028 126896 200080 126948
rect 221096 126896 221148 126948
rect 223488 126896 223540 126948
rect 239220 126896 239272 126948
rect 276664 126896 276716 126948
rect 279148 126896 279200 126948
rect 344560 126896 344612 126948
rect 345664 126896 345716 126948
rect 401692 126896 401744 126948
rect 403624 126896 403676 126948
rect 472440 126896 472492 126948
rect 56508 126828 56560 126880
rect 111340 126828 111392 126880
rect 112536 126828 112588 126880
rect 113180 126828 113232 126880
rect 126244 126828 126296 126880
rect 145840 126828 145892 126880
rect 160008 126828 160060 126880
rect 190276 126828 190328 126880
rect 195244 126828 195296 126880
rect 217508 126828 217560 126880
rect 220084 126828 220136 126880
rect 236552 126828 236604 126880
rect 238024 126828 238076 126880
rect 242900 126828 242952 126880
rect 246304 126828 246356 126880
rect 251916 126828 251968 126880
rect 312820 126828 312872 126880
rect 317420 126828 317472 126880
rect 469772 126828 469824 126880
rect 519544 126828 519596 126880
rect 57888 126760 57940 126812
rect 112260 126760 112312 126812
rect 112444 126760 112496 126812
rect 121276 126760 121328 126812
rect 124128 126760 124180 126812
rect 163044 126760 163096 126812
rect 171048 126760 171100 126812
rect 198372 126760 198424 126812
rect 202696 126760 202748 126812
rect 223856 126760 223908 126812
rect 224868 126760 224920 126812
rect 240140 126760 240192 126812
rect 242808 126760 242860 126812
rect 253756 126760 253808 126812
rect 256608 126760 256660 126812
rect 264612 126760 264664 126812
rect 285588 126760 285640 126812
rect 287336 126760 287388 126812
rect 440700 126760 440752 126812
rect 450544 126760 450596 126812
rect 466092 126760 466144 126812
rect 517520 126760 517572 126812
rect 29644 126692 29696 126744
rect 89536 126692 89588 126744
rect 117228 126692 117280 126744
rect 157616 126692 157668 126744
rect 162768 126692 162820 126744
rect 192944 126692 192996 126744
rect 193128 126692 193180 126744
rect 215668 126692 215720 126744
rect 216588 126692 216640 126744
rect 233792 126692 233844 126744
rect 238668 126692 238720 126744
rect 250996 126692 251048 126744
rect 253204 126692 253256 126744
rect 261944 126692 261996 126744
rect 448888 126692 448940 126744
rect 14464 126624 14516 126676
rect 73252 126624 73304 126676
rect 78496 126624 78548 126676
rect 127624 126624 127676 126676
rect 152556 126624 152608 126676
rect 153936 126624 153988 126676
rect 158628 126624 158680 126676
rect 189356 126624 189408 126676
rect 191748 126624 191800 126676
rect 214748 126624 214800 126676
rect 217968 126624 218020 126676
rect 234712 126624 234764 126676
rect 235908 126624 235960 126676
rect 249248 126624 249300 126676
rect 250444 126624 250496 126676
rect 259184 126624 259236 126676
rect 415308 126624 415360 126676
rect 442264 126624 442316 126676
rect 457076 126624 457128 126676
rect 464344 126624 464396 126676
rect 22744 126556 22796 126608
rect 84108 126556 84160 126608
rect 111708 126556 111760 126608
rect 153016 126556 153068 126608
rect 153108 126556 153160 126608
rect 185676 126556 185728 126608
rect 188988 126556 189040 126608
rect 212908 126556 212960 126608
rect 213828 126556 213880 126608
rect 231952 126556 232004 126608
rect 237288 126556 237340 126608
rect 250168 126556 250220 126608
rect 252468 126556 252520 126608
rect 261024 126556 261076 126608
rect 420736 126556 420788 126608
rect 432604 126556 432656 126608
rect 437112 126556 437164 126608
rect 471336 126556 471388 126608
rect 477040 126692 477092 126744
rect 536104 126692 536156 126744
rect 471520 126624 471572 126676
rect 524420 126624 524472 126676
rect 479524 126556 479576 126608
rect 531320 126556 531372 126608
rect 25504 126488 25556 126540
rect 86868 126488 86920 126540
rect 88248 126488 88300 126540
rect 99564 126488 99616 126540
rect 104808 126488 104860 126540
rect 148508 126488 148560 126540
rect 148968 126488 149020 126540
rect 182088 126488 182140 126540
rect 187608 126488 187660 126540
rect 21364 126420 21416 126472
rect 82268 126420 82320 126472
rect 88984 126420 89036 126472
rect 96620 126420 96672 126472
rect 99288 126420 99340 126472
rect 144000 126420 144052 126472
rect 144828 126420 144880 126472
rect 179328 126420 179380 126472
rect 184756 126420 184808 126472
rect 209320 126420 209372 126472
rect 17224 126352 17276 126404
rect 79600 126352 79652 126404
rect 93768 126352 93820 126404
rect 139492 126352 139544 126404
rect 142068 126352 142120 126404
rect 176660 126352 176712 126404
rect 177948 126352 178000 126404
rect 203892 126352 203944 126404
rect 212448 126488 212500 126540
rect 231032 126488 231084 126540
rect 234528 126488 234580 126540
rect 247408 126488 247460 126540
rect 249064 126488 249116 126540
rect 258264 126488 258316 126540
rect 267648 126488 267700 126540
rect 272800 126488 272852 126540
rect 399024 126488 399076 126540
rect 418804 126488 418856 126540
rect 419816 126488 419868 126540
rect 456892 126488 456944 126540
rect 459744 126488 459796 126540
rect 471244 126488 471296 126540
rect 478788 126488 478840 126540
rect 533344 126488 533396 126540
rect 209688 126420 209740 126472
rect 228364 126420 228416 126472
rect 231124 126420 231176 126472
rect 244648 126420 244700 126472
rect 246948 126420 247000 126472
rect 257344 126420 257396 126472
rect 409788 126420 409840 126472
rect 429752 126420 429804 126472
rect 434352 126420 434404 126472
rect 484216 126420 484268 126472
rect 547144 126420 547196 126472
rect 211988 126352 212040 126404
rect 225604 126352 225656 126404
rect 229008 126352 229060 126404
rect 243728 126352 243780 126404
rect 245568 126352 245620 126404
rect 256516 126352 256568 126404
rect 260748 126352 260800 126404
rect 268292 126352 268344 126404
rect 332784 126352 332836 126404
rect 336004 126352 336056 126404
rect 388076 126352 388128 126404
rect 407764 126352 407816 126404
rect 428924 126352 428976 126404
rect 467104 126352 467156 126404
rect 486976 126352 487028 126404
rect 543004 126352 543056 126404
rect 7564 126284 7616 126336
rect 72332 126284 72384 126336
rect 75828 126284 75880 126336
rect 125876 126284 125928 126336
rect 130384 126284 130436 126336
rect 165620 126284 165672 126336
rect 166908 126284 166960 126336
rect 195704 126284 195756 126336
rect 195888 126284 195940 126336
rect 218336 126284 218388 126336
rect 220728 126284 220780 126336
rect 237380 126284 237432 126336
rect 241428 126284 241480 126336
rect 252836 126284 252888 126336
rect 255228 126284 255280 126336
rect 263692 126284 263744 126336
rect 350908 126284 350960 126336
rect 359464 126284 359516 126336
rect 377220 126284 377272 126336
rect 389824 126284 389876 126336
rect 393504 126284 393556 126336
rect 421564 126284 421616 126336
rect 423496 126284 423548 126336
rect 461492 126284 461544 126336
rect 470508 126284 470560 126336
rect 475384 126284 475436 126336
rect 482468 126284 482520 126336
rect 539600 126284 539652 126336
rect 11704 126216 11756 126268
rect 75920 126216 75972 126268
rect 78588 126216 78640 126268
rect 128360 126216 128412 126268
rect 137928 126216 137980 126268
rect 173900 126216 173952 126268
rect 180708 126216 180760 126268
rect 206560 126216 206612 126268
rect 206928 126216 206980 126268
rect 226524 126216 226576 126268
rect 227628 126216 227680 126268
rect 241980 126216 242032 126268
rect 244924 126216 244976 126268
rect 255596 126216 255648 126268
rect 267004 126216 267056 126268
rect 271880 126216 271932 126268
rect 273996 126216 274048 126268
rect 277308 126216 277360 126268
rect 303712 126216 303764 126268
rect 306380 126216 306432 126268
rect 315488 126216 315540 126268
rect 318064 126216 318116 126268
rect 357256 126216 357308 126268
rect 375380 126216 375432 126268
rect 379888 126216 379940 126268
rect 400864 126216 400916 126268
rect 404452 126216 404504 126268
rect 436744 126216 436796 126268
rect 442540 126216 442592 126268
rect 482284 126216 482336 126268
rect 492404 126216 492456 126268
rect 568580 126216 568632 126268
rect 63408 126148 63460 126200
rect 116768 126148 116820 126200
rect 144184 126148 144236 126200
rect 168472 126148 168524 126200
rect 169668 126148 169720 126200
rect 70216 126080 70268 126132
rect 122196 126080 122248 126132
rect 148324 126080 148376 126132
rect 68284 126012 68336 126064
rect 114100 126012 114152 126064
rect 151084 126012 151136 126064
rect 58624 125944 58676 125996
rect 102232 125944 102284 125996
rect 50344 125876 50396 125928
rect 91192 125876 91244 125928
rect 164884 126080 164936 126132
rect 171232 126080 171284 126132
rect 173808 126148 173860 126200
rect 201132 126148 201184 126200
rect 202788 126148 202840 126200
rect 222936 126148 222988 126200
rect 226984 126148 227036 126200
rect 241060 126148 241112 126200
rect 251824 126148 251876 126200
rect 260104 126148 260156 126200
rect 456156 126148 456208 126200
rect 476764 126148 476816 126200
rect 483388 126148 483440 126200
rect 529204 126148 529256 126200
rect 173164 126080 173216 126132
rect 186596 126080 186648 126132
rect 186964 126080 187016 126132
rect 210240 126080 210292 126132
rect 211068 126080 211120 126132
rect 230204 126080 230256 126132
rect 231768 126080 231820 126132
rect 245476 126080 245528 126132
rect 277308 126080 277360 126132
rect 280068 126080 280120 126132
rect 472624 126080 472676 126132
rect 477868 126080 477920 126132
rect 522304 126080 522356 126132
rect 180064 126012 180116 126064
rect 196624 126012 196676 126064
rect 198648 126012 198700 126064
rect 220176 126012 220228 126064
rect 222108 126012 222160 126064
rect 238300 126012 238352 126064
rect 462504 126012 462556 126064
rect 504364 126012 504416 126064
rect 510528 126012 510580 126064
rect 533436 126012 533488 126064
rect 172980 125944 173032 125996
rect 181444 125944 181496 125996
rect 202052 125944 202104 125996
rect 204168 125944 204220 125996
rect 224684 125944 224736 125996
rect 233148 125944 233200 125996
rect 246488 125944 246540 125996
rect 260104 125944 260156 125996
rect 262864 125944 262916 125996
rect 451556 125944 451608 125996
rect 483664 125944 483716 125996
rect 486056 125944 486108 125996
rect 526444 125944 526496 125996
rect 167552 125876 167604 125928
rect 184204 125876 184256 125928
rect 204812 125876 204864 125928
rect 208308 125876 208360 125928
rect 227444 125876 227496 125928
rect 491484 125876 491536 125928
rect 507860 125876 507912 125928
rect 520924 125876 520976 125928
rect 53104 125808 53156 125860
rect 77760 125808 77812 125860
rect 178684 125808 178736 125860
rect 192024 125808 192076 125860
rect 205548 125808 205600 125860
rect 215208 125808 215260 125860
rect 232872 125808 232924 125860
rect 262864 125808 262916 125860
rect 269212 125808 269264 125860
rect 270408 125808 270460 125860
rect 275560 125808 275612 125860
rect 505008 125808 505060 125860
rect 213184 125740 213236 125792
rect 229284 125740 229336 125792
rect 259368 125740 259420 125792
rect 266452 125740 266504 125792
rect 269028 125740 269080 125792
rect 273720 125740 273772 125792
rect 309048 125740 309100 125792
rect 313280 125740 313332 125792
rect 219348 125672 219400 125724
rect 235632 125672 235684 125724
rect 264244 125672 264296 125724
rect 267372 125672 267424 125724
rect 271788 125672 271840 125724
rect 276388 125672 276440 125724
rect 280804 125672 280856 125724
rect 282736 125672 282788 125724
rect 282828 125672 282880 125724
rect 284392 125672 284444 125724
rect 301964 125672 302016 125724
rect 303620 125672 303672 125724
rect 308312 125672 308364 125724
rect 311900 125672 311952 125724
rect 319168 125672 319220 125724
rect 322204 125672 322256 125724
rect 326436 125672 326488 125724
rect 331772 125672 331824 125724
rect 333704 125672 333756 125724
rect 334624 125672 334676 125724
rect 337292 125672 337344 125724
rect 340144 125672 340196 125724
rect 348148 125672 348200 125724
rect 353944 125672 353996 125724
rect 356336 125672 356388 125724
rect 357348 125672 357400 125724
rect 369032 125672 369084 125724
rect 371884 125672 371936 125724
rect 445208 125672 445260 125724
rect 447784 125672 447836 125724
rect 72424 125604 72476 125656
rect 74172 125604 74224 125656
rect 39304 125468 39356 125520
rect 75092 125468 75144 125520
rect 32404 125400 32456 125452
rect 81440 125400 81492 125452
rect 66168 125332 66220 125384
rect 118608 125604 118660 125656
rect 129004 125604 129056 125656
rect 132224 125604 132276 125656
rect 133144 125604 133196 125656
rect 137652 125604 137704 125656
rect 183652 125604 183704 125656
rect 184848 125604 184900 125656
rect 206284 125604 206336 125656
rect 207480 125604 207532 125656
rect 242164 125604 242216 125656
rect 248328 125604 248380 125656
rect 249156 125604 249208 125656
rect 254676 125604 254728 125656
rect 262956 125604 263008 125656
rect 265532 125604 265584 125656
rect 268384 125604 268436 125656
rect 270960 125604 271012 125656
rect 273904 125604 273956 125656
rect 274640 125604 274692 125656
rect 278688 125604 278740 125656
rect 281908 125604 281960 125656
rect 282184 125604 282236 125656
rect 283656 125604 283708 125656
rect 288348 125604 288400 125656
rect 289084 125604 289136 125656
rect 289912 125604 289964 125656
rect 290924 125604 290976 125656
rect 292580 125604 292632 125656
rect 293684 125604 293736 125656
rect 297364 125604 297416 125656
rect 298100 125604 298152 125656
rect 298284 125604 298336 125656
rect 299296 125604 299348 125656
rect 300124 125604 300176 125656
rect 300768 125604 300820 125656
rect 301044 125604 301096 125656
rect 302240 125604 302292 125656
rect 302792 125604 302844 125656
rect 305000 125604 305052 125656
rect 305552 125604 305604 125656
rect 306288 125604 306340 125656
rect 306472 125604 306524 125656
rect 309140 125604 309192 125656
rect 310980 125604 311032 125656
rect 311716 125604 311768 125656
rect 313740 125604 313792 125656
rect 314476 125604 314528 125656
rect 316408 125604 316460 125656
rect 317236 125604 317288 125656
rect 318248 125604 318300 125656
rect 318708 125604 318760 125656
rect 320088 125604 320140 125656
rect 320824 125604 320876 125656
rect 321008 125604 321060 125656
rect 321468 125604 321520 125656
rect 321836 125604 321888 125656
rect 322848 125604 322900 125656
rect 323676 125604 323728 125656
rect 324228 125604 324280 125656
rect 324596 125604 324648 125656
rect 325516 125604 325568 125656
rect 327356 125604 327408 125656
rect 328368 125604 328420 125656
rect 329104 125604 329156 125656
rect 329748 125604 329800 125656
rect 330024 125604 330076 125656
rect 331128 125604 331180 125656
rect 331864 125604 331916 125656
rect 332508 125604 332560 125656
rect 334532 125604 334584 125656
rect 335268 125604 335320 125656
rect 335452 125604 335504 125656
rect 336556 125604 336608 125656
rect 338212 125604 338264 125656
rect 339316 125604 339368 125656
rect 340052 125604 340104 125656
rect 340788 125604 340840 125656
rect 340972 125604 341024 125656
rect 342076 125604 342128 125656
rect 342720 125604 342772 125656
rect 343548 125604 343600 125656
rect 345480 125604 345532 125656
rect 346308 125604 346360 125656
rect 349988 125604 350040 125656
rect 350448 125604 350500 125656
rect 352748 125604 352800 125656
rect 353208 125604 353260 125656
rect 353668 125604 353720 125656
rect 354588 125604 354640 125656
rect 355416 125604 355468 125656
rect 356704 125604 356756 125656
rect 358176 125604 358228 125656
rect 358728 125604 358780 125656
rect 359096 125604 359148 125656
rect 360108 125604 360160 125656
rect 360844 125604 360896 125656
rect 361488 125604 361540 125656
rect 361764 125604 361816 125656
rect 362868 125604 362920 125656
rect 363604 125604 363656 125656
rect 364248 125604 364300 125656
rect 364524 125604 364576 125656
rect 365628 125604 365680 125656
rect 366364 125604 366416 125656
rect 367008 125604 367060 125656
rect 367192 125604 367244 125656
rect 368388 125604 368440 125656
rect 369952 125604 370004 125656
rect 371148 125604 371200 125656
rect 371792 125604 371844 125656
rect 372528 125604 372580 125656
rect 372712 125604 372764 125656
rect 373908 125604 373960 125656
rect 374460 125604 374512 125656
rect 375196 125604 375248 125656
rect 381728 125604 381780 125656
rect 382188 125604 382240 125656
rect 382648 125604 382700 125656
rect 383476 125604 383528 125656
rect 384488 125604 384540 125656
rect 384948 125604 385000 125656
rect 385408 125604 385460 125656
rect 386236 125604 386288 125656
rect 387156 125604 387208 125656
rect 387708 125604 387760 125656
rect 389916 125604 389968 125656
rect 390468 125604 390520 125656
rect 390836 125604 390888 125656
rect 392584 125604 392636 125656
rect 392676 125604 392728 125656
rect 393228 125604 393280 125656
rect 395344 125604 395396 125656
rect 395988 125604 396040 125656
rect 396264 125604 396316 125656
rect 397276 125604 397328 125656
rect 398104 125604 398156 125656
rect 398748 125604 398800 125656
rect 400772 125604 400824 125656
rect 401508 125604 401560 125656
rect 403532 125604 403584 125656
rect 404268 125604 404320 125656
rect 406200 125604 406252 125656
rect 407028 125604 407080 125656
rect 408960 125604 409012 125656
rect 409788 125604 409840 125656
rect 411720 125604 411772 125656
rect 412548 125604 412600 125656
rect 413468 125604 413520 125656
rect 413928 125604 413980 125656
rect 414388 125604 414440 125656
rect 415308 125604 415360 125656
rect 416228 125604 416280 125656
rect 416688 125604 416740 125656
rect 417148 125604 417200 125656
rect 418068 125604 418120 125656
rect 418896 125604 418948 125656
rect 419448 125604 419500 125656
rect 421656 125604 421708 125656
rect 422208 125604 422260 125656
rect 422576 125604 422628 125656
rect 423588 125604 423640 125656
rect 424416 125604 424468 125656
rect 424968 125604 425020 125656
rect 425244 125604 425296 125656
rect 426348 125604 426400 125656
rect 427084 125604 427136 125656
rect 427728 125604 427780 125656
rect 428004 125604 428056 125656
rect 429108 125604 429160 125656
rect 429844 125604 429896 125656
rect 430488 125604 430540 125656
rect 430764 125604 430816 125656
rect 431868 125604 431920 125656
rect 432512 125604 432564 125656
rect 433248 125604 433300 125656
rect 433432 125604 433484 125656
rect 434628 125604 434680 125656
rect 435272 125604 435324 125656
rect 436008 125604 436060 125656
rect 436192 125604 436244 125656
rect 437388 125604 437440 125656
rect 438032 125604 438084 125656
rect 439504 125604 439556 125656
rect 443460 125604 443512 125656
rect 444196 125604 444248 125656
rect 446128 125604 446180 125656
rect 446956 125604 447008 125656
rect 447968 125604 448020 125656
rect 448428 125604 448480 125656
rect 450728 125604 450780 125656
rect 451188 125604 451240 125656
rect 453396 125604 453448 125656
rect 453948 125604 454000 125656
rect 454316 125604 454368 125656
rect 455236 125604 455288 125656
rect 458824 125604 458876 125656
rect 459468 125604 459520 125656
rect 461584 125604 461636 125656
rect 462228 125604 462280 125656
rect 464252 125604 464304 125656
rect 464988 125604 465040 125656
rect 465172 125604 465224 125656
rect 466368 125604 466420 125656
rect 467012 125604 467064 125656
rect 467748 125604 467800 125656
rect 467932 125604 467984 125656
rect 469036 125604 469088 125656
rect 479708 125604 479760 125656
rect 480168 125604 480220 125656
rect 480628 125604 480680 125656
rect 485136 125604 485188 125656
rect 485688 125604 485740 125656
rect 487896 125604 487948 125656
rect 488448 125604 488500 125656
rect 490564 125604 490616 125656
rect 491208 125604 491260 125656
rect 493324 125604 493376 125656
rect 493968 125604 494020 125656
rect 496084 125604 496136 125656
rect 496728 125604 496780 125656
rect 498752 125604 498804 125656
rect 499488 125604 499540 125656
rect 501512 125604 501564 125656
rect 502248 125604 502300 125656
rect 504180 125604 504232 125656
rect 505008 125604 505060 125656
rect 506940 125604 506992 125656
rect 507768 125604 507820 125656
rect 509608 125604 509660 125656
rect 510528 125604 510580 125656
rect 511448 125604 511500 125656
rect 511908 125604 511960 125656
rect 512368 125604 512420 125656
rect 513288 125604 513340 125656
rect 514208 125604 514260 125656
rect 514668 125604 514720 125656
rect 515404 125604 515456 125656
rect 516048 125604 516100 125656
rect 507860 125400 507912 125452
rect 550640 125400 550692 125452
rect 536840 125332 536892 125384
rect 33784 125264 33836 125316
rect 85028 125264 85080 125316
rect 475200 125264 475252 125316
rect 529940 125264 529992 125316
rect 18604 125196 18656 125248
rect 69572 125196 69624 125248
rect 481640 125196 481692 125248
rect 538220 125196 538272 125248
rect 62028 125128 62080 125180
rect 115848 125128 115900 125180
rect 488816 125128 488868 125180
rect 547880 125128 547932 125180
rect 55128 125060 55180 125112
rect 110420 125060 110472 125112
rect 494244 125060 494296 125112
rect 554780 125060 554832 125112
rect 52368 124992 52420 125044
rect 107660 124992 107712 125044
rect 496912 124992 496964 125044
rect 557540 124992 557592 125044
rect 48228 124924 48280 124976
rect 104992 124924 105044 124976
rect 499672 124924 499724 124976
rect 561680 124924 561732 124976
rect 4804 124856 4856 124908
rect 70492 124856 70544 124908
rect 111616 124856 111668 124908
rect 152556 124856 152608 124908
rect 502432 124856 502484 124908
rect 564532 124856 564584 124908
rect 41328 123564 41380 123616
rect 88248 123564 88300 123616
rect 37188 123496 37240 123548
rect 88984 123496 89036 123548
rect 35164 123428 35216 123480
rect 94136 123428 94188 123480
rect 507676 123428 507728 123480
rect 572812 123428 572864 123480
rect 455236 90312 455288 90364
rect 502340 90312 502392 90364
rect 3516 88952 3568 89004
rect 67640 88952 67692 89004
rect 447784 88952 447836 89004
rect 490012 88952 490064 89004
rect 533436 50328 533488 50380
rect 575480 50328 575532 50380
rect 84108 48968 84160 49020
rect 129004 48968 129056 49020
rect 102048 26868 102100 26920
rect 126244 26868 126296 26920
rect 126888 26868 126940 26920
rect 164240 26868 164292 26920
rect 459468 26868 459520 26920
rect 507860 26868 507912 26920
rect 91008 18572 91060 18624
rect 133144 18572 133196 18624
rect 133788 15920 133840 15972
rect 169760 15920 169812 15972
rect 86868 15852 86920 15904
rect 134156 15852 134208 15904
rect 439504 15852 439556 15904
rect 481732 15852 481784 15904
rect 115848 11704 115900 11756
rect 155960 11704 156012 11756
rect 386236 11704 386288 11756
rect 412640 11704 412692 11756
rect 450544 11704 450596 11756
rect 484768 11704 484820 11756
rect 77116 10276 77168 10328
rect 125692 10276 125744 10328
rect 426256 10276 426308 10328
rect 465816 10276 465868 10328
rect 469036 10276 469088 10328
rect 520280 10276 520332 10328
rect 519544 9596 519596 9648
rect 526628 9596 526680 9648
rect 444196 8984 444248 9036
rect 488816 8984 488868 9036
rect 130568 8916 130620 8968
rect 144184 8916 144236 8968
rect 143540 8848 143592 8900
rect 178132 8916 178184 8968
rect 467748 8916 467800 8968
rect 519544 8916 519596 8968
rect 526444 8916 526496 8968
rect 544384 8916 544436 8968
rect 79692 7624 79744 7676
rect 128452 7624 128504 7676
rect 464344 7624 464396 7676
rect 506480 7624 506532 7676
rect 44272 7556 44324 7608
rect 58624 7556 58676 7608
rect 58440 7488 58492 7540
rect 112536 7556 112588 7608
rect 129372 7556 129424 7608
rect 151084 7556 151136 7608
rect 372528 7556 372580 7608
rect 395344 7556 395396 7608
rect 432604 7556 432656 7608
rect 459192 7556 459244 7608
rect 489736 7556 489788 7608
rect 549076 7556 549128 7608
rect 466368 6196 466420 6248
rect 517152 6196 517204 6248
rect 473268 6128 473320 6180
rect 527824 6128 527876 6180
rect 476764 5448 476816 5500
rect 505376 5448 505428 5500
rect 471244 5380 471296 5432
rect 510068 5380 510120 5432
rect 440148 5312 440200 5364
rect 483020 5312 483072 5364
rect 483664 5312 483716 5364
rect 499396 5312 499448 5364
rect 136456 5244 136508 5296
rect 148324 5244 148376 5296
rect 446956 5244 447008 5296
rect 134156 5176 134208 5228
rect 164884 5176 164936 5228
rect 407764 5176 407816 5228
rect 416688 5176 416740 5228
rect 418804 5176 418856 5228
rect 430856 5176 430908 5228
rect 448428 5176 448480 5228
rect 494704 5176 494756 5228
rect 59636 5108 59688 5160
rect 68284 5108 68336 5160
rect 69112 5108 69164 5160
rect 112444 5108 112496 5160
rect 135352 5108 135404 5160
rect 170404 5108 170456 5160
rect 392584 5108 392636 5160
rect 420184 5108 420236 5160
rect 429844 5108 429896 5160
rect 445024 5108 445076 5160
rect 453948 5108 454000 5160
rect 501788 5108 501840 5160
rect 12348 5040 12400 5092
rect 53104 5040 53156 5092
rect 30104 4972 30156 5024
rect 50344 4972 50396 5024
rect 52552 4972 52604 5024
rect 107844 5040 107896 5092
rect 131764 5040 131816 5092
rect 168656 5040 168708 5092
rect 403624 5040 403676 5092
rect 434444 5040 434496 5092
rect 451188 5040 451240 5092
rect 498200 5040 498252 5092
rect 504364 5040 504416 5092
rect 513564 5040 513616 5092
rect 104900 4972 104952 5024
rect 108120 4972 108172 5024
rect 150532 4972 150584 5024
rect 389824 4972 389876 5024
rect 402520 4972 402572 5024
rect 406936 4972 406988 5024
rect 441436 4972 441488 5024
rect 442264 4972 442316 5024
rect 452108 4972 452160 5024
rect 475384 4972 475436 5024
rect 524236 4972 524288 5024
rect 26516 4904 26568 4956
rect 88432 4904 88484 4956
rect 93952 4904 94004 4956
rect 139676 4904 139728 4956
rect 140044 4904 140096 4956
rect 175280 4904 175332 4956
rect 375196 4904 375248 4956
rect 398932 4904 398984 4956
rect 400864 4904 400916 4956
rect 406016 4904 406068 4956
rect 412456 4904 412508 4956
rect 448612 4904 448664 4956
rect 464988 4904 465040 4956
rect 515956 4904 516008 4956
rect 522304 4904 522356 4956
rect 533712 4904 533764 4956
rect 7656 4836 7708 4888
rect 72424 4836 72476 4888
rect 97448 4836 97500 4888
rect 142344 4836 142396 4888
rect 161296 4836 161348 4888
rect 178684 4836 178736 4888
rect 383476 4836 383528 4888
rect 409604 4836 409656 4888
rect 417976 4836 418028 4888
rect 455696 4836 455748 4888
rect 462228 4836 462280 4888
rect 512460 4836 512512 4888
rect 529204 4836 529256 4888
rect 540796 4836 540848 4888
rect 4068 4768 4120 4820
rect 70400 4768 70452 4820
rect 72608 4768 72660 4820
rect 122104 4768 122156 4820
rect 128176 4768 128228 4820
rect 165712 4768 165764 4820
rect 371884 4768 371936 4820
rect 391756 4768 391808 4820
rect 397276 4768 397328 4820
rect 427268 4768 427320 4820
rect 431776 4768 431828 4820
rect 473452 4768 473504 4820
rect 475936 4768 475988 4820
rect 531320 4768 531372 4820
rect 536104 4768 536156 4820
rect 541992 4768 542044 4820
rect 547144 4768 547196 4820
rect 552664 4768 552716 4820
rect 50896 4700 50948 4752
rect 479524 4700 479576 4752
rect 495900 4700 495952 4752
rect 471336 4632 471388 4684
rect 480536 4632 480588 4684
rect 492312 4564 492364 4616
rect 421564 4428 421616 4480
rect 423772 4428 423824 4480
rect 483020 4224 483072 4276
rect 484032 4224 484084 4276
rect 126980 4156 127032 4208
rect 130384 4156 130436 4208
rect 436744 4156 436796 4208
rect 437940 4156 437992 4208
rect 461584 4156 461636 4208
rect 462780 4156 462832 4208
rect 467104 4156 467156 4208
rect 469864 4156 469916 4208
rect 472624 4156 472676 4208
rect 476948 4156 477000 4208
rect 482284 4156 482336 4208
rect 487620 4156 487672 4208
rect 520924 4156 520976 4208
rect 523040 4156 523092 4208
rect 533344 4156 533396 4208
rect 534908 4156 534960 4208
rect 543004 4156 543056 4208
rect 545488 4156 545540 4208
rect 34796 4088 34848 4140
rect 99748 4088 99800 4140
rect 102232 4088 102284 4140
rect 146392 4088 146444 4140
rect 163688 4088 163740 4140
rect 193220 4088 193272 4140
rect 219256 4088 219308 4140
rect 220084 4088 220136 4140
rect 286600 4088 286652 4140
rect 287152 4088 287204 4140
rect 296628 4088 296680 4140
rect 297272 4088 297324 4140
rect 304908 4088 304960 4140
rect 307944 4088 307996 4140
rect 331864 4088 331916 4140
rect 336280 4088 336332 4140
rect 336648 4088 336700 4140
rect 349252 4088 349304 4140
rect 356704 4088 356756 4140
rect 374092 4088 374144 4140
rect 375288 4088 375340 4140
rect 400036 4088 400088 4140
rect 400128 4088 400180 4140
rect 432052 4088 432104 4140
rect 38384 4020 38436 4072
rect 96712 4020 96764 4072
rect 103336 4020 103388 4072
rect 146300 4020 146352 4072
rect 164884 4020 164936 4072
rect 194692 4020 194744 4072
rect 242900 4020 242952 4072
rect 249156 4020 249208 4072
rect 253480 4020 253532 4072
rect 260104 4020 260156 4072
rect 273628 4020 273680 4072
rect 277492 4020 277544 4072
rect 325516 4020 325568 4072
rect 333888 4020 333940 4072
rect 339408 4020 339460 4072
rect 352840 4020 352892 4072
rect 354588 4020 354640 4072
rect 371700 4020 371752 4072
rect 373816 4020 373868 4072
rect 397736 4020 397788 4072
rect 402888 4020 402940 4072
rect 21824 3952 21876 4004
rect 33784 3952 33836 4004
rect 39580 3952 39632 4004
rect 98000 3952 98052 4004
rect 17040 3884 17092 3936
rect 32404 3884 32456 3936
rect 35992 3884 36044 3936
rect 93860 3884 93912 3936
rect 102416 3952 102468 4004
rect 105728 3952 105780 4004
rect 149152 3952 149204 4004
rect 155408 3952 155460 4004
rect 186412 3952 186464 4004
rect 324228 3952 324280 4004
rect 332692 3952 332744 4004
rect 342076 3952 342128 4004
rect 355232 3952 355284 4004
rect 361488 3952 361540 4004
rect 381176 3952 381228 4004
rect 382188 3952 382240 4004
rect 99840 3884 99892 3936
rect 144920 3884 144972 3936
rect 151820 3884 151872 3936
rect 183652 3884 183704 3936
rect 200304 3884 200356 3936
rect 220912 3884 220964 3936
rect 328368 3884 328420 3936
rect 337476 3884 337528 3936
rect 345664 3884 345716 3936
rect 359924 3884 359976 3936
rect 360108 3884 360160 3936
rect 378876 3884 378928 3936
rect 379428 3884 379480 3936
rect 404820 3884 404872 3936
rect 5264 3816 5316 3868
rect 7564 3816 7616 3868
rect 31300 3816 31352 3868
rect 91284 3816 91336 3868
rect 91560 3816 91612 3868
rect 138020 3816 138072 3868
rect 156604 3816 156656 3868
rect 187700 3816 187752 3868
rect 193220 3816 193272 3868
rect 215392 3816 215444 3868
rect 332508 3816 332560 3868
rect 343364 3816 343416 3868
rect 343548 3816 343600 3868
rect 357532 3816 357584 3868
rect 358728 3816 358780 3868
rect 377680 3816 377732 3868
rect 378048 3816 378100 3868
rect 403624 3816 403676 3868
rect 407028 3952 407080 4004
rect 437388 4088 437440 4140
rect 479340 4088 479392 4140
rect 498016 4088 498068 4140
rect 559748 4088 559800 4140
rect 435548 4020 435600 4072
rect 436008 4020 436060 4072
rect 478144 4020 478196 4072
rect 495256 4020 495308 4072
rect 556160 4020 556212 4072
rect 433156 3952 433208 4004
rect 440332 3952 440384 4004
rect 441528 3952 441580 4004
rect 486424 3952 486476 4004
rect 502248 3952 502300 4004
rect 564440 3952 564492 4004
rect 405648 3884 405700 3936
rect 439136 3884 439188 3936
rect 444288 3884 444340 3936
rect 489920 3884 489972 3936
rect 505008 3884 505060 3936
rect 568028 3884 568080 3936
rect 408224 3816 408276 3868
rect 408316 3816 408368 3868
rect 442632 3816 442684 3868
rect 447048 3816 447100 3868
rect 493508 3816 493560 3868
rect 500776 3816 500828 3868
rect 563244 3816 563296 3868
rect 14740 3748 14792 3800
rect 17224 3748 17276 3800
rect 32404 3748 32456 3800
rect 92480 3748 92532 3800
rect 92756 3748 92808 3800
rect 93768 3748 93820 3800
rect 95148 3748 95200 3800
rect 140780 3748 140832 3800
rect 149520 3748 149572 3800
rect 176844 3748 176896 3800
rect 180248 3748 180300 3800
rect 180708 3748 180760 3800
rect 196808 3748 196860 3800
rect 218152 3748 218204 3800
rect 322848 3748 322900 3800
rect 330392 3748 330444 3800
rect 331128 3748 331180 3800
rect 340972 3748 341024 3800
rect 342168 3748 342220 3800
rect 356336 3748 356388 3800
rect 362868 3748 362920 3800
rect 382372 3748 382424 3800
rect 383568 3748 383620 3800
rect 410800 3748 410852 3800
rect 411168 3748 411220 3800
rect 446220 3748 446272 3800
rect 449716 3748 449768 3800
rect 497096 3748 497148 3800
rect 503536 3748 503588 3800
rect 566832 3748 566884 3800
rect 25320 3680 25372 3732
rect 19432 3612 19484 3664
rect 6460 3544 6512 3596
rect 14464 3544 14516 3596
rect 2872 3476 2924 3528
rect 4804 3476 4856 3528
rect 18604 3544 18656 3596
rect 23020 3544 23072 3596
rect 27712 3612 27764 3664
rect 29644 3612 29696 3664
rect 33600 3612 33652 3664
rect 35164 3612 35216 3664
rect 1676 3408 1728 3460
rect 18236 3476 18288 3528
rect 21364 3476 21416 3528
rect 24216 3476 24268 3528
rect 25504 3476 25556 3528
rect 76104 3544 76156 3596
rect 82912 3544 82964 3596
rect 84476 3680 84528 3732
rect 123300 3680 123352 3732
rect 132592 3680 132644 3732
rect 136732 3680 136784 3732
rect 149060 3680 149112 3732
rect 150624 3680 150676 3732
rect 183560 3680 183612 3732
rect 189724 3680 189776 3732
rect 212632 3680 212684 3732
rect 317328 3680 317380 3732
rect 324412 3680 324464 3732
rect 329748 3680 329800 3732
rect 339868 3680 339920 3732
rect 340788 3680 340840 3732
rect 354036 3680 354088 3732
rect 354496 3680 354548 3732
rect 372896 3680 372948 3732
rect 380808 3680 380860 3732
rect 407212 3680 407264 3732
rect 413928 3680 413980 3732
rect 418068 3680 418120 3732
rect 87052 3544 87104 3596
rect 85764 3476 85816 3528
rect 95240 3612 95292 3664
rect 98644 3612 98696 3664
rect 99288 3612 99340 3664
rect 101036 3612 101088 3664
rect 102048 3612 102100 3664
rect 142160 3612 142212 3664
rect 147128 3612 147180 3664
rect 87972 3544 88024 3596
rect 135260 3544 135312 3596
rect 145932 3544 145984 3596
rect 174268 3612 174320 3664
rect 181444 3612 181496 3664
rect 182548 3612 182600 3664
rect 188528 3612 188580 3664
rect 188988 3612 189040 3664
rect 180984 3544 181036 3596
rect 186136 3544 186188 3596
rect 89720 3476 89772 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 11152 3408 11204 3460
rect 75000 3408 75052 3460
rect 75828 3408 75880 3460
rect 76196 3408 76248 3460
rect 77116 3408 77168 3460
rect 77392 3408 77444 3460
rect 78496 3408 78548 3460
rect 83280 3408 83332 3460
rect 84108 3408 84160 3460
rect 85672 3408 85724 3460
rect 89168 3408 89220 3460
rect 132960 3476 133012 3528
rect 133788 3476 133840 3528
rect 141240 3476 141292 3528
rect 142068 3476 142120 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 173164 3476 173216 3528
rect 173808 3476 173860 3528
rect 123484 3408 123536 3460
rect 124128 3408 124180 3460
rect 124680 3408 124732 3460
rect 125324 3408 125376 3460
rect 125876 3408 125928 3460
rect 126888 3408 126940 3460
rect 127072 3408 127124 3460
rect 133880 3408 133932 3460
rect 138848 3408 138900 3460
rect 174084 3408 174136 3460
rect 176660 3476 176712 3528
rect 177948 3476 178000 3528
rect 179512 3476 179564 3528
rect 183744 3476 183796 3528
rect 184848 3476 184900 3528
rect 184940 3476 184992 3528
rect 186964 3476 187016 3528
rect 208492 3612 208544 3664
rect 277124 3612 277176 3664
rect 280344 3612 280396 3664
rect 321468 3612 321520 3664
rect 329196 3612 329248 3664
rect 331036 3612 331088 3664
rect 342168 3612 342220 3664
rect 346308 3612 346360 3664
rect 361120 3612 361172 3664
rect 362776 3612 362828 3664
rect 383568 3612 383620 3664
rect 387708 3612 387760 3664
rect 415492 3612 415544 3664
rect 416596 3612 416648 3664
rect 419448 3612 419500 3664
rect 449808 3680 449860 3732
rect 452568 3680 452620 3732
rect 500592 3680 500644 3732
rect 507768 3680 507820 3732
rect 571524 3680 571576 3732
rect 201500 3476 201552 3528
rect 202788 3476 202840 3528
rect 205088 3476 205140 3528
rect 205548 3476 205600 3528
rect 179052 3408 179104 3460
rect 205732 3408 205784 3460
rect 8760 3340 8812 3392
rect 39304 3340 39356 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 51356 3340 51408 3392
rect 52368 3340 52420 3392
rect 103612 3340 103664 3392
rect 110512 3340 110564 3392
rect 111708 3340 111760 3392
rect 112812 3340 112864 3392
rect 154580 3340 154632 3392
rect 157800 3340 157852 3392
rect 158628 3340 158680 3392
rect 158904 3340 158956 3392
rect 160008 3340 160060 3392
rect 160100 3340 160152 3392
rect 190552 3340 190604 3392
rect 190828 3340 190880 3392
rect 191748 3340 191800 3392
rect 192024 3340 192076 3392
rect 193128 3340 193180 3392
rect 194416 3340 194468 3392
rect 195244 3340 195296 3392
rect 197912 3340 197964 3392
rect 198648 3340 198700 3392
rect 199108 3340 199160 3392
rect 200028 3340 200080 3392
rect 211160 3544 211212 3596
rect 206192 3476 206244 3528
rect 206928 3476 206980 3528
rect 208584 3476 208636 3528
rect 209688 3476 209740 3528
rect 213368 3476 213420 3528
rect 213828 3476 213880 3528
rect 214472 3476 214524 3528
rect 215208 3476 215260 3528
rect 215668 3476 215720 3528
rect 216588 3476 216640 3528
rect 218060 3476 218112 3528
rect 219348 3476 219400 3528
rect 222752 3476 222804 3528
rect 223488 3476 223540 3528
rect 223948 3476 224000 3528
rect 224868 3476 224920 3528
rect 226340 3476 226392 3528
rect 227628 3476 227680 3528
rect 231032 3476 231084 3528
rect 231768 3476 231820 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 234620 3476 234672 3528
rect 242164 3544 242216 3596
rect 247592 3544 247644 3596
rect 249064 3544 249116 3596
rect 241704 3476 241756 3528
rect 242808 3476 242860 3528
rect 244096 3476 244148 3528
rect 244924 3476 244976 3528
rect 246396 3476 246448 3528
rect 246948 3476 247000 3528
rect 248788 3476 248840 3528
rect 250444 3476 250496 3528
rect 252376 3476 252428 3528
rect 253204 3476 253256 3528
rect 254676 3476 254728 3528
rect 255228 3476 255280 3528
rect 255872 3476 255924 3528
rect 256608 3476 256660 3528
rect 257068 3476 257120 3528
rect 262956 3544 263008 3596
rect 292580 3544 292632 3596
rect 293684 3544 293736 3596
rect 314476 3544 314528 3596
rect 319720 3544 319772 3596
rect 328276 3544 328328 3596
rect 338672 3544 338724 3596
rect 343456 3544 343508 3596
rect 358728 3544 358780 3596
rect 360016 3544 360068 3596
rect 379980 3544 380032 3596
rect 386328 3544 386380 3596
rect 414296 3544 414348 3596
rect 415308 3544 415360 3596
rect 421380 3544 421432 3596
rect 454500 3612 454552 3664
rect 458088 3612 458140 3664
rect 507676 3612 507728 3664
rect 509148 3612 509200 3664
rect 573916 3612 573968 3664
rect 261760 3476 261812 3528
rect 262864 3476 262916 3528
rect 266544 3476 266596 3528
rect 267648 3476 267700 3528
rect 267740 3476 267792 3528
rect 269028 3476 269080 3528
rect 271236 3476 271288 3528
rect 271788 3476 271840 3528
rect 276020 3476 276072 3528
rect 277308 3476 277360 3528
rect 281908 3476 281960 3528
rect 282828 3476 282880 3528
rect 283104 3476 283156 3528
rect 284484 3476 284536 3528
rect 288992 3476 289044 3528
rect 289728 3476 289780 3528
rect 293960 3476 294012 3528
rect 294880 3476 294932 3528
rect 295340 3476 295392 3528
rect 296076 3476 296128 3528
rect 300768 3476 300820 3528
rect 301964 3476 302016 3528
rect 318156 3476 318208 3528
rect 322112 3476 322164 3528
rect 325608 3476 325660 3528
rect 335084 3476 335136 3528
rect 229836 3408 229888 3460
rect 231124 3408 231176 3460
rect 238116 3408 238168 3460
rect 238668 3408 238720 3460
rect 251180 3408 251232 3460
rect 252468 3408 252520 3460
rect 259460 3408 259512 3460
rect 264244 3408 264296 3460
rect 265348 3408 265400 3460
rect 267004 3408 267056 3460
rect 306288 3408 306340 3460
rect 309048 3408 309100 3460
rect 314568 3408 314620 3460
rect 320916 3408 320968 3460
rect 322756 3408 322808 3460
rect 331588 3408 331640 3460
rect 334624 3408 334676 3460
rect 345756 3476 345808 3528
rect 346216 3476 346268 3528
rect 362316 3476 362368 3528
rect 365536 3476 365588 3528
rect 387156 3476 387208 3528
rect 389088 3476 389140 3528
rect 417884 3476 417936 3528
rect 422208 3476 422260 3528
rect 453304 3544 453356 3596
rect 455328 3544 455380 3596
rect 504180 3544 504232 3596
rect 506388 3544 506440 3596
rect 570328 3544 570380 3596
rect 336556 3408 336608 3460
rect 348056 3408 348108 3460
rect 349068 3408 349120 3460
rect 365812 3408 365864 3460
rect 368296 3408 368348 3460
rect 390652 3408 390704 3460
rect 391848 3408 391900 3460
rect 424968 3408 425020 3460
rect 456892 3476 456944 3528
rect 460848 3476 460900 3528
rect 511264 3476 511316 3528
rect 511908 3476 511960 3528
rect 577412 3476 577464 3528
rect 460388 3408 460440 3460
rect 463608 3408 463660 3460
rect 514760 3408 514812 3460
rect 516048 3408 516100 3460
rect 583392 3408 583444 3460
rect 227536 3340 227588 3392
rect 238024 3340 238076 3392
rect 279516 3340 279568 3392
rect 280804 3340 280856 3392
rect 311808 3340 311860 3392
rect 317328 3340 317380 3392
rect 318708 3340 318760 3392
rect 325608 3340 325660 3392
rect 339316 3340 339368 3392
rect 351644 3340 351696 3392
rect 353208 3340 353260 3392
rect 370596 3340 370648 3392
rect 371056 3340 371108 3392
rect 394240 3340 394292 3392
rect 397368 3340 397420 3392
rect 428464 3340 428516 3392
rect 474556 3340 474608 3392
rect 499488 3340 499540 3392
rect 560852 3340 560904 3392
rect 28908 3272 28960 3324
rect 43076 3272 43128 3324
rect 41880 3204 41932 3256
rect 572 3136 624 3188
rect 3424 3136 3476 3188
rect 45468 3136 45520 3188
rect 96252 3272 96304 3324
rect 106924 3272 106976 3324
rect 142436 3272 142488 3324
rect 166080 3272 166132 3324
rect 166908 3272 166960 3324
rect 171968 3272 172020 3324
rect 200212 3272 200264 3324
rect 209780 3272 209832 3324
rect 213184 3272 213236 3324
rect 262956 3272 263008 3324
rect 269396 3272 269448 3324
rect 287796 3272 287848 3324
rect 288348 3272 288400 3324
rect 310428 3272 310480 3324
rect 315028 3272 315080 3324
rect 320824 3272 320876 3324
rect 328000 3272 328052 3324
rect 335268 3272 335320 3324
rect 346952 3272 347004 3324
rect 357348 3272 357400 3324
rect 375288 3272 375340 3324
rect 376668 3272 376720 3324
rect 401324 3272 401376 3324
rect 401508 3272 401560 3324
rect 433248 3272 433300 3324
rect 434628 3272 434680 3324
rect 109316 3204 109368 3256
rect 152004 3204 152056 3256
rect 100852 3136 100904 3188
rect 115204 3136 115256 3188
rect 115848 3136 115900 3188
rect 116400 3136 116452 3188
rect 117228 3136 117280 3188
rect 154672 3204 154724 3256
rect 168380 3204 168432 3256
rect 197452 3204 197504 3256
rect 216864 3204 216916 3256
rect 217968 3204 218020 3256
rect 258264 3204 258316 3256
rect 259368 3204 259420 3256
rect 307668 3204 307720 3256
rect 311440 3204 311492 3256
rect 317236 3204 317288 3256
rect 323308 3204 323360 3256
rect 340144 3204 340196 3256
rect 350448 3204 350500 3256
rect 351828 3204 351880 3256
rect 369400 3204 369452 3256
rect 373908 3204 373960 3256
rect 396540 3204 396592 3256
rect 404268 3204 404320 3256
rect 409788 3204 409840 3256
rect 436468 3204 436520 3256
rect 471060 3272 471112 3324
rect 496728 3272 496780 3324
rect 557356 3272 557408 3324
rect 475752 3204 475804 3256
rect 493968 3204 494020 3256
rect 553768 3204 553820 3256
rect 50160 3068 50212 3120
rect 106280 3068 106332 3120
rect 114008 3068 114060 3120
rect 154212 3136 154264 3188
rect 173072 3136 173124 3188
rect 175464 3136 175516 3188
rect 202972 3136 203024 3188
rect 207388 3136 207440 3188
rect 208308 3136 208360 3188
rect 239312 3136 239364 3188
rect 246304 3136 246356 3188
rect 280712 3136 280764 3188
rect 282184 3136 282236 3188
rect 311716 3136 311768 3188
rect 316224 3136 316276 3188
rect 347688 3136 347740 3188
rect 363512 3136 363564 3188
rect 371148 3136 371200 3188
rect 393044 3136 393096 3188
rect 394608 3136 394660 3188
rect 422576 3136 422628 3188
rect 423588 3136 423640 3188
rect 424876 3136 424928 3188
rect 427728 3136 427780 3188
rect 463976 3136 464028 3188
rect 491208 3136 491260 3188
rect 550272 3136 550324 3188
rect 117596 3068 117648 3120
rect 126060 3068 126112 3120
rect 160192 3068 160244 3120
rect 167184 3068 167236 3120
rect 180064 3068 180116 3120
rect 181444 3068 181496 3120
rect 206284 3068 206336 3120
rect 221556 3068 221608 3120
rect 222108 3068 222160 3120
rect 350356 3068 350408 3120
rect 367008 3068 367060 3120
rect 368388 3068 368440 3120
rect 389456 3068 389508 3120
rect 398748 3068 398800 3120
rect 429660 3068 429712 3120
rect 430488 3068 430540 3120
rect 9956 3000 10008 3052
rect 11704 3000 11756 3052
rect 20628 3000 20680 3052
rect 22744 3000 22796 3052
rect 46664 3000 46716 3052
rect 53748 3000 53800 3052
rect 109040 3000 109092 3052
rect 56048 2932 56100 2984
rect 56508 2932 56560 2984
rect 57244 2932 57296 2984
rect 57888 2932 57940 2984
rect 64328 2932 64380 2984
rect 64788 2932 64840 2984
rect 65524 2932 65576 2984
rect 66168 2932 66220 2984
rect 60832 2864 60884 2916
rect 114744 2932 114796 2984
rect 120264 3000 120316 3052
rect 122288 3000 122340 3052
rect 161572 3000 161624 3052
rect 177856 3000 177908 3052
rect 184204 3000 184256 3052
rect 225144 3000 225196 3052
rect 226984 3000 227036 3052
rect 240508 3000 240560 3052
rect 241428 3000 241480 3052
rect 249984 3000 250036 3052
rect 251824 3000 251876 3052
rect 272432 3000 272484 3052
rect 273996 3000 274048 3052
rect 274824 3000 274876 3052
rect 276664 3000 276716 3052
rect 322204 3000 322256 3052
rect 326804 3000 326856 3052
rect 353944 3000 353996 3052
rect 364616 3000 364668 3052
rect 366916 3000 366968 3052
rect 388260 3000 388312 3052
rect 393228 3000 393280 3052
rect 429108 3000 429160 3052
rect 468668 3068 468720 3120
rect 488448 3068 488500 3120
rect 546684 3068 546736 3120
rect 467472 3000 467524 3052
rect 485688 3000 485740 3052
rect 543188 3000 543240 3052
rect 119896 2932 119948 2984
rect 126060 2932 126112 2984
rect 157432 2932 157484 2984
rect 182272 2932 182324 2984
rect 264152 2932 264204 2984
rect 268384 2932 268436 2984
rect 365628 2932 365680 2984
rect 385960 2932 386012 2984
rect 395988 2932 396040 2984
rect 426164 2932 426216 2984
rect 461584 2932 461636 2984
rect 480168 2932 480220 2984
rect 536104 2932 536156 2984
rect 48964 2796 49016 2848
rect 50896 2796 50948 2848
rect 66720 2796 66772 2848
rect 67916 2796 67968 2848
rect 118976 2864 119028 2916
rect 121092 2864 121144 2916
rect 160468 2864 160520 2916
rect 268844 2864 268896 2916
rect 273904 2864 273956 2916
rect 284300 2864 284352 2916
rect 285680 2864 285732 2916
rect 336004 2864 336056 2916
rect 344560 2864 344612 2916
rect 364248 2864 364300 2916
rect 384764 2864 384816 2916
rect 390468 2864 390520 2916
rect 418988 2864 419040 2916
rect 450912 2864 450964 2916
rect 474648 2864 474700 2916
rect 529020 2864 529072 2916
rect 118792 2796 118844 2848
rect 158812 2796 158864 2848
rect 359464 2796 359516 2848
rect 368204 2796 368256 2848
rect 384948 2796 385000 2848
rect 411904 2796 411956 2848
rect 443828 2796 443880 2848
rect 469128 2796 469180 2848
rect 521844 2796 521896 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700670 73016 703520
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 105464 699718 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 170324 699718 170352 703520
rect 202800 700126 202828 703520
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 218992 700058 219020 703520
rect 218980 700052 219032 700058
rect 218980 699994 219032 700000
rect 235184 699718 235212 703520
rect 267660 702434 267688 703520
rect 267568 702406 267688 702434
rect 263508 700868 263560 700874
rect 263508 700810 263560 700816
rect 251088 700596 251140 700602
rect 251088 700538 251140 700544
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 4804 578332 4856 578338
rect 4804 578274 4856 578280
rect 3884 575204 3936 575210
rect 3884 575146 3936 575152
rect 3792 574864 3844 574870
rect 3792 574806 3844 574812
rect 3700 574728 3752 574734
rect 3700 574670 3752 574676
rect 3608 574456 3660 574462
rect 3608 574398 3660 574404
rect 3516 574252 3568 574258
rect 3516 574194 3568 574200
rect 3424 574184 3476 574190
rect 3424 574126 3476 574132
rect 3240 528556 3292 528562
rect 3240 528498 3292 528504
rect 3252 527921 3280 528498
rect 3238 527912 3294 527921
rect 3238 527847 3294 527856
rect 3332 516112 3384 516118
rect 3332 516054 3384 516060
rect 3344 514865 3372 516054
rect 3330 514856 3386 514865
rect 3330 514791 3386 514800
rect 3332 476060 3384 476066
rect 3332 476002 3384 476008
rect 3344 475697 3372 476002
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3332 463684 3384 463690
rect 3332 463626 3384 463632
rect 3344 462641 3372 463626
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 2832 358456 2834 358465
rect 2778 358391 2834 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 188873 3464 574126
rect 3528 293185 3556 574194
rect 3620 397497 3648 574398
rect 3712 449585 3740 574670
rect 3804 501809 3832 574806
rect 3896 553897 3924 575146
rect 3976 575068 4028 575074
rect 3976 575010 4028 575016
rect 3988 566953 4016 575010
rect 3974 566944 4030 566953
rect 3974 566879 4030 566888
rect 3882 553888 3938 553897
rect 3882 553823 3938 553832
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 449576 3754 449585
rect 3698 449511 3754 449520
rect 3606 397488 3662 397497
rect 3606 397423 3662 397432
rect 4816 358494 4844 578274
rect 14464 578264 14516 578270
rect 14464 578206 14516 578212
rect 11704 576224 11756 576230
rect 11704 576166 11756 576172
rect 11716 528562 11744 576166
rect 11704 528556 11756 528562
rect 11704 528498 11756 528504
rect 4804 358488 4856 358494
rect 4804 358430 4856 358436
rect 14476 306338 14504 578206
rect 106200 577862 106228 699654
rect 171060 577998 171088 699654
rect 235816 670812 235868 670818
rect 235816 670754 235868 670760
rect 227628 643136 227680 643142
rect 227628 643078 227680 643084
rect 223488 616888 223540 616894
rect 223488 616830 223540 616836
rect 216588 590708 216640 590714
rect 216588 590650 216640 590656
rect 216600 578202 216628 590650
rect 215760 578196 215812 578202
rect 215760 578138 215812 578144
rect 216588 578196 216640 578202
rect 216588 578138 216640 578144
rect 171048 577992 171100 577998
rect 171048 577934 171100 577940
rect 106188 577856 106240 577862
rect 106188 577798 106240 577804
rect 53104 577652 53156 577658
rect 53104 577594 53156 577600
rect 21362 577144 21418 577153
rect 21362 577079 21418 577088
rect 17224 576972 17276 576978
rect 17224 576914 17276 576920
rect 14464 306332 14516 306338
rect 14464 306274 14516 306280
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 17236 255270 17264 576914
rect 18604 576904 18656 576910
rect 18604 576846 18656 576852
rect 17224 255264 17276 255270
rect 17224 255206 17276 255212
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 18616 202842 18644 576846
rect 18604 202836 18656 202842
rect 18604 202778 18656 202784
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 21376 150414 21404 577079
rect 36544 576496 36596 576502
rect 36544 576438 36596 576444
rect 25504 575952 25556 575958
rect 25504 575894 25556 575900
rect 25516 423638 25544 575894
rect 36556 476066 36584 576438
rect 39304 576156 39356 576162
rect 39304 576098 39356 576104
rect 36544 476060 36596 476066
rect 36544 476002 36596 476008
rect 25504 423632 25556 423638
rect 25504 423574 25556 423580
rect 39316 411262 39344 576098
rect 47584 575748 47636 575754
rect 47584 575690 47636 575696
rect 39304 411256 39356 411262
rect 39304 411198 39356 411204
rect 47596 215286 47624 575690
rect 51724 575612 51776 575618
rect 51724 575554 51776 575560
rect 50344 575544 50396 575550
rect 50344 575486 50396 575492
rect 47584 215280 47636 215286
rect 47584 215222 47636 215228
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 21364 150408 21416 150414
rect 21364 150350 21416 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 50356 137970 50384 575486
rect 51736 164218 51764 575554
rect 53116 463690 53144 577594
rect 184388 577584 184440 577590
rect 184388 577526 184440 577532
rect 172428 577448 172480 577454
rect 172428 577390 172480 577396
rect 160836 577380 160888 577386
rect 160836 577322 160888 577328
rect 148968 577244 149020 577250
rect 148968 577186 149020 577192
rect 137284 577176 137336 577182
rect 137284 577118 137336 577124
rect 125324 577108 125376 577114
rect 125324 577050 125376 577056
rect 121368 577040 121420 577046
rect 113822 577008 113878 577017
rect 121368 576982 121420 576988
rect 113822 576943 113878 576952
rect 66904 576564 66956 576570
rect 66904 576506 66956 576512
rect 57244 576428 57296 576434
rect 57244 576370 57296 576376
rect 54484 575340 54536 575346
rect 54484 575282 54536 575288
rect 54496 516118 54524 575282
rect 54484 516112 54536 516118
rect 54484 516054 54536 516060
rect 53104 463684 53156 463690
rect 53104 463626 53156 463632
rect 57256 346390 57284 576370
rect 61384 576292 61436 576298
rect 61384 576234 61436 576240
rect 58624 574796 58676 574802
rect 58624 574738 58676 574744
rect 57244 346384 57296 346390
rect 57244 346326 57296 346332
rect 58636 241466 58664 574738
rect 61396 320142 61424 576234
rect 65524 576088 65576 576094
rect 65524 576030 65576 576036
rect 61384 320136 61436 320142
rect 61384 320078 61436 320084
rect 65536 267714 65564 576030
rect 66916 372570 66944 576506
rect 113836 575498 113864 576943
rect 121380 575770 121408 576982
rect 113528 575470 113864 575498
rect 121334 575742 121408 575770
rect 121334 575484 121362 575742
rect 125336 575498 125364 577050
rect 129464 575816 129516 575822
rect 129464 575758 129516 575764
rect 129476 575498 129504 575758
rect 133420 575680 133472 575686
rect 133420 575622 133472 575628
rect 133432 575498 133460 575622
rect 137296 575498 137324 577118
rect 141240 576020 141292 576026
rect 141240 575962 141292 575968
rect 141252 575498 141280 575962
rect 148980 575498 149008 577186
rect 153016 576360 153068 576366
rect 153016 576302 153068 576308
rect 153028 575498 153056 576302
rect 156972 575884 157024 575890
rect 156972 575826 157024 575832
rect 156984 575498 157012 575826
rect 160848 575498 160876 577322
rect 168748 577312 168800 577318
rect 168748 577254 168800 577260
rect 168760 575498 168788 577254
rect 172440 575498 172468 577390
rect 184400 575498 184428 577526
rect 211896 576768 211948 576774
rect 211896 576710 211948 576716
rect 199936 576700 199988 576706
rect 199936 576642 199988 576648
rect 188344 576632 188396 576638
rect 188344 576574 188396 576580
rect 188356 575498 188384 576574
rect 199948 575498 199976 576642
rect 211908 575498 211936 576710
rect 215772 575498 215800 578138
rect 219348 577516 219400 577522
rect 219348 577458 219400 577464
rect 219360 575770 219388 577458
rect 219360 575742 219434 575770
rect 125212 575470 125364 575498
rect 129168 575470 129504 575498
rect 133124 575470 133460 575498
rect 136988 575470 137324 575498
rect 140944 575470 141280 575498
rect 148764 575470 149008 575498
rect 152720 575470 153056 575498
rect 156676 575470 157012 575498
rect 160540 575470 160876 575498
rect 168452 575470 168788 575498
rect 172316 575470 172468 575498
rect 184092 575470 184428 575498
rect 188048 575470 188384 575498
rect 199824 575470 199976 575498
rect 211600 575470 211936 575498
rect 215464 575470 215800 575498
rect 219406 575484 219434 575742
rect 223500 575498 223528 616830
rect 227640 575498 227668 643078
rect 231768 630692 231820 630698
rect 231768 630634 231820 630640
rect 231780 576854 231808 630634
rect 235828 578202 235856 670754
rect 235356 578196 235408 578202
rect 235356 578138 235408 578144
rect 235816 578196 235868 578202
rect 235816 578138 235868 578144
rect 231596 576826 231808 576854
rect 231596 575498 231624 576826
rect 235368 575498 235396 578138
rect 235920 578134 235948 699654
rect 240048 696992 240100 696998
rect 240048 696934 240100 696940
rect 240060 578202 240088 696934
rect 244188 683256 244240 683262
rect 244188 683198 244240 683204
rect 244200 578202 244228 683198
rect 239312 578196 239364 578202
rect 239312 578138 239364 578144
rect 240048 578196 240100 578202
rect 240048 578138 240100 578144
rect 243268 578196 243320 578202
rect 243268 578138 243320 578144
rect 244188 578196 244240 578202
rect 244188 578138 244240 578144
rect 235908 578128 235960 578134
rect 235908 578070 235960 578076
rect 239324 575498 239352 578138
rect 243280 575498 243308 578138
rect 246948 577720 247000 577726
rect 246948 577662 247000 577668
rect 246960 575498 246988 577662
rect 251100 575498 251128 700538
rect 255228 700528 255280 700534
rect 255228 700470 255280 700476
rect 255240 576854 255268 700470
rect 263520 578202 263548 700810
rect 267568 699854 267596 702406
rect 267648 700800 267700 700806
rect 267648 700742 267700 700748
rect 267556 699848 267608 699854
rect 267556 699790 267608 699796
rect 267660 578202 267688 700742
rect 278688 700256 278740 700262
rect 278688 700198 278740 700204
rect 274548 700188 274600 700194
rect 274548 700130 274600 700136
rect 262864 578196 262916 578202
rect 262864 578138 262916 578144
rect 263508 578196 263560 578202
rect 263508 578138 263560 578144
rect 266820 578196 266872 578202
rect 266820 578138 266872 578144
rect 267648 578196 267700 578202
rect 267648 578138 267700 578144
rect 258908 577788 258960 577794
rect 258908 577730 258960 577736
rect 255148 576826 255268 576854
rect 255148 575498 255176 576826
rect 258920 575498 258948 577730
rect 262876 575498 262904 578138
rect 266832 575498 266860 578138
rect 270408 577924 270460 577930
rect 270408 577866 270460 577872
rect 270420 575770 270448 577866
rect 223284 575470 223528 575498
rect 227240 575470 227668 575498
rect 231196 575470 231624 575498
rect 235060 575470 235396 575498
rect 239016 575470 239352 575498
rect 242972 575470 243308 575498
rect 246836 575470 246988 575498
rect 250792 575470 251128 575498
rect 254748 575470 255176 575498
rect 258612 575470 258948 575498
rect 262568 575470 262904 575498
rect 266524 575470 266860 575498
rect 270374 575742 270448 575770
rect 270374 575484 270402 575742
rect 274560 575498 274588 700130
rect 278700 576854 278728 700198
rect 283852 699786 283880 703520
rect 291108 699984 291160 699990
rect 291108 699926 291160 699932
rect 286968 699916 287020 699922
rect 286968 699858 287020 699864
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 282460 578196 282512 578202
rect 282460 578138 282512 578144
rect 278608 576826 278728 576854
rect 278608 575498 278636 576826
rect 282472 575498 282500 578138
rect 286980 578066 287008 699858
rect 291120 578202 291148 699926
rect 296720 699848 296772 699854
rect 296720 699790 296772 699796
rect 296732 596174 296760 699790
rect 296732 596146 297496 596174
rect 290280 578196 290332 578202
rect 290280 578138 290332 578144
rect 291108 578196 291160 578202
rect 291108 578138 291160 578144
rect 293868 578196 293920 578202
rect 293868 578138 293920 578144
rect 286416 578060 286468 578066
rect 286416 578002 286468 578008
rect 286968 578060 287020 578066
rect 286968 578002 287020 578008
rect 286428 575498 286456 578002
rect 290292 575498 290320 578138
rect 293880 575770 293908 578138
rect 293880 575742 293954 575770
rect 274344 575470 274588 575498
rect 278208 575470 278636 575498
rect 282164 575470 282500 575498
rect 286120 575470 286456 575498
rect 289984 575470 290320 575498
rect 293926 575484 293954 575742
rect 297468 575498 297496 596146
rect 299492 578202 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 324320 701004 324372 701010
rect 324320 700946 324372 700952
rect 320180 700936 320232 700942
rect 320180 700878 320232 700884
rect 309140 700120 309192 700126
rect 309140 700062 309192 700068
rect 300860 699780 300912 699786
rect 300860 699722 300912 699728
rect 300872 596174 300900 699722
rect 309152 596174 309180 700062
rect 313280 700052 313332 700058
rect 313280 699994 313332 700000
rect 300872 596146 301360 596174
rect 309152 596146 309272 596174
rect 299480 578196 299532 578202
rect 299480 578138 299532 578144
rect 301332 575498 301360 596146
rect 305368 578128 305420 578134
rect 305368 578070 305420 578076
rect 305380 575498 305408 578070
rect 309244 575498 309272 596146
rect 313292 575498 313320 699994
rect 320192 596174 320220 700878
rect 324332 596174 324360 700946
rect 332520 699922 332548 703520
rect 336740 700732 336792 700738
rect 336740 700674 336792 700680
rect 332600 700664 332652 700670
rect 332600 700606 332652 700612
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 332612 596174 332640 700606
rect 320192 596146 320956 596174
rect 324332 596146 324912 596174
rect 332612 596146 332732 596174
rect 317420 577992 317472 577998
rect 317420 577934 317472 577940
rect 317432 575770 317460 577934
rect 317432 575742 317506 575770
rect 297468 575470 297896 575498
rect 301332 575470 301760 575498
rect 305380 575470 305716 575498
rect 309244 575470 309672 575498
rect 313292 575470 313536 575498
rect 317478 575484 317506 575742
rect 320928 575498 320956 596146
rect 324884 575498 324912 596146
rect 328920 577856 328972 577862
rect 328920 577798 328972 577804
rect 328932 575498 328960 577798
rect 332704 575498 332732 596146
rect 336752 575498 336780 700674
rect 340880 700460 340932 700466
rect 340880 700402 340932 700408
rect 340892 575498 340920 700402
rect 347780 700392 347832 700398
rect 347780 700334 347832 700340
rect 343640 700324 343692 700330
rect 343640 700266 343692 700272
rect 343652 596174 343680 700266
rect 347792 596174 347820 700334
rect 348804 699990 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 351920 683188 351972 683194
rect 351920 683130 351972 683136
rect 351932 596174 351960 683130
rect 360200 670744 360252 670750
rect 360200 670686 360252 670692
rect 356060 656940 356112 656946
rect 356060 656882 356112 656888
rect 356072 596174 356100 656882
rect 343652 596146 344508 596174
rect 347792 596146 348464 596174
rect 351932 596146 352420 596174
rect 356072 596146 356284 596174
rect 344480 575498 344508 596146
rect 348436 575498 348464 596146
rect 352392 575498 352420 596146
rect 356256 575498 356284 596146
rect 360212 575498 360240 670686
rect 364352 578066 364380 702406
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 364432 632120 364484 632126
rect 364432 632062 364484 632068
rect 364340 578060 364392 578066
rect 364340 578002 364392 578008
rect 364444 575498 364472 632062
rect 371240 618316 371292 618322
rect 371240 618258 371292 618264
rect 367100 605872 367152 605878
rect 367100 605814 367152 605820
rect 367112 596174 367140 605814
rect 371252 596174 371280 618258
rect 367112 596146 368060 596174
rect 371252 596146 372016 596174
rect 368032 575498 368060 596146
rect 371988 575498 372016 596146
rect 375840 579692 375892 579698
rect 375840 579634 375892 579640
rect 375852 575498 375880 579634
rect 429212 577930 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 430856 578332 430908 578338
rect 430856 578274 430908 578280
rect 429200 577924 429252 577930
rect 429200 577866 429252 577872
rect 407396 577652 407448 577658
rect 407396 577594 407448 577600
rect 399484 576496 399536 576502
rect 399484 576438 399536 576444
rect 387800 576224 387852 576230
rect 387800 576166 387852 576172
rect 387812 575498 387840 576166
rect 399496 575498 399524 576438
rect 407408 575498 407436 577594
rect 423036 576564 423088 576570
rect 423036 576506 423088 576512
rect 419080 576156 419132 576162
rect 419080 576098 419132 576104
rect 411260 575952 411312 575958
rect 411260 575894 411312 575900
rect 411272 575498 411300 575894
rect 419092 575498 419120 576098
rect 423048 575498 423076 576506
rect 426992 576428 427044 576434
rect 426992 576370 427044 576376
rect 427004 575498 427032 576370
rect 430868 575498 430896 578274
rect 442632 578264 442684 578270
rect 442632 578206 442684 578212
rect 434812 576292 434864 576298
rect 434812 576234 434864 576240
rect 434824 575498 434852 576234
rect 442644 575498 442672 578206
rect 494072 577794 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 494060 577788 494112 577794
rect 494060 577730 494112 577736
rect 558932 577726 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 558920 577720 558972 577726
rect 558920 577662 558972 577668
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 538864 577584 538916 577590
rect 538864 577526 538916 577532
rect 537484 577448 537536 577454
rect 537484 577390 537536 577396
rect 536104 577380 536156 577386
rect 536104 577322 536156 577328
rect 533344 577244 533396 577250
rect 533344 577186 533396 577192
rect 530584 577176 530636 577182
rect 477958 577144 478014 577153
rect 530584 577118 530636 577124
rect 477958 577079 478014 577088
rect 529204 577108 529256 577114
rect 454408 576972 454460 576978
rect 454408 576914 454460 576920
rect 446588 576088 446640 576094
rect 446588 576030 446640 576036
rect 446600 575498 446628 576030
rect 454420 575498 454448 576914
rect 466460 576904 466512 576910
rect 466460 576846 466512 576852
rect 466472 575770 466500 576846
rect 458686 575748 458738 575754
rect 466472 575742 466546 575770
rect 458686 575690 458738 575696
rect 320928 575470 321356 575498
rect 324884 575470 325312 575498
rect 328932 575470 329268 575498
rect 332704 575470 333132 575498
rect 336752 575470 337088 575498
rect 340892 575470 341044 575498
rect 344480 575470 344908 575498
rect 348436 575470 348864 575498
rect 352392 575470 352820 575498
rect 356256 575470 356684 575498
rect 360212 575470 360640 575498
rect 364444 575470 364596 575498
rect 368032 575470 368460 575498
rect 371988 575470 372416 575498
rect 375852 575470 376280 575498
rect 387812 575470 388056 575498
rect 399496 575470 399832 575498
rect 407408 575470 407744 575498
rect 411272 575470 411608 575498
rect 419092 575470 419428 575498
rect 423048 575470 423384 575498
rect 427004 575470 427340 575498
rect 430868 575470 431204 575498
rect 434824 575470 435160 575498
rect 442644 575470 442980 575498
rect 446600 575470 446936 575498
rect 454420 575470 454756 575498
rect 458698 575484 458726 575690
rect 466518 575484 466546 575742
rect 470140 575612 470192 575618
rect 470140 575554 470192 575560
rect 470152 575498 470180 575554
rect 474004 575544 474056 575550
rect 470152 575470 470488 575498
rect 477972 575498 478000 577079
rect 529204 577050 529256 577056
rect 526442 577008 526498 577017
rect 526442 576943 526498 576952
rect 519544 576768 519596 576774
rect 519544 576710 519596 576716
rect 518164 576700 518216 576706
rect 518164 576642 518216 576648
rect 516784 576632 516836 576638
rect 516784 576574 516836 576580
rect 474056 575492 474352 575498
rect 474004 575486 474352 575492
rect 474016 575470 474352 575486
rect 477972 575470 478308 575498
rect 395632 575346 395968 575362
rect 395620 575340 395968 575346
rect 395672 575334 395968 575340
rect 395620 575282 395672 575288
rect 207940 575272 207992 575278
rect 207644 575220 207940 575226
rect 207644 575214 207992 575220
rect 207644 575198 207980 575214
rect 379900 575210 380236 575226
rect 379888 575204 380236 575210
rect 379940 575198 380236 575204
rect 379888 575146 379940 575152
rect 203984 575136 204036 575142
rect 203688 575084 203984 575090
rect 203688 575078 204036 575084
rect 203688 575062 204024 575078
rect 383856 575074 384192 575090
rect 391860 575074 392012 575090
rect 403452 575074 403788 575090
rect 415412 575074 415564 575090
rect 438872 575074 439116 575090
rect 450556 575074 450892 575090
rect 462332 575074 462668 575090
rect 383844 575068 384192 575074
rect 383896 575062 384192 575068
rect 391848 575068 392012 575074
rect 383844 575010 383896 575016
rect 391900 575062 392012 575068
rect 403440 575068 403788 575074
rect 391848 575010 391900 575016
rect 403492 575062 403788 575068
rect 415400 575068 415564 575074
rect 403440 575010 403492 575016
rect 415452 575062 415564 575068
rect 438860 575068 439116 575074
rect 415400 575010 415452 575016
rect 438912 575062 439116 575068
rect 450544 575068 450892 575074
rect 438860 575010 438912 575016
rect 450596 575062 450892 575068
rect 462320 575068 462668 575074
rect 450544 575010 450596 575016
rect 462372 575062 462668 575068
rect 462320 575010 462372 575016
rect 195980 575000 196032 575006
rect 70214 574968 70270 574977
rect 73894 574968 73950 574977
rect 70270 574926 70380 574954
rect 70214 574903 70270 574912
rect 78402 574968 78458 574977
rect 73950 574926 74244 574954
rect 78200 574926 78402 574954
rect 73894 574903 73950 574912
rect 82358 574968 82414 574977
rect 82064 574926 82358 574954
rect 78402 574903 78458 574912
rect 86314 574968 86370 574977
rect 86020 574926 86314 574954
rect 82358 574903 82414 574912
rect 90270 574968 90326 574977
rect 89976 574926 90270 574954
rect 86314 574903 86370 574912
rect 90270 574903 90326 574912
rect 93674 574968 93730 574977
rect 97630 574968 97686 574977
rect 93730 574926 93840 574954
rect 93674 574903 93730 574912
rect 101954 574968 102010 574977
rect 97686 574926 97796 574954
rect 101752 574926 101954 574954
rect 97630 574903 97686 574912
rect 105910 574968 105966 574977
rect 105616 574926 105910 574954
rect 101954 574903 102010 574912
rect 109572 574938 109908 574954
rect 117392 574938 117728 574954
rect 144900 574938 145052 574954
rect 164496 574938 164832 574954
rect 176272 574938 176608 574954
rect 180136 574938 180472 574954
rect 191912 574938 192248 574954
rect 195868 574948 195980 574954
rect 195868 574942 196032 574948
rect 481914 574968 481970 574977
rect 109572 574932 109920 574938
rect 109572 574926 109868 574932
rect 105910 574903 105966 574912
rect 117392 574932 117740 574938
rect 117392 574926 117688 574932
rect 109868 574874 109920 574880
rect 144900 574932 145064 574938
rect 144900 574926 145012 574932
rect 117688 574874 117740 574880
rect 164496 574932 164844 574938
rect 164496 574926 164792 574932
rect 145012 574874 145064 574880
rect 176272 574932 176620 574938
rect 176272 574926 176568 574932
rect 164792 574874 164844 574880
rect 180136 574932 180484 574938
rect 180136 574926 180432 574932
rect 176568 574874 176620 574880
rect 191912 574932 192260 574938
rect 191912 574926 192208 574932
rect 180432 574874 180484 574880
rect 195868 574926 196020 574942
rect 485870 574968 485926 574977
rect 481970 574926 482264 574954
rect 481914 574903 481970 574912
rect 489918 574968 489974 574977
rect 485926 574926 486128 574954
rect 485870 574903 485926 574912
rect 493690 574968 493746 574977
rect 489974 574926 490084 574954
rect 489918 574903 489974 574912
rect 497554 574968 497610 574977
rect 493746 574926 494040 574954
rect 493690 574903 493746 574912
rect 501510 574968 501566 574977
rect 497610 574926 497904 574954
rect 497554 574903 497610 574912
rect 505466 574968 505522 574977
rect 501566 574926 501860 574954
rect 501510 574903 501566 574912
rect 509330 574968 509386 574977
rect 505522 574926 505816 574954
rect 505466 574903 505522 574912
rect 513930 574968 513986 574977
rect 509386 574926 509680 574954
rect 513636 574926 513930 574954
rect 509330 574903 509386 574912
rect 513930 574903 513986 574912
rect 192208 574874 192260 574880
rect 516796 458182 516824 576574
rect 518176 511970 518204 576642
rect 519556 564398 519584 576710
rect 525064 576360 525116 576366
rect 525064 576302 525116 576308
rect 522304 576020 522356 576026
rect 522304 575962 522356 575968
rect 520924 575816 520976 575822
rect 520924 575758 520976 575764
rect 519544 564392 519596 564398
rect 519544 564334 519596 564340
rect 518164 511964 518216 511970
rect 518164 511906 518216 511912
rect 516784 458176 516836 458182
rect 516784 458118 516836 458124
rect 66904 372564 66956 372570
rect 66904 372506 66956 372512
rect 65524 267708 65576 267714
rect 65524 267650 65576 267656
rect 58624 241460 58676 241466
rect 58624 241402 58676 241408
rect 520936 206990 520964 575758
rect 522316 245614 522344 575962
rect 525076 299470 525104 576302
rect 525064 299464 525116 299470
rect 525064 299406 525116 299412
rect 522304 245608 522356 245614
rect 522304 245550 522356 245556
rect 520924 206984 520976 206990
rect 520924 206926 520976 206932
rect 51724 164212 51776 164218
rect 51724 164154 51776 164160
rect 526456 139398 526484 576943
rect 529216 179382 529244 577050
rect 530596 219434 530624 577118
rect 533356 259418 533384 577186
rect 536116 313274 536144 577322
rect 537496 365702 537524 577390
rect 538876 419490 538904 577526
rect 580184 577522 580212 577623
rect 580172 577516 580224 577522
rect 580172 577458 580224 577464
rect 551284 577312 551336 577318
rect 551284 577254 551336 577260
rect 543004 577040 543056 577046
rect 543004 576982 543056 576988
rect 540244 574320 540296 574326
rect 540244 574262 540296 574268
rect 538864 419484 538916 419490
rect 538864 419426 538916 419432
rect 537484 365696 537536 365702
rect 537484 365638 537536 365644
rect 536104 313268 536156 313274
rect 536104 313210 536156 313216
rect 533344 259412 533396 259418
rect 533344 259354 533396 259360
rect 530584 219428 530636 219434
rect 530584 219370 530636 219376
rect 529204 179376 529256 179382
rect 529204 179318 529256 179324
rect 540256 153202 540284 574262
rect 543016 193186 543044 576982
rect 548524 575884 548576 575890
rect 548524 575826 548576 575832
rect 544384 575680 544436 575686
rect 544384 575622 544436 575628
rect 544396 233238 544424 575622
rect 547144 574592 547196 574598
rect 547144 574534 547196 574540
rect 547156 273222 547184 574534
rect 548536 325650 548564 575826
rect 551296 379506 551324 577254
rect 580816 575272 580868 575278
rect 580816 575214 580868 575220
rect 580632 575000 580684 575006
rect 580632 574942 580684 574948
rect 580540 574660 580592 574666
rect 580540 574602 580592 574608
rect 580448 574524 580500 574530
rect 580448 574466 580500 574472
rect 580356 574388 580408 574394
rect 580356 574330 580408 574336
rect 580264 574116 580316 574122
rect 580264 574058 580316 574064
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 579712 419484 579764 419490
rect 579712 419426 579764 419432
rect 579724 418305 579752 419426
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 551284 379500 551336 379506
rect 551284 379442 551336 379448
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 579988 365696 580040 365702
rect 579988 365638 580040 365644
rect 580000 365129 580028 365638
rect 579986 365120 580042 365129
rect 579986 365055 580042 365064
rect 548524 325644 548576 325650
rect 548524 325586 548576 325592
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 547144 273216 547196 273222
rect 547144 273158 547196 273164
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 544384 233232 544436 233238
rect 544384 233174 544436 233180
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 579896 219428 579948 219434
rect 579896 219370 579948 219376
rect 579908 219065 579936 219370
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 543004 193180 543056 193186
rect 543004 193122 543056 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 579988 179376 580040 179382
rect 579988 179318 580040 179324
rect 580000 179217 580028 179318
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580276 165889 580304 574058
rect 580368 351937 580396 574330
rect 580460 404977 580488 574466
rect 580552 431633 580580 574602
rect 580644 471481 580672 574942
rect 580724 574932 580776 574938
rect 580724 574874 580776 574880
rect 580736 484673 580764 574874
rect 580828 524521 580856 575214
rect 580908 575136 580960 575142
rect 580908 575078 580960 575084
rect 580920 537849 580948 575078
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580814 524512 580870 524521
rect 580814 524447 580870 524456
rect 580722 484664 580778 484673
rect 580722 484599 580778 484608
rect 580630 471472 580686 471481
rect 580630 471407 580686 471416
rect 580538 431624 580594 431633
rect 580538 431559 580594 431568
rect 580446 404968 580502 404977
rect 580446 404903 580502 404912
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580262 165880 580318 165889
rect 580262 165815 580318 165824
rect 540244 153196 540296 153202
rect 540244 153138 540296 153144
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 526444 139392 526496 139398
rect 580172 139392 580224 139398
rect 526444 139334 526496 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 50344 137964 50396 137970
rect 50344 137906 50396 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 67652 128438 68816 128466
rect 64788 126948 64840 126954
rect 64788 126890 64840 126896
rect 56508 126880 56560 126886
rect 56508 126822 56560 126828
rect 29644 126744 29696 126750
rect 29644 126686 29696 126692
rect 14464 126676 14516 126682
rect 14464 126618 14516 126624
rect 7564 126336 7616 126342
rect 7564 126278 7616 126284
rect 4804 124908 4856 124914
rect 4804 124850 4856 124856
rect 3422 111752 3478 111761
rect 3422 111687 3478 111696
rect 3436 110673 3464 111687
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3516 89004 3568 89010
rect 3516 88946 3568 88952
rect 3422 85504 3478 85513
rect 3422 85439 3478 85448
rect 3436 84697 3464 85439
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3528 84194 3556 88946
rect 3436 84166 3556 84194
rect 3238 59256 3294 59265
rect 3238 59191 3294 59200
rect 3252 58585 3280 59191
rect 3238 58576 3294 58585
rect 3238 58511 3294 58520
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 572 3188 624 3194
rect 572 3130 624 3136
rect 584 480 612 3130
rect 1688 480 1716 3402
rect 2884 480 2912 3470
rect 3436 3194 3464 84166
rect 3514 33144 3570 33153
rect 3514 33079 3570 33088
rect 3528 32473 3556 33079
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3514 20632 3570 20641
rect 3514 20567 3570 20576
rect 3528 19417 3556 20567
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 4080 480 4108 4762
rect 4816 3534 4844 124850
rect 7576 3874 7604 126278
rect 11704 126268 11756 126274
rect 11704 126210 11756 126216
rect 7656 4888 7708 4894
rect 7656 4830 7708 4836
rect 5264 3868 5316 3874
rect 5264 3810 5316 3816
rect 7564 3868 7616 3874
rect 7564 3810 7616 3816
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5276 480 5304 3810
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6472 480 6500 3538
rect 7668 480 7696 4830
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 480 8800 3334
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9968 480 9996 2994
rect 11164 480 11192 3402
rect 11716 3058 11744 126210
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 12360 480 12388 5034
rect 14476 3602 14504 126618
rect 22744 126608 22796 126614
rect 22744 126550 22796 126556
rect 21364 126472 21416 126478
rect 21364 126414 21416 126420
rect 17224 126404 17276 126410
rect 17224 126346 17276 126352
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 14740 3800 14792 3806
rect 14740 3742 14792 3748
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 13542 3360 13598 3369
rect 13542 3295 13598 3304
rect 13556 480 13584 3295
rect 14752 480 14780 3742
rect 15934 3496 15990 3505
rect 15934 3431 15990 3440
rect 15948 480 15976 3431
rect 17052 480 17080 3878
rect 17236 3806 17264 126346
rect 18604 125248 18656 125254
rect 18604 125190 18656 125196
rect 17224 3800 17276 3806
rect 17224 3742 17276 3748
rect 18616 3602 18644 125190
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 480 18276 3470
rect 19444 480 19472 3606
rect 21376 3534 21404 126414
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20640 480 20668 2994
rect 21836 480 21864 3946
rect 22756 3058 22784 126550
rect 25504 126540 25556 126546
rect 25504 126482 25556 126488
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 23032 480 23060 3538
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24228 480 24256 3470
rect 25332 480 25360 3674
rect 25516 3534 25544 126482
rect 26516 4956 26568 4962
rect 26516 4898 26568 4904
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 26528 480 26556 4898
rect 29656 3670 29684 126686
rect 50344 125928 50396 125934
rect 50344 125870 50396 125876
rect 39304 125520 39356 125526
rect 39304 125462 39356 125468
rect 32404 125452 32456 125458
rect 32404 125394 32456 125400
rect 30104 5024 30156 5030
rect 30104 4966 30156 4972
rect 27712 3664 27764 3670
rect 27712 3606 27764 3612
rect 29644 3664 29696 3670
rect 29644 3606 29696 3612
rect 27724 480 27752 3606
rect 28908 3324 28960 3330
rect 28908 3266 28960 3272
rect 28920 480 28948 3266
rect 30116 480 30144 4966
rect 32416 3942 32444 125394
rect 33784 125316 33836 125322
rect 33784 125258 33836 125264
rect 33796 4010 33824 125258
rect 37188 123548 37240 123554
rect 37188 123490 37240 123496
rect 35164 123480 35216 123486
rect 35164 123422 35216 123428
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 33784 4004 33836 4010
rect 33784 3946 33836 3952
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 31300 3868 31352 3874
rect 31300 3810 31352 3816
rect 31312 480 31340 3810
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32416 480 32444 3742
rect 33600 3664 33652 3670
rect 33600 3606 33652 3612
rect 33612 480 33640 3606
rect 34808 480 34836 4082
rect 35176 3670 35204 123422
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 35164 3664 35216 3670
rect 35164 3606 35216 3612
rect 36004 480 36032 3878
rect 37200 480 37228 123490
rect 38384 4072 38436 4078
rect 38384 4014 38436 4020
rect 38396 480 38424 4014
rect 39316 3398 39344 125462
rect 48228 124976 48280 124982
rect 48228 124918 48280 124924
rect 41328 123616 41380 123622
rect 41328 123558 41380 123564
rect 39580 4004 39632 4010
rect 39580 3946 39632 3952
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 39592 480 39620 3946
rect 41340 3398 41368 123558
rect 44272 7608 44324 7614
rect 44272 7550 44324 7556
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 40696 480 40724 3334
rect 43076 3324 43128 3330
rect 43076 3266 43128 3272
rect 41880 3256 41932 3262
rect 41880 3198 41932 3204
rect 41892 480 41920 3198
rect 43088 480 43116 3266
rect 44284 480 44312 7550
rect 48240 6914 48268 124918
rect 47872 6886 48268 6914
rect 45468 3188 45520 3194
rect 45468 3130 45520 3136
rect 45480 480 45508 3130
rect 46664 3052 46716 3058
rect 46664 2994 46716 3000
rect 46676 480 46704 2994
rect 47872 480 47900 6886
rect 50356 5030 50384 125870
rect 53104 125860 53156 125866
rect 53104 125802 53156 125808
rect 52368 125044 52420 125050
rect 52368 124986 52420 124992
rect 50344 5024 50396 5030
rect 50344 4966 50396 4972
rect 50896 4752 50948 4758
rect 50896 4694 50948 4700
rect 50160 3120 50212 3126
rect 50160 3062 50212 3068
rect 48964 2848 49016 2854
rect 48964 2790 49016 2796
rect 48976 480 49004 2790
rect 50172 480 50200 3062
rect 50908 2854 50936 4694
rect 52380 3398 52408 124986
rect 53116 5098 53144 125802
rect 55128 125112 55180 125118
rect 55128 125054 55180 125060
rect 55140 6914 55168 125054
rect 54956 6886 55168 6914
rect 53104 5092 53156 5098
rect 53104 5034 53156 5040
rect 52552 5024 52604 5030
rect 52552 4966 52604 4972
rect 51356 3392 51408 3398
rect 51356 3334 51408 3340
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 50896 2848 50948 2854
rect 50896 2790 50948 2796
rect 51368 480 51396 3334
rect 52564 480 52592 4966
rect 53748 3052 53800 3058
rect 53748 2994 53800 3000
rect 53760 480 53788 2994
rect 54956 480 54984 6886
rect 56520 2990 56548 126822
rect 57888 126812 57940 126818
rect 57888 126754 57940 126760
rect 57900 2990 57928 126754
rect 63408 126200 63460 126206
rect 63408 126142 63460 126148
rect 58624 125996 58676 126002
rect 58624 125938 58676 125944
rect 58636 7614 58664 125938
rect 62028 125180 62080 125186
rect 62028 125122 62080 125128
rect 58624 7608 58676 7614
rect 58624 7550 58676 7556
rect 58440 7540 58492 7546
rect 58440 7482 58492 7488
rect 56048 2984 56100 2990
rect 56048 2926 56100 2932
rect 56508 2984 56560 2990
rect 56508 2926 56560 2932
rect 57244 2984 57296 2990
rect 57244 2926 57296 2932
rect 57888 2984 57940 2990
rect 57888 2926 57940 2932
rect 56060 480 56088 2926
rect 57256 480 57284 2926
rect 58452 480 58480 7482
rect 59636 5160 59688 5166
rect 59636 5102 59688 5108
rect 59648 480 59676 5102
rect 60832 2916 60884 2922
rect 60832 2858 60884 2864
rect 60844 480 60872 2858
rect 62040 480 62068 125122
rect 63420 6914 63448 126142
rect 63236 6886 63448 6914
rect 63236 480 63264 6886
rect 64800 2990 64828 126890
rect 66168 125384 66220 125390
rect 66168 125326 66220 125332
rect 66180 2990 66208 125326
rect 67652 89010 67680 128438
rect 69630 128194 69658 128452
rect 70550 128330 70578 128452
rect 69584 128166 69658 128194
rect 70504 128302 70578 128330
rect 68284 126064 68336 126070
rect 68284 126006 68336 126012
rect 67640 89004 67692 89010
rect 67640 88946 67692 88952
rect 68296 5166 68324 126006
rect 69584 125254 69612 128166
rect 70216 126132 70268 126138
rect 70216 126074 70268 126080
rect 69572 125248 69624 125254
rect 69572 125190 69624 125196
rect 70228 16574 70256 126074
rect 70504 124914 70532 128302
rect 71470 128194 71498 128452
rect 72390 128194 72418 128452
rect 73310 128194 73338 128452
rect 74230 128194 74258 128452
rect 75150 128194 75178 128452
rect 75978 128194 76006 128452
rect 76898 128194 76926 128452
rect 77818 128194 77846 128452
rect 70688 128166 71498 128194
rect 72344 128166 72418 128194
rect 73264 128166 73338 128194
rect 74184 128166 74258 128194
rect 75104 128166 75178 128194
rect 75932 128166 76006 128194
rect 76116 128166 76926 128194
rect 77772 128166 77846 128194
rect 78738 128194 78766 128452
rect 79658 128194 79686 128452
rect 80578 128194 80606 128452
rect 81498 128194 81526 128452
rect 82326 128194 82354 128452
rect 83246 128194 83274 128452
rect 84166 128194 84194 128452
rect 85086 128194 85114 128452
rect 86006 128194 86034 128452
rect 86926 128194 86954 128452
rect 87846 128194 87874 128452
rect 88674 128194 88702 128452
rect 89594 128194 89622 128452
rect 90514 128194 90542 128452
rect 91434 128330 91462 128452
rect 78738 128166 78812 128194
rect 70492 124908 70544 124914
rect 70492 124850 70544 124856
rect 70688 122834 70716 128166
rect 72344 126342 72372 128166
rect 73264 126682 73292 128166
rect 73252 126676 73304 126682
rect 73252 126618 73304 126624
rect 72332 126336 72384 126342
rect 72332 126278 72384 126284
rect 74184 125662 74212 128166
rect 72424 125656 72476 125662
rect 72424 125598 72476 125604
rect 74172 125656 74224 125662
rect 74172 125598 74224 125604
rect 70412 122806 70716 122834
rect 70228 16546 70348 16574
rect 68284 5160 68336 5166
rect 68284 5102 68336 5108
rect 69112 5160 69164 5166
rect 69112 5102 69164 5108
rect 64328 2984 64380 2990
rect 64328 2926 64380 2932
rect 64788 2984 64840 2990
rect 64788 2926 64840 2932
rect 65524 2984 65576 2990
rect 65524 2926 65576 2932
rect 66168 2984 66220 2990
rect 66168 2926 66220 2932
rect 64340 480 64368 2926
rect 65536 480 65564 2926
rect 66720 2848 66772 2854
rect 66720 2790 66772 2796
rect 67916 2848 67968 2854
rect 67916 2790 67968 2796
rect 66732 480 66760 2790
rect 67928 480 67956 2790
rect 69124 480 69152 5102
rect 70320 480 70348 16546
rect 70412 4826 70440 122806
rect 72436 4894 72464 125598
rect 75104 125526 75132 128166
rect 75828 126336 75880 126342
rect 75828 126278 75880 126284
rect 75092 125520 75144 125526
rect 75092 125462 75144 125468
rect 72424 4888 72476 4894
rect 72424 4830 72476 4836
rect 70400 4820 70452 4826
rect 70400 4762 70452 4768
rect 72608 4820 72660 4826
rect 72608 4762 72660 4768
rect 71502 3632 71558 3641
rect 71502 3567 71558 3576
rect 71516 480 71544 3567
rect 72620 480 72648 4762
rect 73802 3768 73858 3777
rect 73802 3703 73858 3712
rect 73816 480 73844 3703
rect 75840 3466 75868 126278
rect 75932 126274 75960 128166
rect 75920 126268 75972 126274
rect 75920 126210 75972 126216
rect 76116 3602 76144 128166
rect 77772 125866 77800 128166
rect 78496 126676 78548 126682
rect 78496 126618 78548 126624
rect 77760 125860 77812 125866
rect 77760 125802 77812 125808
rect 77116 10328 77168 10334
rect 77116 10270 77168 10276
rect 76104 3596 76156 3602
rect 76104 3538 76156 3544
rect 77128 3466 77156 10270
rect 78508 3466 78536 126618
rect 78588 126268 78640 126274
rect 78588 126210 78640 126216
rect 75000 3460 75052 3466
rect 75000 3402 75052 3408
rect 75828 3460 75880 3466
rect 75828 3402 75880 3408
rect 76196 3460 76248 3466
rect 76196 3402 76248 3408
rect 77116 3460 77168 3466
rect 77116 3402 77168 3408
rect 77392 3460 77444 3466
rect 77392 3402 77444 3408
rect 78496 3460 78548 3466
rect 78496 3402 78548 3408
rect 75012 480 75040 3402
rect 76208 480 76236 3402
rect 77404 480 77432 3402
rect 78600 480 78628 126210
rect 78784 3233 78812 128166
rect 79612 128166 79686 128194
rect 80072 128166 80606 128194
rect 81452 128166 81526 128194
rect 82280 128166 82354 128194
rect 82924 128166 83274 128194
rect 84120 128166 84194 128194
rect 85040 128166 85114 128194
rect 85776 128166 86034 128194
rect 86880 128166 86954 128194
rect 87064 128166 87874 128194
rect 88444 128166 88702 128194
rect 89548 128166 89622 128194
rect 89732 128166 90542 128194
rect 91204 128302 91462 128330
rect 79612 126410 79640 128166
rect 79600 126404 79652 126410
rect 79600 126346 79652 126352
rect 79692 7676 79744 7682
rect 79692 7618 79744 7624
rect 78770 3224 78826 3233
rect 78770 3159 78826 3168
rect 79704 480 79732 7618
rect 80072 3369 80100 128166
rect 81452 125458 81480 128166
rect 82280 126478 82308 128166
rect 82268 126472 82320 126478
rect 82268 126414 82320 126420
rect 81440 125452 81492 125458
rect 81440 125394 81492 125400
rect 82924 3602 82952 128166
rect 84120 126614 84148 128166
rect 84108 126608 84160 126614
rect 84108 126550 84160 126556
rect 85040 125322 85068 128166
rect 85028 125316 85080 125322
rect 85028 125258 85080 125264
rect 84108 49020 84160 49026
rect 84108 48962 84160 48968
rect 82912 3596 82964 3602
rect 82912 3538 82964 3544
rect 80886 3496 80942 3505
rect 84120 3466 84148 48962
rect 84476 3732 84528 3738
rect 84476 3674 84528 3680
rect 80886 3431 80942 3440
rect 83280 3460 83332 3466
rect 80058 3360 80114 3369
rect 80058 3295 80114 3304
rect 80900 480 80928 3431
rect 83280 3402 83332 3408
rect 84108 3460 84160 3466
rect 84108 3402 84160 3408
rect 82082 3360 82138 3369
rect 82082 3295 82138 3304
rect 82096 480 82124 3295
rect 83292 480 83320 3402
rect 84488 480 84516 3674
rect 85776 3534 85804 128166
rect 86880 126546 86908 128166
rect 86868 126540 86920 126546
rect 86868 126482 86920 126488
rect 86868 15904 86920 15910
rect 86868 15846 86920 15852
rect 85764 3528 85816 3534
rect 85764 3470 85816 3476
rect 85672 3460 85724 3466
rect 85672 3402 85724 3408
rect 85684 480 85712 3402
rect 86880 480 86908 15846
rect 87064 3602 87092 128166
rect 88248 126540 88300 126546
rect 88248 126482 88300 126488
rect 88260 123622 88288 126482
rect 88248 123616 88300 123622
rect 88248 123558 88300 123564
rect 88444 4962 88472 128166
rect 89548 126750 89576 128166
rect 89536 126744 89588 126750
rect 89536 126686 89588 126692
rect 88984 126472 89036 126478
rect 88984 126414 89036 126420
rect 88996 123554 89024 126414
rect 88984 123548 89036 123554
rect 88984 123490 89036 123496
rect 88432 4956 88484 4962
rect 88432 4898 88484 4904
rect 87052 3596 87104 3602
rect 87052 3538 87104 3544
rect 87972 3596 88024 3602
rect 87972 3538 88024 3544
rect 87984 480 88012 3538
rect 89732 3534 89760 128166
rect 91204 125934 91232 128302
rect 92354 128194 92382 128452
rect 93274 128194 93302 128452
rect 91296 128166 92382 128194
rect 92492 128166 93302 128194
rect 93860 128240 93912 128246
rect 94194 128194 94222 128452
rect 95022 128246 95050 128452
rect 93860 128182 93912 128188
rect 91192 125928 91244 125934
rect 91192 125870 91244 125876
rect 91008 18624 91060 18630
rect 91008 18566 91060 18572
rect 91020 3534 91048 18566
rect 91296 3874 91324 128166
rect 91284 3868 91336 3874
rect 91284 3810 91336 3816
rect 91560 3868 91612 3874
rect 91560 3810 91612 3816
rect 89720 3528 89772 3534
rect 89720 3470 89772 3476
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 89168 3460 89220 3466
rect 89168 3402 89220 3408
rect 89180 480 89208 3402
rect 90376 480 90404 3470
rect 91572 480 91600 3810
rect 92492 3806 92520 128166
rect 93768 126404 93820 126410
rect 93768 126346 93820 126352
rect 93780 3806 93808 126346
rect 93872 3942 93900 128182
rect 94148 128166 94222 128194
rect 95010 128240 95062 128246
rect 95942 128194 95970 128452
rect 96862 128330 96890 128452
rect 95010 128182 95062 128188
rect 95252 128166 95970 128194
rect 96632 128302 96890 128330
rect 94148 123486 94176 128166
rect 94136 123480 94188 123486
rect 94136 123422 94188 123428
rect 93952 4956 94004 4962
rect 93952 4898 94004 4904
rect 93860 3936 93912 3942
rect 93860 3878 93912 3884
rect 92480 3800 92532 3806
rect 92480 3742 92532 3748
rect 92756 3800 92808 3806
rect 92756 3742 92808 3748
rect 93768 3800 93820 3806
rect 93768 3742 93820 3748
rect 92768 480 92796 3742
rect 93964 480 93992 4898
rect 95148 3800 95200 3806
rect 95148 3742 95200 3748
rect 95160 480 95188 3742
rect 95252 3670 95280 128166
rect 96632 126478 96660 128302
rect 97782 128194 97810 128452
rect 98702 128194 98730 128452
rect 99622 128194 99650 128452
rect 100542 128194 100570 128452
rect 101370 128194 101398 128452
rect 102290 128194 102318 128452
rect 103210 128194 103238 128452
rect 104130 128194 104158 128452
rect 105050 128330 105078 128452
rect 96724 128166 97810 128194
rect 98012 128166 98730 128194
rect 99576 128166 99650 128194
rect 99760 128166 100570 128194
rect 100864 128166 101398 128194
rect 102244 128166 102318 128194
rect 102428 128166 103238 128194
rect 103624 128166 104158 128194
rect 105004 128302 105078 128330
rect 96620 126472 96672 126478
rect 96620 126414 96672 126420
rect 96724 4078 96752 128166
rect 97448 4888 97500 4894
rect 97448 4830 97500 4836
rect 96712 4072 96764 4078
rect 96712 4014 96764 4020
rect 95240 3664 95292 3670
rect 95240 3606 95292 3612
rect 96252 3324 96304 3330
rect 96252 3266 96304 3272
rect 96264 480 96292 3266
rect 97460 480 97488 4830
rect 98012 4010 98040 128166
rect 99576 126546 99604 128166
rect 99564 126540 99616 126546
rect 99564 126482 99616 126488
rect 99288 126472 99340 126478
rect 99288 126414 99340 126420
rect 98000 4004 98052 4010
rect 98000 3946 98052 3952
rect 99300 3670 99328 126414
rect 99760 4146 99788 128166
rect 99748 4140 99800 4146
rect 99748 4082 99800 4088
rect 99840 3936 99892 3942
rect 99840 3878 99892 3884
rect 98644 3664 98696 3670
rect 98644 3606 98696 3612
rect 99288 3664 99340 3670
rect 99288 3606 99340 3612
rect 98656 480 98684 3606
rect 99852 480 99880 3878
rect 100864 3194 100892 128166
rect 102244 126002 102272 128166
rect 102232 125996 102284 126002
rect 102232 125938 102284 125944
rect 102048 26920 102100 26926
rect 102048 26862 102100 26868
rect 102060 3670 102088 26862
rect 102232 4140 102284 4146
rect 102232 4082 102284 4088
rect 101036 3664 101088 3670
rect 101036 3606 101088 3612
rect 102048 3664 102100 3670
rect 102048 3606 102100 3612
rect 100852 3188 100904 3194
rect 100852 3130 100904 3136
rect 101048 480 101076 3606
rect 102244 480 102272 4082
rect 102428 4010 102456 128166
rect 103336 4072 103388 4078
rect 103336 4014 103388 4020
rect 102416 4004 102468 4010
rect 102416 3946 102468 3952
rect 103348 480 103376 4014
rect 103624 3398 103652 128166
rect 104808 126540 104860 126546
rect 104808 126482 104860 126488
rect 104820 6914 104848 126482
rect 105004 124982 105032 128302
rect 105970 128194 105998 128452
rect 106890 128194 106918 128452
rect 107718 128194 107746 128452
rect 108638 128194 108666 128452
rect 109558 128194 109586 128452
rect 110478 128194 110506 128452
rect 111398 128194 111426 128452
rect 112318 128194 112346 128452
rect 113238 128194 113266 128452
rect 114158 128194 114186 128452
rect 114986 128194 115014 128452
rect 115906 128194 115934 128452
rect 116826 128194 116854 128452
rect 117746 128194 117774 128452
rect 118666 128194 118694 128452
rect 119586 128194 119614 128452
rect 120506 128194 120534 128452
rect 121334 128194 121362 128452
rect 122254 128194 122282 128452
rect 123174 128194 123202 128452
rect 124094 128194 124122 128452
rect 125014 128194 125042 128452
rect 105188 128166 105998 128194
rect 106292 128166 106918 128194
rect 107672 128166 107746 128194
rect 107856 128166 108666 128194
rect 109052 128166 109586 128194
rect 110432 128166 110506 128194
rect 111352 128166 111426 128194
rect 112272 128166 112346 128194
rect 113192 128166 113266 128194
rect 114112 128166 114186 128194
rect 114756 128166 115014 128194
rect 115860 128166 115934 128194
rect 116780 128166 116854 128194
rect 117700 128166 117774 128194
rect 118620 128166 118694 128194
rect 118988 128166 119614 128194
rect 120276 128166 120534 128194
rect 121288 128166 121362 128194
rect 122208 128166 122282 128194
rect 122944 128166 123202 128194
rect 124048 128166 124122 128194
rect 124232 128166 125042 128194
rect 125692 128240 125744 128246
rect 125934 128194 125962 128452
rect 126854 128246 126882 128452
rect 125692 128182 125744 128188
rect 104992 124976 105044 124982
rect 104992 124918 105044 124924
rect 105188 122834 105216 128166
rect 104544 6886 104848 6914
rect 104912 122806 105216 122834
rect 103612 3392 103664 3398
rect 103612 3334 103664 3340
rect 104544 480 104572 6886
rect 104912 5030 104940 122806
rect 104900 5024 104952 5030
rect 104900 4966 104952 4972
rect 105728 4004 105780 4010
rect 105728 3946 105780 3952
rect 105740 480 105768 3946
rect 106292 3126 106320 128166
rect 107672 125050 107700 128166
rect 107660 125044 107712 125050
rect 107660 124986 107712 124992
rect 107856 5098 107884 128166
rect 107844 5092 107896 5098
rect 107844 5034 107896 5040
rect 108120 5024 108172 5030
rect 108120 4966 108172 4972
rect 106924 3324 106976 3330
rect 106924 3266 106976 3272
rect 106280 3120 106332 3126
rect 106280 3062 106332 3068
rect 106936 480 106964 3266
rect 108132 480 108160 4966
rect 109052 3058 109080 128166
rect 110432 125118 110460 128166
rect 111352 126886 111380 128166
rect 111340 126880 111392 126886
rect 111340 126822 111392 126828
rect 112272 126818 112300 128166
rect 113192 126886 113220 128166
rect 112536 126880 112588 126886
rect 112536 126822 112588 126828
rect 113180 126880 113232 126886
rect 113180 126822 113232 126828
rect 112260 126812 112312 126818
rect 112260 126754 112312 126760
rect 112444 126812 112496 126818
rect 112444 126754 112496 126760
rect 111708 126608 111760 126614
rect 111708 126550 111760 126556
rect 110420 125112 110472 125118
rect 110420 125054 110472 125060
rect 111616 124908 111668 124914
rect 111616 124850 111668 124856
rect 110512 3392 110564 3398
rect 110512 3334 110564 3340
rect 109316 3256 109368 3262
rect 109316 3198 109368 3204
rect 109040 3052 109092 3058
rect 109040 2994 109092 3000
rect 109328 480 109356 3198
rect 110524 480 110552 3334
rect 111628 480 111656 124850
rect 111720 3398 111748 126550
rect 112456 5166 112484 126754
rect 112548 7614 112576 126822
rect 114112 126070 114140 128166
rect 114100 126064 114152 126070
rect 114100 126006 114152 126012
rect 112536 7608 112588 7614
rect 112536 7550 112588 7556
rect 112444 5160 112496 5166
rect 112444 5102 112496 5108
rect 111708 3392 111760 3398
rect 111708 3334 111760 3340
rect 112812 3392 112864 3398
rect 112812 3334 112864 3340
rect 112824 480 112852 3334
rect 114008 3120 114060 3126
rect 114008 3062 114060 3068
rect 114020 480 114048 3062
rect 114756 2990 114784 128166
rect 115860 125186 115888 128166
rect 116780 126206 116808 128166
rect 117700 126954 117728 128166
rect 117688 126948 117740 126954
rect 117688 126890 117740 126896
rect 117228 126744 117280 126750
rect 117228 126686 117280 126692
rect 116768 126200 116820 126206
rect 116768 126142 116820 126148
rect 115848 125180 115900 125186
rect 115848 125122 115900 125128
rect 115848 11756 115900 11762
rect 115848 11698 115900 11704
rect 115860 3194 115888 11698
rect 117240 3194 117268 126686
rect 118620 125662 118648 128166
rect 118608 125656 118660 125662
rect 118608 125598 118660 125604
rect 115204 3188 115256 3194
rect 115204 3130 115256 3136
rect 115848 3188 115900 3194
rect 115848 3130 115900 3136
rect 116400 3188 116452 3194
rect 116400 3130 116452 3136
rect 117228 3188 117280 3194
rect 117228 3130 117280 3136
rect 114744 2984 114796 2990
rect 114744 2926 114796 2932
rect 115216 480 115244 3130
rect 116412 480 116440 3130
rect 117596 3120 117648 3126
rect 117596 3062 117648 3068
rect 117608 480 117636 3062
rect 118988 2922 119016 128166
rect 120276 3058 120304 128166
rect 121288 126818 121316 128166
rect 122104 126948 122156 126954
rect 122104 126890 122156 126896
rect 121276 126812 121328 126818
rect 121276 126754 121328 126760
rect 122116 4826 122144 126890
rect 122208 126138 122236 128166
rect 122196 126132 122248 126138
rect 122196 126074 122248 126080
rect 122104 4820 122156 4826
rect 122104 4762 122156 4768
rect 122944 3641 122972 128166
rect 124048 126954 124076 128166
rect 124036 126948 124088 126954
rect 124036 126890 124088 126896
rect 124128 126812 124180 126818
rect 124128 126754 124180 126760
rect 123300 3732 123352 3738
rect 123300 3674 123352 3680
rect 123312 3641 123340 3674
rect 122930 3632 122986 3641
rect 122930 3567 122986 3576
rect 123298 3632 123354 3641
rect 123298 3567 123354 3576
rect 124140 3466 124168 126754
rect 124232 3777 124260 128166
rect 125508 126948 125560 126954
rect 125508 126890 125560 126896
rect 125520 6914 125548 126890
rect 125704 10334 125732 128182
rect 125888 128166 125962 128194
rect 126842 128240 126894 128246
rect 127682 128194 127710 128452
rect 128602 128330 128630 128452
rect 126842 128182 126894 128188
rect 127636 128166 127710 128194
rect 128372 128302 128630 128330
rect 125888 126342 125916 128166
rect 126244 126880 126296 126886
rect 126244 126822 126296 126828
rect 125876 126336 125928 126342
rect 125876 126278 125928 126284
rect 126256 26926 126284 126822
rect 127636 126682 127664 128166
rect 127624 126676 127676 126682
rect 127624 126618 127676 126624
rect 128372 126274 128400 128302
rect 129522 128194 129550 128452
rect 130442 128194 130470 128452
rect 131362 128194 131390 128452
rect 132282 128194 132310 128452
rect 133202 128194 133230 128452
rect 134030 128194 134058 128452
rect 134950 128194 134978 128452
rect 135870 128194 135898 128452
rect 136790 128194 136818 128452
rect 137710 128194 137738 128452
rect 138630 128194 138658 128452
rect 139550 128194 139578 128452
rect 140378 128194 140406 128452
rect 141298 128194 141326 128452
rect 142218 128194 142246 128452
rect 143138 128194 143166 128452
rect 144058 128194 144086 128452
rect 144978 128194 145006 128452
rect 145898 128194 145926 128452
rect 128464 128166 129550 128194
rect 129844 128166 130470 128194
rect 131224 128166 131390 128194
rect 132236 128166 132310 128194
rect 132604 128166 133230 128194
rect 133892 128166 134058 128194
rect 134168 128166 134978 128194
rect 135272 128166 135898 128194
rect 136744 128166 136818 128194
rect 137664 128166 137738 128194
rect 138032 128166 138658 128194
rect 139504 128166 139578 128194
rect 139688 128166 140406 128194
rect 140792 128166 141326 128194
rect 142172 128166 142246 128194
rect 142356 128166 143166 128194
rect 144012 128166 144086 128194
rect 144932 128166 145006 128194
rect 145852 128166 145926 128194
rect 146300 128240 146352 128246
rect 146726 128194 146754 128452
rect 147646 128246 147674 128452
rect 146300 128182 146352 128188
rect 128360 126268 128412 126274
rect 128360 126210 128412 126216
rect 126244 26920 126296 26926
rect 126244 26862 126296 26868
rect 126888 26920 126940 26926
rect 126888 26862 126940 26868
rect 125692 10328 125744 10334
rect 125692 10270 125744 10276
rect 125336 6886 125548 6914
rect 124218 3768 124274 3777
rect 124218 3703 124274 3712
rect 125336 3466 125364 6886
rect 126900 3466 126928 26862
rect 128464 7682 128492 128166
rect 129004 125656 129056 125662
rect 129004 125598 129056 125604
rect 129016 49026 129044 125598
rect 129004 49020 129056 49026
rect 129004 48962 129056 48968
rect 128452 7676 128504 7682
rect 128452 7618 128504 7624
rect 129372 7608 129424 7614
rect 129372 7550 129424 7556
rect 128176 4820 128228 4826
rect 128176 4762 128228 4768
rect 126980 4208 127032 4214
rect 126980 4150 127032 4156
rect 123484 3460 123536 3466
rect 123484 3402 123536 3408
rect 124128 3460 124180 3466
rect 124128 3402 124180 3408
rect 124680 3460 124732 3466
rect 124680 3402 124732 3408
rect 125324 3460 125376 3466
rect 125324 3402 125376 3408
rect 125876 3460 125928 3466
rect 125876 3402 125928 3408
rect 126888 3460 126940 3466
rect 126888 3402 126940 3408
rect 120264 3052 120316 3058
rect 120264 2994 120316 3000
rect 122288 3052 122340 3058
rect 122288 2994 122340 3000
rect 119896 2984 119948 2990
rect 119896 2926 119948 2932
rect 118976 2916 119028 2922
rect 118976 2858 119028 2864
rect 118792 2848 118844 2854
rect 118792 2790 118844 2796
rect 118804 480 118832 2790
rect 119908 480 119936 2926
rect 121092 2916 121144 2922
rect 121092 2858 121144 2864
rect 121104 480 121132 2858
rect 122300 480 122328 2994
rect 123496 480 123524 3402
rect 124692 480 124720 3402
rect 125888 480 125916 3402
rect 126060 3120 126112 3126
rect 126060 3062 126112 3068
rect 126072 2990 126100 3062
rect 126060 2984 126112 2990
rect 126060 2926 126112 2932
rect 126992 480 127020 4150
rect 127070 3632 127126 3641
rect 127070 3567 127126 3576
rect 127084 3466 127112 3567
rect 127072 3460 127124 3466
rect 127072 3402 127124 3408
rect 128188 480 128216 4762
rect 129384 480 129412 7550
rect 129844 3505 129872 128166
rect 130384 126336 130436 126342
rect 130384 126278 130436 126284
rect 130396 4214 130424 126278
rect 130568 8968 130620 8974
rect 130568 8910 130620 8916
rect 130384 4208 130436 4214
rect 130384 4150 130436 4156
rect 129830 3496 129886 3505
rect 129830 3431 129886 3440
rect 130580 480 130608 8910
rect 131224 3369 131252 128166
rect 132236 125662 132264 128166
rect 132224 125656 132276 125662
rect 132224 125598 132276 125604
rect 131764 5092 131816 5098
rect 131764 5034 131816 5040
rect 131210 3360 131266 3369
rect 131210 3295 131266 3304
rect 131776 480 131804 5034
rect 132604 3738 132632 128166
rect 133144 125656 133196 125662
rect 133144 125598 133196 125604
rect 133156 18630 133184 125598
rect 133144 18624 133196 18630
rect 133144 18566 133196 18572
rect 133788 15972 133840 15978
rect 133788 15914 133840 15920
rect 132592 3732 132644 3738
rect 132592 3674 132644 3680
rect 133800 3534 133828 15914
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 132972 480 133000 3470
rect 133892 3466 133920 128166
rect 134168 15910 134196 128166
rect 134156 15904 134208 15910
rect 134156 15846 134208 15852
rect 134156 5228 134208 5234
rect 134156 5170 134208 5176
rect 133880 3460 133932 3466
rect 133880 3402 133932 3408
rect 134168 480 134196 5170
rect 135272 3602 135300 128166
rect 136456 5296 136508 5302
rect 136456 5238 136508 5244
rect 135352 5160 135404 5166
rect 135352 5102 135404 5108
rect 135260 3596 135312 3602
rect 135260 3538 135312 3544
rect 135364 2666 135392 5102
rect 135272 2638 135392 2666
rect 135272 480 135300 2638
rect 136468 480 136496 5238
rect 136744 3738 136772 128166
rect 137664 125662 137692 128166
rect 137928 126268 137980 126274
rect 137928 126210 137980 126216
rect 137652 125656 137704 125662
rect 137652 125598 137704 125604
rect 137940 6914 137968 126210
rect 137664 6886 137968 6914
rect 136732 3732 136784 3738
rect 136732 3674 136784 3680
rect 137664 480 137692 6886
rect 138032 3874 138060 128166
rect 139504 126410 139532 128166
rect 139492 126404 139544 126410
rect 139492 126346 139544 126352
rect 139688 4962 139716 128166
rect 139676 4956 139728 4962
rect 139676 4898 139728 4904
rect 140044 4956 140096 4962
rect 140044 4898 140096 4904
rect 138020 3868 138072 3874
rect 138020 3810 138072 3816
rect 138848 3460 138900 3466
rect 138848 3402 138900 3408
rect 138860 480 138888 3402
rect 140056 480 140084 4898
rect 140792 3806 140820 128166
rect 142068 126404 142120 126410
rect 142068 126346 142120 126352
rect 140780 3800 140832 3806
rect 140780 3742 140832 3748
rect 142080 3534 142108 126346
rect 142172 3670 142200 128166
rect 142356 4894 142384 128166
rect 144012 126478 144040 128166
rect 144000 126472 144052 126478
rect 144000 126414 144052 126420
rect 144828 126472 144880 126478
rect 144828 126414 144880 126420
rect 144184 126200 144236 126206
rect 144184 126142 144236 126148
rect 144196 8974 144224 126142
rect 144184 8968 144236 8974
rect 144184 8910 144236 8916
rect 143540 8900 143592 8906
rect 143540 8842 143592 8848
rect 142344 4888 142396 4894
rect 142344 4830 142396 4836
rect 142160 3664 142212 3670
rect 142160 3606 142212 3612
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 142068 3528 142120 3534
rect 142068 3470 142120 3476
rect 141252 480 141280 3470
rect 142436 3324 142488 3330
rect 142436 3266 142488 3272
rect 142448 480 142476 3266
rect 143552 480 143580 8842
rect 144840 6914 144868 126414
rect 144748 6886 144868 6914
rect 144748 480 144776 6886
rect 144932 3942 144960 128166
rect 145852 126886 145880 128166
rect 145840 126880 145892 126886
rect 145840 126822 145892 126828
rect 146312 4078 146340 128182
rect 146404 128166 146754 128194
rect 147634 128240 147686 128246
rect 148566 128194 148594 128452
rect 147634 128182 147686 128188
rect 148520 128166 148594 128194
rect 149060 128240 149112 128246
rect 149486 128194 149514 128452
rect 150406 128246 150434 128452
rect 149060 128182 149112 128188
rect 146404 4146 146432 128166
rect 148520 126546 148548 128166
rect 148508 126540 148560 126546
rect 148508 126482 148560 126488
rect 148968 126540 149020 126546
rect 148968 126482 149020 126488
rect 148324 126132 148376 126138
rect 148324 126074 148376 126080
rect 148336 5302 148364 126074
rect 148324 5296 148376 5302
rect 148324 5238 148376 5244
rect 146392 4140 146444 4146
rect 146392 4082 146444 4088
rect 146300 4072 146352 4078
rect 146300 4014 146352 4020
rect 144920 3936 144972 3942
rect 144920 3878 144972 3884
rect 147128 3664 147180 3670
rect 147128 3606 147180 3612
rect 145932 3596 145984 3602
rect 145932 3538 145984 3544
rect 145944 480 145972 3538
rect 147140 480 147168 3606
rect 148980 3534 149008 126482
rect 149072 3738 149100 128182
rect 149164 128166 149514 128194
rect 150394 128240 150446 128246
rect 151326 128194 151354 128452
rect 152246 128194 152274 128452
rect 153074 128194 153102 128452
rect 153994 128194 154022 128452
rect 154914 128194 154942 128452
rect 155834 128194 155862 128452
rect 156754 128194 156782 128452
rect 150394 128182 150446 128188
rect 150544 128166 151354 128194
rect 152016 128166 152274 128194
rect 153028 128166 153102 128194
rect 153948 128166 154022 128194
rect 154592 128166 154942 128194
rect 155052 128166 155862 128194
rect 155972 128166 156782 128194
rect 157432 128240 157484 128246
rect 157674 128194 157702 128452
rect 158594 128246 158622 128452
rect 157432 128182 157484 128188
rect 149164 4010 149192 128166
rect 150544 5030 150572 128166
rect 151084 126064 151136 126070
rect 151084 126006 151136 126012
rect 151096 7614 151124 126006
rect 151084 7608 151136 7614
rect 151084 7550 151136 7556
rect 150532 5024 150584 5030
rect 150532 4966 150584 4972
rect 149152 4004 149204 4010
rect 149152 3946 149204 3952
rect 151820 3936 151872 3942
rect 151820 3878 151872 3884
rect 149520 3800 149572 3806
rect 149520 3742 149572 3748
rect 149060 3732 149112 3738
rect 149060 3674 149112 3680
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 148336 480 148364 3470
rect 149532 480 149560 3742
rect 150624 3732 150676 3738
rect 150624 3674 150676 3680
rect 150636 480 150664 3674
rect 151832 480 151860 3878
rect 152016 3262 152044 128166
rect 152556 126676 152608 126682
rect 152556 126618 152608 126624
rect 152568 124914 152596 126618
rect 153028 126614 153056 128166
rect 153948 126682 153976 128166
rect 153936 126676 153988 126682
rect 153936 126618 153988 126624
rect 153016 126608 153068 126614
rect 153016 126550 153068 126556
rect 153108 126608 153160 126614
rect 153108 126550 153160 126556
rect 152556 124908 152608 124914
rect 152556 124850 152608 124856
rect 153120 6914 153148 126550
rect 153028 6886 153148 6914
rect 152004 3256 152056 3262
rect 152004 3198 152056 3204
rect 153028 480 153056 6886
rect 154592 3398 154620 128166
rect 155052 122834 155080 128166
rect 154684 122806 155080 122834
rect 154580 3392 154632 3398
rect 154580 3334 154632 3340
rect 154684 3262 154712 122806
rect 155972 11762 156000 128166
rect 155960 11756 156012 11762
rect 155960 11698 156012 11704
rect 155408 4004 155460 4010
rect 155408 3946 155460 3952
rect 154672 3256 154724 3262
rect 154672 3198 154724 3204
rect 154212 3188 154264 3194
rect 154212 3130 154264 3136
rect 154224 480 154252 3130
rect 155420 480 155448 3946
rect 156604 3868 156656 3874
rect 156604 3810 156656 3816
rect 156616 480 156644 3810
rect 157444 2990 157472 128182
rect 157628 128166 157702 128194
rect 158582 128240 158634 128246
rect 159514 128194 159542 128452
rect 160342 128194 160370 128452
rect 161262 128194 161290 128452
rect 162182 128194 162210 128452
rect 163102 128194 163130 128452
rect 164022 128194 164050 128452
rect 164942 128194 164970 128452
rect 165862 128330 165890 128452
rect 158582 128182 158634 128188
rect 158824 128166 159542 128194
rect 160204 128166 160370 128194
rect 160480 128166 161290 128194
rect 161584 128166 162210 128194
rect 163056 128166 163130 128194
rect 163976 128166 164050 128194
rect 164252 128166 164970 128194
rect 165632 128302 165890 128330
rect 157628 126750 157656 128166
rect 157616 126744 157668 126750
rect 157616 126686 157668 126692
rect 158628 126676 158680 126682
rect 158628 126618 158680 126624
rect 158640 3398 158668 126618
rect 157800 3392 157852 3398
rect 157800 3334 157852 3340
rect 158628 3392 158680 3398
rect 158628 3334 158680 3340
rect 157432 2984 157484 2990
rect 157432 2926 157484 2932
rect 157812 480 157840 3334
rect 158824 2854 158852 128166
rect 160008 126880 160060 126886
rect 160008 126822 160060 126828
rect 160020 3398 160048 126822
rect 158904 3392 158956 3398
rect 158904 3334 158956 3340
rect 160008 3392 160060 3398
rect 160008 3334 160060 3340
rect 160100 3392 160152 3398
rect 160100 3334 160152 3340
rect 158812 2848 158864 2854
rect 158812 2790 158864 2796
rect 158916 480 158944 3334
rect 160112 480 160140 3334
rect 160204 3126 160232 128166
rect 160192 3120 160244 3126
rect 160192 3062 160244 3068
rect 160480 2922 160508 128166
rect 161296 4888 161348 4894
rect 161296 4830 161348 4836
rect 160468 2916 160520 2922
rect 160468 2858 160520 2864
rect 161308 480 161336 4830
rect 161584 3058 161612 128166
rect 163056 126818 163084 128166
rect 163976 126954 164004 128166
rect 163964 126948 164016 126954
rect 163964 126890 164016 126896
rect 163044 126812 163096 126818
rect 163044 126754 163096 126760
rect 162768 126744 162820 126750
rect 162768 126686 162820 126692
rect 162780 6914 162808 126686
rect 164252 26926 164280 128166
rect 165632 126342 165660 128302
rect 166690 128194 166718 128452
rect 167610 128194 167638 128452
rect 168530 128194 168558 128452
rect 169450 128194 169478 128452
rect 170370 128194 170398 128452
rect 171290 128194 171318 128452
rect 172210 128194 172238 128452
rect 173038 128194 173066 128452
rect 173958 128194 173986 128452
rect 174878 128194 174906 128452
rect 175798 128194 175826 128452
rect 176718 128194 176746 128452
rect 177638 128194 177666 128452
rect 178558 128194 178586 128452
rect 179386 128194 179414 128452
rect 180306 128194 180334 128452
rect 181226 128194 181254 128452
rect 182146 128194 182174 128452
rect 183066 128194 183094 128452
rect 183986 128194 184014 128452
rect 184906 128194 184934 128452
rect 185734 128194 185762 128452
rect 165724 128166 166718 128194
rect 167564 128166 167638 128194
rect 168484 128166 168558 128194
rect 168668 128166 169478 128194
rect 169772 128166 170398 128194
rect 171244 128166 171318 128194
rect 172164 128166 172238 128194
rect 172992 128166 173066 128194
rect 173912 128166 173986 128194
rect 174096 128166 174906 128194
rect 175292 128166 175826 128194
rect 176672 128166 176746 128194
rect 176856 128166 177666 128194
rect 178144 128166 178586 128194
rect 179340 128166 179414 128194
rect 179524 128166 180334 128194
rect 180996 128166 181254 128194
rect 182100 128166 182174 128194
rect 182284 128166 183094 128194
rect 183572 128166 184014 128194
rect 184860 128166 184934 128194
rect 185688 128166 185762 128194
rect 186412 128240 186464 128246
rect 186654 128194 186682 128452
rect 187574 128246 187602 128452
rect 186412 128182 186464 128188
rect 165620 126336 165672 126342
rect 165620 126278 165672 126284
rect 164884 126132 164936 126138
rect 164884 126074 164936 126080
rect 164240 26920 164292 26926
rect 164240 26862 164292 26868
rect 162504 6886 162808 6914
rect 161572 3052 161624 3058
rect 161572 2994 161624 3000
rect 162504 480 162532 6886
rect 164896 5234 164924 126074
rect 164884 5228 164936 5234
rect 164884 5170 164936 5176
rect 165724 4826 165752 128166
rect 166908 126336 166960 126342
rect 166908 126278 166960 126284
rect 165712 4820 165764 4826
rect 165712 4762 165764 4768
rect 163688 4140 163740 4146
rect 163688 4082 163740 4088
rect 163700 480 163728 4082
rect 164884 4072 164936 4078
rect 164884 4014 164936 4020
rect 164896 480 164924 4014
rect 166920 3330 166948 126278
rect 167564 125934 167592 128166
rect 168484 126206 168512 128166
rect 168472 126200 168524 126206
rect 168472 126142 168524 126148
rect 167552 125928 167604 125934
rect 167552 125870 167604 125876
rect 168668 5098 168696 128166
rect 169668 126200 169720 126206
rect 169668 126142 169720 126148
rect 169680 6914 169708 126142
rect 169772 15978 169800 128166
rect 170404 126948 170456 126954
rect 170404 126890 170456 126896
rect 169760 15972 169812 15978
rect 169760 15914 169812 15920
rect 169588 6886 169708 6914
rect 168656 5092 168708 5098
rect 168656 5034 168708 5040
rect 166080 3324 166132 3330
rect 166080 3266 166132 3272
rect 166908 3324 166960 3330
rect 166908 3266 166960 3272
rect 166092 480 166120 3266
rect 168380 3256 168432 3262
rect 168380 3198 168432 3204
rect 167184 3120 167236 3126
rect 167184 3062 167236 3068
rect 167196 480 167224 3062
rect 168392 480 168420 3198
rect 169588 480 169616 6886
rect 170416 5166 170444 126890
rect 171048 126812 171100 126818
rect 171048 126754 171100 126760
rect 171060 6914 171088 126754
rect 171244 126138 171272 128166
rect 172164 126954 172192 128166
rect 172152 126948 172204 126954
rect 172152 126890 172204 126896
rect 171232 126132 171284 126138
rect 171232 126074 171284 126080
rect 172992 126002 173020 128166
rect 173912 126274 173940 128166
rect 173900 126268 173952 126274
rect 173900 126210 173952 126216
rect 173808 126200 173860 126206
rect 173808 126142 173860 126148
rect 173164 126132 173216 126138
rect 173164 126074 173216 126080
rect 172980 125996 173032 126002
rect 172980 125938 173032 125944
rect 173176 6914 173204 126074
rect 170784 6886 171088 6914
rect 173084 6886 173204 6914
rect 170404 5160 170456 5166
rect 170404 5102 170456 5108
rect 170784 480 170812 6886
rect 171968 3324 172020 3330
rect 171968 3266 172020 3272
rect 171980 480 172008 3266
rect 173084 3194 173112 6886
rect 173820 3534 173848 126142
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 173072 3188 173124 3194
rect 173072 3130 173124 3136
rect 173176 480 173204 3470
rect 174096 3466 174124 128166
rect 175292 4962 175320 128166
rect 176672 126410 176700 128166
rect 176660 126404 176712 126410
rect 176660 126346 176712 126352
rect 175280 4956 175332 4962
rect 175280 4898 175332 4904
rect 176856 3806 176884 128166
rect 177948 126404 178000 126410
rect 177948 126346 178000 126352
rect 176844 3800 176896 3806
rect 176844 3742 176896 3748
rect 174268 3664 174320 3670
rect 174268 3606 174320 3612
rect 174084 3460 174136 3466
rect 174084 3402 174136 3408
rect 174280 480 174308 3606
rect 177960 3534 177988 126346
rect 178144 8974 178172 128166
rect 179340 126478 179368 128166
rect 179328 126472 179380 126478
rect 179328 126414 179380 126420
rect 178684 125860 178736 125866
rect 178684 125802 178736 125808
rect 178132 8968 178184 8974
rect 178132 8910 178184 8916
rect 178696 4894 178724 125802
rect 178684 4888 178736 4894
rect 178684 4830 178736 4836
rect 179524 3534 179552 128166
rect 180708 126268 180760 126274
rect 180708 126210 180760 126216
rect 180064 126064 180116 126070
rect 180064 126006 180116 126012
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 177948 3528 178000 3534
rect 177948 3470 178000 3476
rect 179512 3528 179564 3534
rect 179512 3470 179564 3476
rect 175464 3188 175516 3194
rect 175464 3130 175516 3136
rect 175476 480 175504 3130
rect 176672 480 176700 3470
rect 179052 3460 179104 3466
rect 179052 3402 179104 3408
rect 177856 3052 177908 3058
rect 177856 2994 177908 3000
rect 177868 480 177896 2994
rect 179064 480 179092 3402
rect 180076 3126 180104 126006
rect 180720 3806 180748 126210
rect 180248 3800 180300 3806
rect 180248 3742 180300 3748
rect 180708 3800 180760 3806
rect 180708 3742 180760 3748
rect 180064 3120 180116 3126
rect 180064 3062 180116 3068
rect 180260 480 180288 3742
rect 180996 3602 181024 128166
rect 182100 126546 182128 128166
rect 182088 126540 182140 126546
rect 182088 126482 182140 126488
rect 181444 125996 181496 126002
rect 181444 125938 181496 125944
rect 181456 3670 181484 125938
rect 181444 3664 181496 3670
rect 181444 3606 181496 3612
rect 180984 3596 181036 3602
rect 180984 3538 181036 3544
rect 181444 3120 181496 3126
rect 181444 3062 181496 3068
rect 181456 480 181484 3062
rect 182284 2990 182312 128166
rect 183572 3738 183600 128166
rect 184756 126472 184808 126478
rect 184756 126414 184808 126420
rect 184204 125928 184256 125934
rect 184204 125870 184256 125876
rect 183652 125656 183704 125662
rect 183652 125598 183704 125604
rect 183664 3942 183692 125598
rect 183652 3936 183704 3942
rect 183652 3878 183704 3884
rect 183560 3732 183612 3738
rect 183560 3674 183612 3680
rect 182548 3664 182600 3670
rect 182548 3606 182600 3612
rect 182272 2984 182324 2990
rect 182272 2926 182324 2932
rect 182560 480 182588 3606
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 183756 480 183784 3470
rect 184216 3058 184244 125870
rect 184768 122834 184796 126414
rect 184860 125662 184888 128166
rect 185688 126614 185716 128166
rect 185676 126608 185728 126614
rect 185676 126550 185728 126556
rect 184848 125656 184900 125662
rect 184848 125598 184900 125604
rect 184768 122806 184888 122834
rect 184860 3534 184888 122806
rect 186424 4010 186452 128182
rect 186608 128166 186682 128194
rect 187562 128240 187614 128246
rect 188494 128194 188522 128452
rect 189414 128194 189442 128452
rect 190334 128194 190362 128452
rect 191254 128194 191282 128452
rect 192082 128194 192110 128452
rect 193002 128194 193030 128452
rect 193922 128194 193950 128452
rect 194842 128194 194870 128452
rect 195762 128194 195790 128452
rect 196682 128194 196710 128452
rect 197602 128194 197630 128452
rect 198430 128194 198458 128452
rect 199350 128194 199378 128452
rect 187562 128182 187614 128188
rect 187712 128166 188522 128194
rect 189368 128166 189442 128194
rect 190288 128166 190362 128194
rect 190564 128166 191282 128194
rect 192036 128166 192110 128194
rect 192956 128166 193030 128194
rect 193232 128166 193950 128194
rect 194704 128166 194870 128194
rect 195716 128166 195790 128194
rect 196636 128166 196710 128194
rect 197464 128166 197630 128194
rect 198384 128166 198458 128194
rect 199304 128166 199378 128194
rect 200270 128194 200298 128452
rect 201190 128194 201218 128452
rect 202110 128194 202138 128452
rect 203030 128194 203058 128452
rect 203950 128194 203978 128452
rect 204870 128194 204898 128452
rect 200270 128166 200344 128194
rect 186608 126138 186636 128166
rect 187608 126540 187660 126546
rect 187608 126482 187660 126488
rect 186596 126132 186648 126138
rect 186596 126074 186648 126080
rect 186964 126132 187016 126138
rect 186964 126074 187016 126080
rect 186412 4004 186464 4010
rect 186412 3946 186464 3952
rect 186136 3596 186188 3602
rect 186136 3538 186188 3544
rect 184848 3528 184900 3534
rect 184848 3470 184900 3476
rect 184940 3528 184992 3534
rect 184940 3470 184992 3476
rect 184204 3052 184256 3058
rect 184204 2994 184256 3000
rect 184952 480 184980 3470
rect 186148 480 186176 3538
rect 186976 3534 187004 126074
rect 187620 6914 187648 126482
rect 187344 6886 187648 6914
rect 186964 3528 187016 3534
rect 186964 3470 187016 3476
rect 187344 480 187372 6886
rect 187712 3874 187740 128166
rect 189368 126682 189396 128166
rect 190288 126886 190316 128166
rect 190276 126880 190328 126886
rect 190276 126822 190328 126828
rect 189356 126676 189408 126682
rect 189356 126618 189408 126624
rect 188988 126608 189040 126614
rect 188988 126550 189040 126556
rect 187700 3868 187752 3874
rect 187700 3810 187752 3816
rect 189000 3670 189028 126550
rect 189724 3732 189776 3738
rect 189724 3674 189776 3680
rect 188528 3664 188580 3670
rect 188528 3606 188580 3612
rect 188988 3664 189040 3670
rect 188988 3606 189040 3612
rect 188540 480 188568 3606
rect 189736 480 189764 3674
rect 190564 3398 190592 128166
rect 191748 126676 191800 126682
rect 191748 126618 191800 126624
rect 191760 3398 191788 126618
rect 192036 125866 192064 128166
rect 192956 126750 192984 128166
rect 192944 126744 192996 126750
rect 192944 126686 192996 126692
rect 193128 126744 193180 126750
rect 193128 126686 193180 126692
rect 192024 125860 192076 125866
rect 192024 125802 192076 125808
rect 193140 3398 193168 126686
rect 193232 4146 193260 128166
rect 193220 4140 193272 4146
rect 193220 4082 193272 4088
rect 194704 4078 194732 128166
rect 195244 126880 195296 126886
rect 195244 126822 195296 126828
rect 194692 4072 194744 4078
rect 194692 4014 194744 4020
rect 193220 3868 193272 3874
rect 193220 3810 193272 3816
rect 190552 3392 190604 3398
rect 190552 3334 190604 3340
rect 190828 3392 190880 3398
rect 190828 3334 190880 3340
rect 191748 3392 191800 3398
rect 191748 3334 191800 3340
rect 192024 3392 192076 3398
rect 192024 3334 192076 3340
rect 193128 3392 193180 3398
rect 193128 3334 193180 3340
rect 190840 480 190868 3334
rect 192036 480 192064 3334
rect 193232 480 193260 3810
rect 195256 3398 195284 126822
rect 195716 126342 195744 128166
rect 195704 126336 195756 126342
rect 195704 126278 195756 126284
rect 195888 126336 195940 126342
rect 195888 126278 195940 126284
rect 195900 6914 195928 126278
rect 196636 126070 196664 128166
rect 196624 126064 196676 126070
rect 196624 126006 196676 126012
rect 195624 6886 195928 6914
rect 194416 3392 194468 3398
rect 194416 3334 194468 3340
rect 195244 3392 195296 3398
rect 195244 3334 195296 3340
rect 194428 480 194456 3334
rect 195624 480 195652 6886
rect 196808 3800 196860 3806
rect 196808 3742 196860 3748
rect 196820 480 196848 3742
rect 197464 3262 197492 128166
rect 198384 126818 198412 128166
rect 199304 126954 199332 128166
rect 199292 126948 199344 126954
rect 199292 126890 199344 126896
rect 200028 126948 200080 126954
rect 200028 126890 200080 126896
rect 198372 126812 198424 126818
rect 198372 126754 198424 126760
rect 198648 126064 198700 126070
rect 198648 126006 198700 126012
rect 198660 3398 198688 126006
rect 200040 3398 200068 126890
rect 200316 6914 200344 128166
rect 201144 128166 201218 128194
rect 202064 128166 202138 128194
rect 202984 128166 203058 128194
rect 203904 128166 203978 128194
rect 204824 128166 204898 128194
rect 205698 128194 205726 128452
rect 206618 128194 206646 128452
rect 207538 128194 207566 128452
rect 205698 128166 205772 128194
rect 201144 126206 201172 128166
rect 201132 126200 201184 126206
rect 201132 126142 201184 126148
rect 202064 126002 202092 128166
rect 202696 126812 202748 126818
rect 202696 126754 202748 126760
rect 202052 125996 202104 126002
rect 202052 125938 202104 125944
rect 200224 6886 200344 6914
rect 197912 3392 197964 3398
rect 197912 3334 197964 3340
rect 198648 3392 198700 3398
rect 198648 3334 198700 3340
rect 199108 3392 199160 3398
rect 199108 3334 199160 3340
rect 200028 3392 200080 3398
rect 200028 3334 200080 3340
rect 197452 3256 197504 3262
rect 197452 3198 197504 3204
rect 197924 480 197952 3334
rect 199120 480 199148 3334
rect 200224 3330 200252 6886
rect 200304 3936 200356 3942
rect 200304 3878 200356 3884
rect 200212 3324 200264 3330
rect 200212 3266 200264 3272
rect 200316 480 200344 3878
rect 201500 3528 201552 3534
rect 201500 3470 201552 3476
rect 201512 480 201540 3470
rect 202708 480 202736 126754
rect 202788 126200 202840 126206
rect 202788 126142 202840 126148
rect 202800 3534 202828 126142
rect 202788 3528 202840 3534
rect 202788 3470 202840 3476
rect 202984 3194 203012 128166
rect 203904 126410 203932 128166
rect 203892 126404 203944 126410
rect 203892 126346 203944 126352
rect 204168 125996 204220 126002
rect 204168 125938 204220 125944
rect 204180 6914 204208 125938
rect 204824 125934 204852 128166
rect 204812 125928 204864 125934
rect 204812 125870 204864 125876
rect 205548 125860 205600 125866
rect 205548 125802 205600 125808
rect 203904 6886 204208 6914
rect 202972 3188 203024 3194
rect 202972 3130 203024 3136
rect 203904 480 203932 6886
rect 205560 3534 205588 125802
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 205100 480 205128 3470
rect 205744 3466 205772 128166
rect 206572 128166 206646 128194
rect 207492 128166 207566 128194
rect 208458 128194 208486 128452
rect 209378 128194 209406 128452
rect 210298 128194 210326 128452
rect 211218 128194 211246 128452
rect 212046 128194 212074 128452
rect 208458 128166 208532 128194
rect 206572 126274 206600 128166
rect 206560 126268 206612 126274
rect 206560 126210 206612 126216
rect 206928 126268 206980 126274
rect 206928 126210 206980 126216
rect 206284 125656 206336 125662
rect 206284 125598 206336 125604
rect 206192 3528 206244 3534
rect 206192 3470 206244 3476
rect 205732 3460 205784 3466
rect 205732 3402 205784 3408
rect 206204 480 206232 3470
rect 206296 3126 206324 125598
rect 206940 3534 206968 126210
rect 207492 125662 207520 128166
rect 208308 125928 208360 125934
rect 208308 125870 208360 125876
rect 207480 125656 207532 125662
rect 207480 125598 207532 125604
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 208320 3194 208348 125870
rect 208504 3670 208532 128166
rect 209332 128166 209406 128194
rect 210252 128166 210326 128194
rect 211172 128166 211246 128194
rect 212000 128166 212074 128194
rect 212632 128240 212684 128246
rect 212966 128194 212994 128452
rect 213886 128246 213914 128452
rect 212632 128182 212684 128188
rect 209332 126478 209360 128166
rect 209320 126472 209372 126478
rect 209320 126414 209372 126420
rect 209688 126472 209740 126478
rect 209688 126414 209740 126420
rect 208492 3664 208544 3670
rect 208492 3606 208544 3612
rect 209700 3534 209728 126414
rect 210252 126138 210280 128166
rect 210240 126132 210292 126138
rect 210240 126074 210292 126080
rect 211068 126132 211120 126138
rect 211068 126074 211120 126080
rect 211080 6914 211108 126074
rect 210988 6886 211108 6914
rect 208584 3528 208636 3534
rect 208584 3470 208636 3476
rect 209688 3528 209740 3534
rect 209688 3470 209740 3476
rect 207388 3188 207440 3194
rect 207388 3130 207440 3136
rect 208308 3188 208360 3194
rect 208308 3130 208360 3136
rect 206284 3120 206336 3126
rect 206284 3062 206336 3068
rect 207400 480 207428 3130
rect 208596 480 208624 3470
rect 209780 3324 209832 3330
rect 209780 3266 209832 3272
rect 209792 480 209820 3266
rect 210988 480 211016 6886
rect 211172 3602 211200 128166
rect 212000 126410 212028 128166
rect 212448 126540 212500 126546
rect 212448 126482 212500 126488
rect 211988 126404 212040 126410
rect 211988 126346 212040 126352
rect 212460 6914 212488 126482
rect 212184 6886 212488 6914
rect 211160 3596 211212 3602
rect 211160 3538 211212 3544
rect 212184 480 212212 6886
rect 212644 3738 212672 128182
rect 212920 128166 212994 128194
rect 213874 128240 213926 128246
rect 214806 128194 214834 128452
rect 213874 128182 213926 128188
rect 214760 128166 214834 128194
rect 215392 128240 215444 128246
rect 215726 128194 215754 128452
rect 216646 128246 216674 128452
rect 215392 128182 215444 128188
rect 212920 126614 212948 128166
rect 214760 126682 214788 128166
rect 214748 126676 214800 126682
rect 214748 126618 214800 126624
rect 212908 126608 212960 126614
rect 212908 126550 212960 126556
rect 213828 126608 213880 126614
rect 213828 126550 213880 126556
rect 213184 125792 213236 125798
rect 213184 125734 213236 125740
rect 212632 3732 212684 3738
rect 212632 3674 212684 3680
rect 213196 3330 213224 125734
rect 213840 3534 213868 126550
rect 215208 125860 215260 125866
rect 215208 125802 215260 125808
rect 215220 3534 215248 125802
rect 215404 3874 215432 128182
rect 215680 128166 215754 128194
rect 216634 128240 216686 128246
rect 217566 128194 217594 128452
rect 216634 128182 216686 128188
rect 217520 128166 217594 128194
rect 218152 128240 218204 128246
rect 218394 128194 218422 128452
rect 219314 128246 219342 128452
rect 218152 128182 218204 128188
rect 215680 126750 215708 128166
rect 217520 126886 217548 128166
rect 217508 126880 217560 126886
rect 217508 126822 217560 126828
rect 215668 126744 215720 126750
rect 215668 126686 215720 126692
rect 216588 126744 216640 126750
rect 216588 126686 216640 126692
rect 215392 3868 215444 3874
rect 215392 3810 215444 3816
rect 216600 3534 216628 126686
rect 217968 126676 218020 126682
rect 217968 126618 218020 126624
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213828 3528 213880 3534
rect 213828 3470 213880 3476
rect 214472 3528 214524 3534
rect 214472 3470 214524 3476
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 213184 3324 213236 3330
rect 213184 3266 213236 3272
rect 213380 480 213408 3470
rect 214484 480 214512 3470
rect 215680 480 215708 3470
rect 217980 3262 218008 126618
rect 218164 3806 218192 128182
rect 218348 128166 218422 128194
rect 219302 128240 219354 128246
rect 220234 128194 220262 128452
rect 219302 128182 219354 128188
rect 220188 128166 220262 128194
rect 220912 128240 220964 128246
rect 221154 128194 221182 128452
rect 222074 128246 222102 128452
rect 220912 128182 220964 128188
rect 218348 126342 218376 128166
rect 220084 126880 220136 126886
rect 220084 126822 220136 126828
rect 218336 126336 218388 126342
rect 218336 126278 218388 126284
rect 219348 125724 219400 125730
rect 219348 125666 219400 125672
rect 219256 4140 219308 4146
rect 219256 4082 219308 4088
rect 218152 3800 218204 3806
rect 218152 3742 218204 3748
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 216864 3256 216916 3262
rect 216864 3198 216916 3204
rect 217968 3256 218020 3262
rect 217968 3198 218020 3204
rect 216876 480 216904 3198
rect 218072 480 218100 3470
rect 219268 480 219296 4082
rect 219360 3534 219388 125666
rect 220096 4146 220124 126822
rect 220188 126070 220216 128166
rect 220728 126336 220780 126342
rect 220728 126278 220780 126284
rect 220176 126064 220228 126070
rect 220176 126006 220228 126012
rect 220740 6914 220768 126278
rect 220464 6886 220768 6914
rect 220084 4140 220136 4146
rect 220084 4082 220136 4088
rect 219348 3528 219400 3534
rect 219348 3470 219400 3476
rect 220464 480 220492 6886
rect 220924 3942 220952 128182
rect 221108 128166 221182 128194
rect 222062 128240 222114 128246
rect 222994 128194 223022 128452
rect 223914 128194 223942 128452
rect 224742 128194 224770 128452
rect 225662 128194 225690 128452
rect 226582 128194 226610 128452
rect 227502 128194 227530 128452
rect 228422 128194 228450 128452
rect 229342 128194 229370 128452
rect 230262 128194 230290 128452
rect 231090 128194 231118 128452
rect 232010 128194 232038 128452
rect 232930 128194 232958 128452
rect 233850 128194 233878 128452
rect 234770 128194 234798 128452
rect 235690 128194 235718 128452
rect 236610 128194 236638 128452
rect 237438 128194 237466 128452
rect 238358 128194 238386 128452
rect 239278 128194 239306 128452
rect 240198 128194 240226 128452
rect 241118 128194 241146 128452
rect 242038 128194 242066 128452
rect 242958 128194 242986 128452
rect 243786 128194 243814 128452
rect 244706 128194 244734 128452
rect 245626 128194 245654 128452
rect 246546 128194 246574 128452
rect 247466 128194 247494 128452
rect 248386 128194 248414 128452
rect 249306 128194 249334 128452
rect 250226 128194 250254 128452
rect 251054 128194 251082 128452
rect 251974 128194 252002 128452
rect 252894 128194 252922 128452
rect 253814 128194 253842 128452
rect 254734 128194 254762 128452
rect 255654 128194 255682 128452
rect 256574 128194 256602 128452
rect 257402 128194 257430 128452
rect 258322 128194 258350 128452
rect 259242 128194 259270 128452
rect 260162 128194 260190 128452
rect 261082 128194 261110 128452
rect 262002 128194 262030 128452
rect 262922 128194 262950 128452
rect 263750 128194 263778 128452
rect 264670 128194 264698 128452
rect 265590 128194 265618 128452
rect 266510 128194 266538 128452
rect 267430 128194 267458 128452
rect 268350 128194 268378 128452
rect 269270 128194 269298 128452
rect 270098 128194 270126 128452
rect 271018 128194 271046 128452
rect 271938 128194 271966 128452
rect 272858 128194 272886 128452
rect 273778 128194 273806 128452
rect 274698 128194 274726 128452
rect 275618 128194 275646 128452
rect 276446 128194 276474 128452
rect 277366 128194 277394 128452
rect 278286 128194 278314 128452
rect 279206 128194 279234 128452
rect 280126 128194 280154 128452
rect 281046 128194 281074 128452
rect 281966 128194 281994 128452
rect 282794 128194 282822 128452
rect 283714 128194 283742 128452
rect 284634 128330 284662 128452
rect 222062 128182 222114 128188
rect 222948 128166 223022 128194
rect 223868 128166 223942 128194
rect 224696 128166 224770 128194
rect 225616 128166 225690 128194
rect 226536 128166 226610 128194
rect 227456 128166 227530 128194
rect 228376 128166 228450 128194
rect 229296 128166 229370 128194
rect 230216 128166 230290 128194
rect 231044 128166 231118 128194
rect 231964 128166 232038 128194
rect 232884 128166 232958 128194
rect 233804 128166 233878 128194
rect 234724 128166 234798 128194
rect 235644 128166 235718 128194
rect 236564 128166 236638 128194
rect 237392 128166 237466 128194
rect 238312 128166 238386 128194
rect 239232 128166 239306 128194
rect 240152 128166 240226 128194
rect 241072 128166 241146 128194
rect 241992 128166 242066 128194
rect 242912 128166 242986 128194
rect 243740 128166 243814 128194
rect 244660 128166 244734 128194
rect 245488 128166 245654 128194
rect 246500 128166 246574 128194
rect 247420 128166 247494 128194
rect 248340 128166 248414 128194
rect 249260 128166 249334 128194
rect 250180 128166 250254 128194
rect 251008 128166 251082 128194
rect 251928 128166 252002 128194
rect 252848 128166 252922 128194
rect 253768 128166 253842 128194
rect 254688 128166 254762 128194
rect 255608 128166 255682 128194
rect 256528 128166 256602 128194
rect 257356 128166 257430 128194
rect 258276 128166 258350 128194
rect 259196 128166 259270 128194
rect 260116 128166 260190 128194
rect 261036 128166 261110 128194
rect 261956 128166 262030 128194
rect 262876 128166 262950 128194
rect 263704 128166 263778 128194
rect 264624 128166 264698 128194
rect 265544 128166 265618 128194
rect 266464 128166 266538 128194
rect 267384 128166 267458 128194
rect 268304 128166 268378 128194
rect 269224 128166 269298 128194
rect 269408 128166 270126 128194
rect 270972 128166 271046 128194
rect 271892 128166 271966 128194
rect 272812 128166 272886 128194
rect 273732 128166 273806 128194
rect 274652 128166 274726 128194
rect 275572 128166 275646 128194
rect 276400 128166 276474 128194
rect 277320 128166 277394 128194
rect 277504 128166 278314 128194
rect 279160 128166 279234 128194
rect 280080 128166 280154 128194
rect 280356 128166 281074 128194
rect 281920 128166 281994 128194
rect 282748 128166 282822 128194
rect 283668 128166 283742 128194
rect 284404 128302 284662 128330
rect 221108 126954 221136 128166
rect 221096 126948 221148 126954
rect 221096 126890 221148 126896
rect 222948 126206 222976 128166
rect 223488 126948 223540 126954
rect 223488 126890 223540 126896
rect 222936 126200 222988 126206
rect 222936 126142 222988 126148
rect 222108 126064 222160 126070
rect 222108 126006 222160 126012
rect 220912 3936 220964 3942
rect 220912 3878 220964 3884
rect 222120 3126 222148 126006
rect 223500 3534 223528 126890
rect 223868 126818 223896 128166
rect 223856 126812 223908 126818
rect 223856 126754 223908 126760
rect 224696 126002 224724 128166
rect 224868 126812 224920 126818
rect 224868 126754 224920 126760
rect 224684 125996 224736 126002
rect 224684 125938 224736 125944
rect 224880 3534 224908 126754
rect 225616 126410 225644 128166
rect 225604 126404 225656 126410
rect 225604 126346 225656 126352
rect 226536 126274 226564 128166
rect 226524 126268 226576 126274
rect 226524 126210 226576 126216
rect 226984 126200 227036 126206
rect 226984 126142 227036 126148
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 221556 3120 221608 3126
rect 221556 3062 221608 3068
rect 222108 3120 222160 3126
rect 222108 3062 222160 3068
rect 221568 480 221596 3062
rect 222764 480 222792 3470
rect 223960 480 223988 3470
rect 225144 3052 225196 3058
rect 225144 2994 225196 3000
rect 225156 480 225184 2994
rect 226352 480 226380 3470
rect 226996 3058 227024 126142
rect 227456 125934 227484 128166
rect 228376 126478 228404 128166
rect 228364 126472 228416 126478
rect 228364 126414 228416 126420
rect 229008 126404 229060 126410
rect 229008 126346 229060 126352
rect 227628 126268 227680 126274
rect 227628 126210 227680 126216
rect 227444 125928 227496 125934
rect 227444 125870 227496 125876
rect 227640 3534 227668 126210
rect 229020 6914 229048 126346
rect 229296 125798 229324 128166
rect 230216 126138 230244 128166
rect 231044 126546 231072 128166
rect 231964 126614 231992 128166
rect 231952 126608 232004 126614
rect 231952 126550 232004 126556
rect 231032 126540 231084 126546
rect 231032 126482 231084 126488
rect 231124 126472 231176 126478
rect 231124 126414 231176 126420
rect 230204 126132 230256 126138
rect 230204 126074 230256 126080
rect 229284 125792 229336 125798
rect 229284 125734 229336 125740
rect 228744 6886 229048 6914
rect 227628 3528 227680 3534
rect 227628 3470 227680 3476
rect 227536 3392 227588 3398
rect 227536 3334 227588 3340
rect 226984 3052 227036 3058
rect 226984 2994 227036 3000
rect 227548 480 227576 3334
rect 228744 480 228772 6886
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 229836 3460 229888 3466
rect 229836 3402 229888 3408
rect 229848 480 229876 3402
rect 231044 480 231072 3470
rect 231136 3466 231164 126414
rect 231768 126132 231820 126138
rect 231768 126074 231820 126080
rect 231780 3534 231808 126074
rect 232884 125866 232912 128166
rect 233804 126750 233832 128166
rect 233792 126744 233844 126750
rect 233792 126686 233844 126692
rect 234724 126682 234752 128166
rect 234712 126676 234764 126682
rect 234712 126618 234764 126624
rect 234528 126540 234580 126546
rect 234528 126482 234580 126488
rect 233148 125996 233200 126002
rect 233148 125938 233200 125944
rect 232872 125860 232924 125866
rect 232872 125802 232924 125808
rect 233160 3534 233188 125938
rect 234540 3534 234568 126482
rect 235644 125730 235672 128166
rect 236564 126886 236592 128166
rect 236552 126880 236604 126886
rect 236552 126822 236604 126828
rect 235908 126676 235960 126682
rect 235908 126618 235960 126624
rect 235632 125724 235684 125730
rect 235632 125666 235684 125672
rect 235920 6914 235948 126618
rect 237288 126608 237340 126614
rect 237288 126550 237340 126556
rect 237300 6914 237328 126550
rect 237392 126342 237420 128166
rect 238024 126880 238076 126886
rect 238024 126822 238076 126828
rect 237380 126336 237432 126342
rect 237380 126278 237432 126284
rect 235828 6886 235948 6914
rect 237024 6886 237328 6914
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 231124 3460 231176 3466
rect 231124 3402 231176 3408
rect 232240 480 232268 3470
rect 233436 480 233464 3470
rect 234632 480 234660 3470
rect 235828 480 235856 6886
rect 237024 480 237052 6886
rect 238036 3398 238064 126822
rect 238312 126070 238340 128166
rect 239232 126954 239260 128166
rect 239220 126948 239272 126954
rect 239220 126890 239272 126896
rect 240152 126818 240180 128166
rect 240140 126812 240192 126818
rect 240140 126754 240192 126760
rect 238668 126744 238720 126750
rect 238668 126686 238720 126692
rect 238300 126064 238352 126070
rect 238300 126006 238352 126012
rect 238680 3466 238708 126686
rect 241072 126206 241100 128166
rect 241428 126336 241480 126342
rect 241428 126278 241480 126284
rect 241060 126200 241112 126206
rect 241060 126142 241112 126148
rect 238116 3460 238168 3466
rect 238116 3402 238168 3408
rect 238668 3460 238720 3466
rect 238668 3402 238720 3408
rect 238024 3392 238076 3398
rect 238024 3334 238076 3340
rect 238128 480 238156 3402
rect 239312 3188 239364 3194
rect 239312 3130 239364 3136
rect 239324 480 239352 3130
rect 241440 3058 241468 126278
rect 241992 126274 242020 128166
rect 242912 126886 242940 128166
rect 242900 126880 242952 126886
rect 242900 126822 242952 126828
rect 242808 126812 242860 126818
rect 242808 126754 242860 126760
rect 241980 126268 242032 126274
rect 241980 126210 242032 126216
rect 242164 125656 242216 125662
rect 242164 125598 242216 125604
rect 242176 3602 242204 125598
rect 242164 3596 242216 3602
rect 242164 3538 242216 3544
rect 242820 3534 242848 126754
rect 243740 126410 243768 128166
rect 244660 126478 244688 128166
rect 244648 126472 244700 126478
rect 244648 126414 244700 126420
rect 243728 126404 243780 126410
rect 243728 126346 243780 126352
rect 244924 126268 244976 126274
rect 244924 126210 244976 126216
rect 242900 4072 242952 4078
rect 242900 4014 242952 4020
rect 241704 3528 241756 3534
rect 241704 3470 241756 3476
rect 242808 3528 242860 3534
rect 242808 3470 242860 3476
rect 240508 3052 240560 3058
rect 240508 2994 240560 3000
rect 241428 3052 241480 3058
rect 241428 2994 241480 3000
rect 240520 480 240548 2994
rect 241716 480 241744 3470
rect 242912 480 242940 4014
rect 244936 3534 244964 126210
rect 245488 126138 245516 128166
rect 246304 126880 246356 126886
rect 246304 126822 246356 126828
rect 245568 126404 245620 126410
rect 245568 126346 245620 126352
rect 245476 126132 245528 126138
rect 245476 126074 245528 126080
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 244924 3528 244976 3534
rect 244924 3470 244976 3476
rect 244108 480 244136 3470
rect 245212 598 245424 626
rect 245212 480 245240 598
rect 245396 490 245424 598
rect 245580 490 245608 126346
rect 246316 3194 246344 126822
rect 246500 126002 246528 128166
rect 247420 126546 247448 128166
rect 247408 126540 247460 126546
rect 247408 126482 247460 126488
rect 246948 126472 247000 126478
rect 246948 126414 247000 126420
rect 246488 125996 246540 126002
rect 246488 125938 246540 125944
rect 246960 3534 246988 126414
rect 248340 125662 248368 128166
rect 249260 126682 249288 128166
rect 249248 126676 249300 126682
rect 249248 126618 249300 126624
rect 250180 126614 250208 128166
rect 251008 126750 251036 128166
rect 251928 126886 251956 128166
rect 251916 126880 251968 126886
rect 251916 126822 251968 126828
rect 250996 126744 251048 126750
rect 250996 126686 251048 126692
rect 250444 126676 250496 126682
rect 250444 126618 250496 126624
rect 250168 126608 250220 126614
rect 250168 126550 250220 126556
rect 249064 126540 249116 126546
rect 249064 126482 249116 126488
rect 248328 125656 248380 125662
rect 248328 125598 248380 125604
rect 249076 3602 249104 126482
rect 249156 125656 249208 125662
rect 249156 125598 249208 125604
rect 249168 4078 249196 125598
rect 249156 4072 249208 4078
rect 249156 4014 249208 4020
rect 247592 3596 247644 3602
rect 247592 3538 247644 3544
rect 249064 3596 249116 3602
rect 249064 3538 249116 3544
rect 246396 3528 246448 3534
rect 246396 3470 246448 3476
rect 246948 3528 247000 3534
rect 246948 3470 247000 3476
rect 246304 3188 246356 3194
rect 246304 3130 246356 3136
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245396 462 245608 490
rect 246408 480 246436 3470
rect 247604 480 247632 3538
rect 250456 3534 250484 126618
rect 252468 126608 252520 126614
rect 252468 126550 252520 126556
rect 251824 126200 251876 126206
rect 251824 126142 251876 126148
rect 248788 3528 248840 3534
rect 248788 3470 248840 3476
rect 250444 3528 250496 3534
rect 250444 3470 250496 3476
rect 248800 480 248828 3470
rect 251180 3460 251232 3466
rect 251180 3402 251232 3408
rect 249984 3052 250036 3058
rect 249984 2994 250036 3000
rect 249996 480 250024 2994
rect 251192 480 251220 3402
rect 251836 3058 251864 126142
rect 252376 3528 252428 3534
rect 252376 3470 252428 3476
rect 251824 3052 251876 3058
rect 251824 2994 251876 3000
rect 252388 480 252416 3470
rect 252480 3466 252508 126550
rect 252848 126342 252876 128166
rect 253768 126818 253796 128166
rect 253756 126812 253808 126818
rect 253756 126754 253808 126760
rect 253204 126744 253256 126750
rect 253204 126686 253256 126692
rect 252836 126336 252888 126342
rect 252836 126278 252888 126284
rect 253216 3534 253244 126686
rect 254688 125662 254716 128166
rect 255228 126336 255280 126342
rect 255228 126278 255280 126284
rect 254676 125656 254728 125662
rect 254676 125598 254728 125604
rect 253480 4072 253532 4078
rect 253480 4014 253532 4020
rect 253204 3528 253256 3534
rect 253204 3470 253256 3476
rect 252468 3460 252520 3466
rect 252468 3402 252520 3408
rect 253492 480 253520 4014
rect 255240 3534 255268 126278
rect 255608 126274 255636 128166
rect 256528 126410 256556 128166
rect 256608 126812 256660 126818
rect 256608 126754 256660 126760
rect 256516 126404 256568 126410
rect 256516 126346 256568 126352
rect 255596 126268 255648 126274
rect 255596 126210 255648 126216
rect 256620 3534 256648 126754
rect 257356 126478 257384 128166
rect 258276 126546 258304 128166
rect 259196 126682 259224 128166
rect 259184 126676 259236 126682
rect 259184 126618 259236 126624
rect 258264 126540 258316 126546
rect 258264 126482 258316 126488
rect 257344 126472 257396 126478
rect 257344 126414 257396 126420
rect 260116 126206 260144 128166
rect 261036 126614 261064 128166
rect 261956 126750 261984 128166
rect 261944 126744 261996 126750
rect 261944 126686 261996 126692
rect 261024 126608 261076 126614
rect 261024 126550 261076 126556
rect 260748 126404 260800 126410
rect 260748 126346 260800 126352
rect 260104 126200 260156 126206
rect 260104 126142 260156 126148
rect 260104 125996 260156 126002
rect 260104 125938 260156 125944
rect 259368 125792 259420 125798
rect 259368 125734 259420 125740
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 255228 3528 255280 3534
rect 255228 3470 255280 3476
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 256608 3528 256660 3534
rect 256608 3470 256660 3476
rect 257068 3528 257120 3534
rect 257068 3470 257120 3476
rect 254688 480 254716 3470
rect 255884 480 255912 3470
rect 257080 480 257108 3470
rect 259380 3262 259408 125734
rect 260116 4078 260144 125938
rect 260760 6914 260788 126346
rect 262876 126002 262904 128166
rect 263704 126342 263732 128166
rect 264624 126818 264652 128166
rect 264612 126812 264664 126818
rect 264612 126754 264664 126760
rect 263692 126336 263744 126342
rect 263692 126278 263744 126284
rect 262864 125996 262916 126002
rect 262864 125938 262916 125944
rect 262864 125860 262916 125866
rect 262864 125802 262916 125808
rect 260668 6886 260788 6914
rect 260104 4072 260156 4078
rect 260104 4014 260156 4020
rect 259460 3460 259512 3466
rect 259460 3402 259512 3408
rect 258264 3256 258316 3262
rect 258264 3198 258316 3204
rect 259368 3256 259420 3262
rect 259368 3198 259420 3204
rect 258276 480 258304 3198
rect 259472 480 259500 3402
rect 260668 480 260696 6886
rect 262876 3534 262904 125802
rect 264244 125724 264296 125730
rect 264244 125666 264296 125672
rect 262956 125656 263008 125662
rect 262956 125598 263008 125604
rect 262968 3602 262996 125598
rect 262956 3596 263008 3602
rect 262956 3538 263008 3544
rect 261760 3528 261812 3534
rect 261760 3470 261812 3476
rect 262864 3528 262916 3534
rect 262864 3470 262916 3476
rect 261772 480 261800 3470
rect 264256 3466 264284 125666
rect 265544 125662 265572 128166
rect 266464 125798 266492 128166
rect 267004 126268 267056 126274
rect 267004 126210 267056 126216
rect 266452 125792 266504 125798
rect 266452 125734 266504 125740
rect 265532 125656 265584 125662
rect 265532 125598 265584 125604
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 264244 3460 264296 3466
rect 264244 3402 264296 3408
rect 265348 3460 265400 3466
rect 265348 3402 265400 3408
rect 262956 3324 263008 3330
rect 262956 3266 263008 3272
rect 262968 480 262996 3266
rect 264152 2984 264204 2990
rect 264152 2926 264204 2932
rect 264164 480 264192 2926
rect 265360 480 265388 3402
rect 266556 480 266584 3470
rect 267016 3466 267044 126210
rect 267384 125730 267412 128166
rect 267648 126540 267700 126546
rect 267648 126482 267700 126488
rect 267372 125724 267424 125730
rect 267372 125666 267424 125672
rect 267660 3534 267688 126482
rect 268304 126410 268332 128166
rect 268292 126404 268344 126410
rect 268292 126346 268344 126352
rect 269224 125866 269252 128166
rect 269212 125860 269264 125866
rect 269212 125802 269264 125808
rect 269028 125792 269080 125798
rect 269028 125734 269080 125740
rect 268384 125656 268436 125662
rect 268384 125598 268436 125604
rect 267648 3528 267700 3534
rect 267648 3470 267700 3476
rect 267740 3528 267792 3534
rect 267740 3470 267792 3476
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 267752 480 267780 3470
rect 268396 2990 268424 125598
rect 269040 3534 269068 125734
rect 269028 3528 269080 3534
rect 269028 3470 269080 3476
rect 269408 3330 269436 128166
rect 270408 125860 270460 125866
rect 270408 125802 270460 125808
rect 269396 3324 269448 3330
rect 269396 3266 269448 3272
rect 268384 2984 268436 2990
rect 268384 2926 268436 2932
rect 268844 2916 268896 2922
rect 268844 2858 268896 2864
rect 268856 480 268884 2858
rect 270052 598 270264 626
rect 270052 480 270080 598
rect 270236 490 270264 598
rect 270420 490 270448 125802
rect 270972 125662 271000 128166
rect 271892 126274 271920 128166
rect 272812 126546 272840 128166
rect 272800 126540 272852 126546
rect 272800 126482 272852 126488
rect 271880 126268 271932 126274
rect 271880 126210 271932 126216
rect 273732 125798 273760 128166
rect 273996 126268 274048 126274
rect 273996 126210 274048 126216
rect 273720 125792 273772 125798
rect 273720 125734 273772 125740
rect 271788 125724 271840 125730
rect 271788 125666 271840 125672
rect 270960 125656 271012 125662
rect 270960 125598 271012 125604
rect 271800 3534 271828 125666
rect 273904 125656 273956 125662
rect 273904 125598 273956 125604
rect 273628 4072 273680 4078
rect 273628 4014 273680 4020
rect 271236 3528 271288 3534
rect 271236 3470 271288 3476
rect 271788 3528 271840 3534
rect 271788 3470 271840 3476
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270236 462 270448 490
rect 271248 480 271276 3470
rect 272432 3052 272484 3058
rect 272432 2994 272484 3000
rect 272444 480 272472 2994
rect 273640 480 273668 4014
rect 273916 2922 273944 125598
rect 274008 3058 274036 126210
rect 274652 125662 274680 128166
rect 275572 125866 275600 128166
rect 275560 125860 275612 125866
rect 275560 125802 275612 125808
rect 276400 125730 276428 128166
rect 276664 126948 276716 126954
rect 276664 126890 276716 126896
rect 276388 125724 276440 125730
rect 276388 125666 276440 125672
rect 274640 125656 274692 125662
rect 274640 125598 274692 125604
rect 276020 3528 276072 3534
rect 276020 3470 276072 3476
rect 273996 3052 274048 3058
rect 273996 2994 274048 3000
rect 274824 3052 274876 3058
rect 274824 2994 274876 3000
rect 273904 2916 273956 2922
rect 273904 2858 273956 2864
rect 274836 480 274864 2994
rect 276032 480 276060 3470
rect 276676 3058 276704 126890
rect 277320 126274 277348 128166
rect 277308 126268 277360 126274
rect 277308 126210 277360 126216
rect 277308 126132 277360 126138
rect 277308 126074 277360 126080
rect 277124 3664 277176 3670
rect 277124 3606 277176 3612
rect 276664 3052 276716 3058
rect 276664 2994 276716 3000
rect 277136 480 277164 3606
rect 277320 3534 277348 126074
rect 277504 4078 277532 128166
rect 279160 126954 279188 128166
rect 279148 126948 279200 126954
rect 279148 126890 279200 126896
rect 280080 126138 280108 128166
rect 280068 126132 280120 126138
rect 280068 126074 280120 126080
rect 278688 125656 278740 125662
rect 278688 125598 278740 125604
rect 277492 4072 277544 4078
rect 277492 4014 277544 4020
rect 277308 3528 277360 3534
rect 277308 3470 277360 3476
rect 278332 598 278544 626
rect 278332 480 278360 598
rect 278516 490 278544 598
rect 278700 490 278728 125598
rect 280356 3670 280384 128166
rect 280804 125724 280856 125730
rect 280804 125666 280856 125672
rect 280344 3664 280396 3670
rect 280344 3606 280396 3612
rect 280816 3398 280844 125666
rect 281920 125662 281948 128166
rect 282748 125730 282776 128166
rect 282736 125724 282788 125730
rect 282736 125666 282788 125672
rect 282828 125724 282880 125730
rect 282828 125666 282880 125672
rect 281908 125656 281960 125662
rect 281908 125598 281960 125604
rect 282184 125656 282236 125662
rect 282184 125598 282236 125604
rect 281908 3528 281960 3534
rect 281908 3470 281960 3476
rect 279516 3392 279568 3398
rect 279516 3334 279568 3340
rect 280804 3392 280856 3398
rect 280804 3334 280856 3340
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 278516 462 278728 490
rect 279528 480 279556 3334
rect 280712 3188 280764 3194
rect 280712 3130 280764 3136
rect 280724 480 280752 3130
rect 281920 480 281948 3470
rect 282196 3194 282224 125598
rect 282840 3534 282868 125666
rect 283668 125662 283696 128166
rect 284404 125730 284432 128302
rect 285554 128194 285582 128452
rect 286474 128194 286502 128452
rect 284496 128166 285582 128194
rect 285692 128166 286502 128194
rect 287152 128240 287204 128246
rect 287394 128194 287422 128452
rect 288314 128246 288342 128452
rect 287152 128182 287204 128188
rect 284392 125724 284444 125730
rect 284392 125666 284444 125672
rect 283656 125656 283708 125662
rect 283656 125598 283708 125604
rect 284496 3534 284524 128166
rect 285588 126812 285640 126818
rect 285588 126754 285640 126760
rect 285600 6914 285628 126754
rect 285416 6886 285628 6914
rect 282828 3528 282880 3534
rect 282828 3470 282880 3476
rect 283104 3528 283156 3534
rect 283104 3470 283156 3476
rect 284484 3528 284536 3534
rect 284484 3470 284536 3476
rect 282184 3188 282236 3194
rect 282184 3130 282236 3136
rect 283116 480 283144 3470
rect 284300 2916 284352 2922
rect 284300 2858 284352 2864
rect 284312 480 284340 2858
rect 285416 480 285444 6886
rect 285692 2922 285720 128166
rect 287164 4146 287192 128182
rect 287348 128166 287422 128194
rect 288302 128240 288354 128246
rect 289142 128194 289170 128452
rect 290062 128194 290090 128452
rect 290982 128194 291010 128452
rect 291902 128194 291930 128452
rect 292822 128194 292850 128452
rect 293742 128194 293770 128452
rect 294662 128194 294690 128452
rect 295582 128194 295610 128452
rect 288302 128182 288354 128188
rect 289096 128166 289170 128194
rect 289832 128166 290090 128194
rect 290936 128166 291010 128194
rect 291212 128166 291930 128194
rect 292684 128166 292850 128194
rect 293696 128166 293770 128194
rect 293972 128166 294690 128194
rect 295352 128166 295610 128194
rect 296410 128194 296438 128452
rect 297330 128194 297358 128452
rect 298250 128194 298278 128452
rect 299170 128194 299198 128452
rect 300090 128194 300118 128452
rect 301010 128194 301038 128452
rect 301930 128194 301958 128452
rect 302758 128194 302786 128452
rect 303678 128194 303706 128452
rect 304598 128194 304626 128452
rect 305518 128194 305546 128452
rect 306438 128194 306466 128452
rect 307358 128194 307386 128452
rect 308278 128194 308306 128452
rect 309106 128194 309134 128452
rect 296410 128166 296668 128194
rect 297330 128166 297404 128194
rect 298250 128166 298324 128194
rect 299170 128166 299428 128194
rect 300090 128166 300164 128194
rect 301010 128166 301084 128194
rect 301930 128166 302004 128194
rect 302758 128166 302832 128194
rect 303678 128166 303752 128194
rect 304598 128166 304948 128194
rect 305518 128166 305592 128194
rect 306438 128166 306512 128194
rect 307358 128166 307708 128194
rect 308278 128166 308352 128194
rect 287348 126818 287376 128166
rect 287336 126812 287388 126818
rect 287336 126754 287388 126760
rect 289096 125662 289124 128166
rect 288348 125656 288400 125662
rect 288348 125598 288400 125604
rect 289084 125656 289136 125662
rect 289832 125610 289860 128166
rect 290936 125662 290964 128166
rect 289084 125598 289136 125604
rect 286600 4140 286652 4146
rect 286600 4082 286652 4088
rect 287152 4140 287204 4146
rect 287152 4082 287204 4088
rect 285680 2916 285732 2922
rect 285680 2858 285732 2864
rect 286612 480 286640 4082
rect 288360 3330 288388 125598
rect 289740 125582 289860 125610
rect 289912 125656 289964 125662
rect 289912 125598 289964 125604
rect 290924 125656 290976 125662
rect 290924 125598 290976 125604
rect 289740 3534 289768 125582
rect 289924 122834 289952 125598
rect 289832 122806 289952 122834
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 287796 3324 287848 3330
rect 287796 3266 287848 3272
rect 288348 3324 288400 3330
rect 288348 3266 288400 3272
rect 287808 480 287836 3266
rect 289004 480 289032 3470
rect 289832 490 289860 122806
rect 291212 16574 291240 128166
rect 292580 125656 292632 125662
rect 292580 125598 292632 125604
rect 291212 16546 291424 16574
rect 290016 598 290228 626
rect 290016 490 290044 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 462 290044 490
rect 290200 480 290228 598
rect 291396 480 291424 16546
rect 292592 3602 292620 125598
rect 292580 3596 292632 3602
rect 292580 3538 292632 3544
rect 292684 3482 292712 128166
rect 293696 125662 293724 128166
rect 293684 125656 293736 125662
rect 293684 125598 293736 125604
rect 293684 3596 293736 3602
rect 293684 3538 293736 3544
rect 292592 3454 292712 3482
rect 292592 480 292620 3454
rect 293696 480 293724 3538
rect 293972 3534 294000 128166
rect 295352 3534 295380 128166
rect 296640 4146 296668 128166
rect 297376 125662 297404 128166
rect 298296 125662 298324 128166
rect 297364 125656 297416 125662
rect 297364 125598 297416 125604
rect 298100 125656 298152 125662
rect 298100 125598 298152 125604
rect 298284 125656 298336 125662
rect 298284 125598 298336 125604
rect 299296 125656 299348 125662
rect 299400 125644 299428 128166
rect 300136 125662 300164 128166
rect 301056 125662 301084 128166
rect 301976 125730 302004 128166
rect 301964 125724 302016 125730
rect 301964 125666 302016 125672
rect 302804 125662 302832 128166
rect 303724 126274 303752 128166
rect 303712 126268 303764 126274
rect 303712 126210 303764 126216
rect 303620 125724 303672 125730
rect 303620 125666 303672 125672
rect 300124 125656 300176 125662
rect 299400 125616 299612 125644
rect 299296 125598 299348 125604
rect 296628 4140 296680 4146
rect 296628 4082 296680 4088
rect 297272 4140 297324 4146
rect 297272 4082 297324 4088
rect 293960 3528 294012 3534
rect 293960 3470 294012 3476
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 295340 3528 295392 3534
rect 295340 3470 295392 3476
rect 296076 3528 296128 3534
rect 296076 3470 296128 3476
rect 294892 480 294920 3470
rect 296088 480 296116 3470
rect 297284 480 297312 4082
rect 298112 490 298140 125598
rect 299308 122834 299336 125598
rect 299308 122806 299428 122834
rect 299400 3482 299428 122806
rect 299584 16574 299612 125616
rect 300124 125598 300176 125604
rect 300768 125656 300820 125662
rect 300768 125598 300820 125604
rect 301044 125656 301096 125662
rect 301044 125598 301096 125604
rect 302240 125656 302292 125662
rect 302240 125598 302292 125604
rect 302792 125656 302844 125662
rect 302792 125598 302844 125604
rect 299584 16546 300716 16574
rect 299400 3454 299704 3482
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3454
rect 300688 3346 300716 16546
rect 300780 3534 300808 125598
rect 302252 16574 302280 125598
rect 303632 16574 303660 125666
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 301964 3528 302016 3534
rect 301964 3470 302016 3476
rect 300688 3318 300808 3346
rect 300780 480 300808 3318
rect 301976 480 302004 3470
rect 303172 480 303200 16546
rect 303908 490 303936 16546
rect 304920 4146 304948 128166
rect 305564 125662 305592 128166
rect 306380 126268 306432 126274
rect 306380 126210 306432 126216
rect 305000 125656 305052 125662
rect 305000 125598 305052 125604
rect 305552 125656 305604 125662
rect 305552 125598 305604 125604
rect 306288 125656 306340 125662
rect 306288 125598 306340 125604
rect 305012 16574 305040 125598
rect 305012 16546 305592 16574
rect 304908 4140 304960 4146
rect 304908 4082 304960 4088
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 16546
rect 306300 3466 306328 125598
rect 306288 3460 306340 3466
rect 306288 3402 306340 3408
rect 306392 490 306420 126210
rect 306484 125662 306512 128166
rect 306472 125656 306524 125662
rect 306472 125598 306524 125604
rect 307680 3262 307708 128166
rect 308324 125730 308352 128166
rect 309060 128166 309134 128194
rect 310026 128194 310054 128452
rect 310946 128194 310974 128452
rect 311866 128194 311894 128452
rect 310026 128166 310468 128194
rect 310946 128166 311020 128194
rect 309060 125798 309088 128166
rect 309048 125792 309100 125798
rect 309048 125734 309100 125740
rect 308312 125724 308364 125730
rect 308312 125666 308364 125672
rect 309140 125656 309192 125662
rect 309140 125598 309192 125604
rect 309152 16574 309180 125598
rect 309152 16546 309824 16574
rect 307944 4140 307996 4146
rect 307944 4082 307996 4088
rect 307668 3256 307720 3262
rect 307668 3198 307720 3204
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 4082
rect 309048 3460 309100 3466
rect 309048 3402 309100 3408
rect 309060 480 309088 3402
rect 309796 490 309824 16546
rect 310440 3330 310468 128166
rect 310992 125662 311020 128166
rect 311820 128166 311894 128194
rect 312786 128194 312814 128452
rect 313706 128194 313734 128452
rect 314626 128194 314654 128452
rect 312786 128166 312860 128194
rect 313706 128166 313780 128194
rect 310980 125656 311032 125662
rect 310980 125598 311032 125604
rect 311716 125656 311768 125662
rect 311716 125598 311768 125604
rect 310428 3324 310480 3330
rect 310428 3266 310480 3272
rect 311440 3256 311492 3262
rect 311440 3198 311492 3204
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 3198
rect 311728 3194 311756 125598
rect 311820 3398 311848 128166
rect 312832 126886 312860 128166
rect 312820 126880 312872 126886
rect 312820 126822 312872 126828
rect 313280 125792 313332 125798
rect 313280 125734 313332 125740
rect 311900 125724 311952 125730
rect 311900 125666 311952 125672
rect 311912 16574 311940 125666
rect 313292 16574 313320 125734
rect 313752 125662 313780 128166
rect 314580 128166 314654 128194
rect 315454 128194 315482 128452
rect 316374 128194 316402 128452
rect 317294 128194 317322 128452
rect 318214 128194 318242 128452
rect 319134 128194 319162 128452
rect 320054 128194 320082 128452
rect 320974 128194 321002 128452
rect 321802 128194 321830 128452
rect 322722 128194 322750 128452
rect 323642 128194 323670 128452
rect 324562 128194 324590 128452
rect 325482 128194 325510 128452
rect 326402 128194 326430 128452
rect 327322 128194 327350 128452
rect 328150 128194 328178 128452
rect 329070 128194 329098 128452
rect 329990 128194 330018 128452
rect 330910 128194 330938 128452
rect 331830 128194 331858 128452
rect 332750 128194 332778 128452
rect 333670 128194 333698 128452
rect 334498 128194 334526 128452
rect 335418 128194 335446 128452
rect 336338 128194 336366 128452
rect 337258 128194 337286 128452
rect 338178 128194 338206 128452
rect 339098 128194 339126 128452
rect 340018 128194 340046 128452
rect 340938 128194 340966 128452
rect 341766 128194 341794 128452
rect 342686 128194 342714 128452
rect 343606 128194 343634 128452
rect 315454 128166 315528 128194
rect 316374 128166 316448 128194
rect 317294 128166 317368 128194
rect 318214 128166 318288 128194
rect 319134 128166 319208 128194
rect 320054 128166 320128 128194
rect 320974 128166 321048 128194
rect 321802 128166 321876 128194
rect 322722 128166 322796 128194
rect 323642 128166 323716 128194
rect 324562 128166 324636 128194
rect 325482 128166 325648 128194
rect 326402 128166 326476 128194
rect 327322 128166 327396 128194
rect 328150 128166 328316 128194
rect 329070 128166 329144 128194
rect 329990 128166 330064 128194
rect 330910 128166 331076 128194
rect 331830 128166 331904 128194
rect 332750 128166 332824 128194
rect 333670 128166 333744 128194
rect 334498 128166 334572 128194
rect 335418 128166 335492 128194
rect 336338 128166 336688 128194
rect 337258 128166 337332 128194
rect 338178 128166 338252 128194
rect 339098 128166 339448 128194
rect 340018 128166 340092 128194
rect 340938 128166 341012 128194
rect 341766 128166 342208 128194
rect 342686 128166 342760 128194
rect 313740 125656 313792 125662
rect 313740 125598 313792 125604
rect 314476 125656 314528 125662
rect 314476 125598 314528 125604
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 311808 3392 311860 3398
rect 311808 3334 311860 3340
rect 311716 3188 311768 3194
rect 311716 3130 311768 3136
rect 312188 490 312216 16546
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 314488 3602 314516 125598
rect 314476 3596 314528 3602
rect 314476 3538 314528 3544
rect 314580 3466 314608 128166
rect 315500 126274 315528 128166
rect 315488 126268 315540 126274
rect 315488 126210 315540 126216
rect 316420 125662 316448 128166
rect 316408 125656 316460 125662
rect 316408 125598 316460 125604
rect 317236 125656 317288 125662
rect 317236 125598 317288 125604
rect 314568 3460 314620 3466
rect 314568 3402 314620 3408
rect 315028 3324 315080 3330
rect 315028 3266 315080 3272
rect 315040 480 315068 3266
rect 317248 3262 317276 125598
rect 317340 3738 317368 128166
rect 317420 126880 317472 126886
rect 317420 126822 317472 126828
rect 317432 6914 317460 126822
rect 318064 126268 318116 126274
rect 318064 126210 318116 126216
rect 318076 16574 318104 126210
rect 318260 125662 318288 128166
rect 319180 125730 319208 128166
rect 319168 125724 319220 125730
rect 319168 125666 319220 125672
rect 320100 125662 320128 128166
rect 321020 125662 321048 128166
rect 321848 125662 321876 128166
rect 322204 125724 322256 125730
rect 322204 125666 322256 125672
rect 318248 125656 318300 125662
rect 318248 125598 318300 125604
rect 318708 125656 318760 125662
rect 318708 125598 318760 125604
rect 320088 125656 320140 125662
rect 320088 125598 320140 125604
rect 320824 125656 320876 125662
rect 320824 125598 320876 125604
rect 321008 125656 321060 125662
rect 321008 125598 321060 125604
rect 321468 125656 321520 125662
rect 321468 125598 321520 125604
rect 321836 125656 321888 125662
rect 321836 125598 321888 125604
rect 318076 16546 318196 16574
rect 317432 6886 318104 6914
rect 317328 3732 317380 3738
rect 317328 3674 317380 3680
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317236 3256 317288 3262
rect 317236 3198 317288 3204
rect 316224 3188 316276 3194
rect 316224 3130 316276 3136
rect 316236 480 316264 3130
rect 317340 480 317368 3334
rect 318076 490 318104 6886
rect 318168 3534 318196 16546
rect 318156 3528 318208 3534
rect 318156 3470 318208 3476
rect 318720 3398 318748 125598
rect 319720 3596 319772 3602
rect 319720 3538 319772 3544
rect 318708 3392 318760 3398
rect 318708 3334 318760 3340
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 3538
rect 320836 3330 320864 125598
rect 321480 3670 321508 125598
rect 321468 3664 321520 3670
rect 321468 3606 321520 3612
rect 322112 3528 322164 3534
rect 322112 3470 322164 3476
rect 320916 3460 320968 3466
rect 320916 3402 320968 3408
rect 320824 3324 320876 3330
rect 320824 3266 320876 3272
rect 320928 480 320956 3402
rect 322124 480 322152 3470
rect 322216 3058 322244 125666
rect 322768 3466 322796 128166
rect 323688 125662 323716 128166
rect 324608 125662 324636 128166
rect 322848 125656 322900 125662
rect 322848 125598 322900 125604
rect 323676 125656 323728 125662
rect 323676 125598 323728 125604
rect 324228 125656 324280 125662
rect 324228 125598 324280 125604
rect 324596 125656 324648 125662
rect 324596 125598 324648 125604
rect 325516 125656 325568 125662
rect 325516 125598 325568 125604
rect 322860 3806 322888 125598
rect 324240 4010 324268 125598
rect 325528 4078 325556 125598
rect 325516 4072 325568 4078
rect 325516 4014 325568 4020
rect 324228 4004 324280 4010
rect 324228 3946 324280 3952
rect 322848 3800 322900 3806
rect 322848 3742 322900 3748
rect 324412 3732 324464 3738
rect 324412 3674 324464 3680
rect 322756 3460 322808 3466
rect 322756 3402 322808 3408
rect 323308 3256 323360 3262
rect 323308 3198 323360 3204
rect 322204 3052 322256 3058
rect 322204 2994 322256 3000
rect 323320 480 323348 3198
rect 324424 480 324452 3674
rect 325620 3534 325648 128166
rect 326448 125730 326476 128166
rect 326436 125724 326488 125730
rect 326436 125666 326488 125672
rect 327368 125662 327396 128166
rect 327356 125656 327408 125662
rect 327356 125598 327408 125604
rect 328288 3602 328316 128166
rect 329116 125662 329144 128166
rect 330036 125662 330064 128166
rect 328368 125656 328420 125662
rect 328368 125598 328420 125604
rect 329104 125656 329156 125662
rect 329104 125598 329156 125604
rect 329748 125656 329800 125662
rect 329748 125598 329800 125604
rect 330024 125656 330076 125662
rect 330024 125598 330076 125604
rect 328380 3942 328408 125598
rect 328368 3936 328420 3942
rect 328368 3878 328420 3884
rect 329760 3738 329788 125598
rect 330392 3800 330444 3806
rect 330392 3742 330444 3748
rect 329748 3732 329800 3738
rect 329748 3674 329800 3680
rect 329196 3664 329248 3670
rect 329196 3606 329248 3612
rect 328276 3596 328328 3602
rect 328276 3538 328328 3544
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 328000 3324 328052 3330
rect 328000 3266 328052 3272
rect 326804 3052 326856 3058
rect 326804 2994 326856 3000
rect 326816 480 326844 2994
rect 328012 480 328040 3266
rect 329208 480 329236 3606
rect 330404 480 330432 3742
rect 331048 3670 331076 128166
rect 331772 125724 331824 125730
rect 331772 125666 331824 125672
rect 331128 125656 331180 125662
rect 331128 125598 331180 125604
rect 331140 3806 331168 125598
rect 331784 122834 331812 125666
rect 331876 125662 331904 128166
rect 332796 126410 332824 128166
rect 332784 126404 332836 126410
rect 332784 126346 332836 126352
rect 333716 125730 333744 128166
rect 333704 125724 333756 125730
rect 333704 125666 333756 125672
rect 334544 125662 334572 128166
rect 334624 125724 334676 125730
rect 334624 125666 334676 125672
rect 331864 125656 331916 125662
rect 331864 125598 331916 125604
rect 332508 125656 332560 125662
rect 332508 125598 332560 125604
rect 334532 125656 334584 125662
rect 334532 125598 334584 125604
rect 331784 122806 331904 122834
rect 331876 4146 331904 122806
rect 331864 4140 331916 4146
rect 331864 4082 331916 4088
rect 332520 3874 332548 125598
rect 333888 4072 333940 4078
rect 333888 4014 333940 4020
rect 332692 4004 332744 4010
rect 332692 3946 332744 3952
rect 332508 3868 332560 3874
rect 332508 3810 332560 3816
rect 331128 3800 331180 3806
rect 331128 3742 331180 3748
rect 331036 3664 331088 3670
rect 331036 3606 331088 3612
rect 331588 3460 331640 3466
rect 331588 3402 331640 3408
rect 331600 480 331628 3402
rect 332704 480 332732 3946
rect 333900 480 333928 4014
rect 334636 3466 334664 125666
rect 335464 125662 335492 128166
rect 336004 126404 336056 126410
rect 336004 126346 336056 126352
rect 335268 125656 335320 125662
rect 335268 125598 335320 125604
rect 335452 125656 335504 125662
rect 335452 125598 335504 125604
rect 335084 3528 335136 3534
rect 335084 3470 335136 3476
rect 334624 3460 334676 3466
rect 334624 3402 334676 3408
rect 335096 480 335124 3470
rect 335280 3330 335308 125598
rect 335268 3324 335320 3330
rect 335268 3266 335320 3272
rect 336016 2922 336044 126346
rect 336556 125656 336608 125662
rect 336556 125598 336608 125604
rect 336280 4140 336332 4146
rect 336280 4082 336332 4088
rect 336004 2916 336056 2922
rect 336004 2858 336056 2864
rect 336292 480 336320 4082
rect 336568 3466 336596 125598
rect 336660 4146 336688 128166
rect 337304 125730 337332 128166
rect 337292 125724 337344 125730
rect 337292 125666 337344 125672
rect 338224 125662 338252 128166
rect 338212 125656 338264 125662
rect 338212 125598 338264 125604
rect 339316 125656 339368 125662
rect 339316 125598 339368 125604
rect 336648 4140 336700 4146
rect 336648 4082 336700 4088
rect 337476 3936 337528 3942
rect 337476 3878 337528 3884
rect 336556 3460 336608 3466
rect 336556 3402 336608 3408
rect 337488 480 337516 3878
rect 338672 3596 338724 3602
rect 338672 3538 338724 3544
rect 338684 480 338712 3538
rect 339328 3398 339356 125598
rect 339420 4078 339448 128166
rect 340064 125662 340092 128166
rect 340144 125724 340196 125730
rect 340144 125666 340196 125672
rect 340052 125656 340104 125662
rect 340052 125598 340104 125604
rect 339408 4072 339460 4078
rect 339408 4014 339460 4020
rect 339868 3732 339920 3738
rect 339868 3674 339920 3680
rect 339316 3392 339368 3398
rect 339316 3334 339368 3340
rect 339880 480 339908 3674
rect 340156 3262 340184 125666
rect 340984 125662 341012 128166
rect 340788 125656 340840 125662
rect 340788 125598 340840 125604
rect 340972 125656 341024 125662
rect 340972 125598 341024 125604
rect 342076 125656 342128 125662
rect 342076 125598 342128 125604
rect 340800 3738 340828 125598
rect 342088 4010 342116 125598
rect 342076 4004 342128 4010
rect 342076 3946 342128 3952
rect 342180 3806 342208 128166
rect 342732 125662 342760 128166
rect 343468 128166 343634 128194
rect 344526 128194 344554 128452
rect 345446 128194 345474 128452
rect 346366 128194 346394 128452
rect 344526 128166 344600 128194
rect 345446 128166 345520 128194
rect 342720 125656 342772 125662
rect 342720 125598 342772 125604
rect 343364 3868 343416 3874
rect 343364 3810 343416 3816
rect 340972 3800 341024 3806
rect 340972 3742 341024 3748
rect 342168 3800 342220 3806
rect 342168 3742 342220 3748
rect 340788 3732 340840 3738
rect 340788 3674 340840 3680
rect 340144 3256 340196 3262
rect 340144 3198 340196 3204
rect 340984 480 341012 3742
rect 342168 3664 342220 3670
rect 342168 3606 342220 3612
rect 342180 480 342208 3606
rect 343376 480 343404 3810
rect 343468 3602 343496 128166
rect 344572 126954 344600 128166
rect 344560 126948 344612 126954
rect 344560 126890 344612 126896
rect 345492 125662 345520 128166
rect 346228 128166 346394 128194
rect 347286 128194 347314 128452
rect 348114 128194 348142 128452
rect 349034 128194 349062 128452
rect 349954 128194 349982 128452
rect 350874 128194 350902 128452
rect 351794 128194 351822 128452
rect 352714 128194 352742 128452
rect 353634 128194 353662 128452
rect 354462 128194 354490 128452
rect 355382 128194 355410 128452
rect 356302 128194 356330 128452
rect 357222 128194 357250 128452
rect 358142 128194 358170 128452
rect 359062 128194 359090 128452
rect 359982 128194 360010 128452
rect 360810 128194 360838 128452
rect 361730 128194 361758 128452
rect 362650 128194 362678 128452
rect 363570 128194 363598 128452
rect 364490 128194 364518 128452
rect 365410 128194 365438 128452
rect 366330 128194 366358 128452
rect 367158 128194 367186 128452
rect 368078 128194 368106 128452
rect 368998 128194 369026 128452
rect 369918 128194 369946 128452
rect 370838 128194 370866 128452
rect 371758 128194 371786 128452
rect 372678 128194 372706 128452
rect 373506 128194 373534 128452
rect 374426 128194 374454 128452
rect 375346 128194 375374 128452
rect 347286 128166 347728 128194
rect 348114 128166 348188 128194
rect 349034 128166 349108 128194
rect 349954 128166 350028 128194
rect 350874 128166 350948 128194
rect 351794 128166 351868 128194
rect 352714 128166 352788 128194
rect 353634 128166 353708 128194
rect 354462 128166 354536 128194
rect 355382 128166 355456 128194
rect 356302 128166 356376 128194
rect 357222 128166 357296 128194
rect 358142 128166 358216 128194
rect 359062 128166 359136 128194
rect 359982 128166 360056 128194
rect 360810 128166 360884 128194
rect 361730 128166 361804 128194
rect 362650 128166 362816 128194
rect 363570 128166 363644 128194
rect 364490 128166 364564 128194
rect 365410 128166 365576 128194
rect 366330 128166 366404 128194
rect 367158 128166 367232 128194
rect 368078 128166 368336 128194
rect 368998 128166 369072 128194
rect 369918 128166 369992 128194
rect 370838 128166 371096 128194
rect 371758 128166 371832 128194
rect 372678 128166 372752 128194
rect 373506 128166 373856 128194
rect 374426 128166 374500 128194
rect 345664 126948 345716 126954
rect 345664 126890 345716 126896
rect 343548 125656 343600 125662
rect 343548 125598 343600 125604
rect 345480 125656 345532 125662
rect 345480 125598 345532 125604
rect 343560 3874 343588 125598
rect 345676 3942 345704 126890
rect 345664 3936 345716 3942
rect 345664 3878 345716 3884
rect 343548 3868 343600 3874
rect 343548 3810 343600 3816
rect 343456 3596 343508 3602
rect 343456 3538 343508 3544
rect 346228 3534 346256 128166
rect 346308 125656 346360 125662
rect 346308 125598 346360 125604
rect 346320 3670 346348 125598
rect 346308 3664 346360 3670
rect 346308 3606 346360 3612
rect 345756 3528 345808 3534
rect 345756 3470 345808 3476
rect 346216 3528 346268 3534
rect 346216 3470 346268 3476
rect 344560 2916 344612 2922
rect 344560 2858 344612 2864
rect 344572 480 344600 2858
rect 345768 480 345796 3470
rect 346952 3324 347004 3330
rect 346952 3266 347004 3272
rect 346964 480 346992 3266
rect 347700 3194 347728 128166
rect 348160 125730 348188 128166
rect 348148 125724 348200 125730
rect 348148 125666 348200 125672
rect 349080 3466 349108 128166
rect 350000 125662 350028 128166
rect 350920 126342 350948 128166
rect 350908 126336 350960 126342
rect 350908 126278 350960 126284
rect 349988 125656 350040 125662
rect 349988 125598 350040 125604
rect 350448 125656 350500 125662
rect 350448 125598 350500 125604
rect 350460 6914 350488 125598
rect 350368 6886 350488 6914
rect 349252 4140 349304 4146
rect 349252 4082 349304 4088
rect 348056 3460 348108 3466
rect 348056 3402 348108 3408
rect 349068 3460 349120 3466
rect 349068 3402 349120 3408
rect 347688 3188 347740 3194
rect 347688 3130 347740 3136
rect 348068 480 348096 3402
rect 349264 480 349292 4082
rect 350368 3126 350396 6886
rect 351644 3392 351696 3398
rect 351644 3334 351696 3340
rect 350448 3256 350500 3262
rect 350448 3198 350500 3204
rect 350356 3120 350408 3126
rect 350356 3062 350408 3068
rect 350460 480 350488 3198
rect 351656 480 351684 3334
rect 351840 3262 351868 128166
rect 352760 125662 352788 128166
rect 353680 125662 353708 128166
rect 353944 125724 353996 125730
rect 353944 125666 353996 125672
rect 352748 125656 352800 125662
rect 352748 125598 352800 125604
rect 353208 125656 353260 125662
rect 353208 125598 353260 125604
rect 353668 125656 353720 125662
rect 353668 125598 353720 125604
rect 352840 4072 352892 4078
rect 352840 4014 352892 4020
rect 351828 3256 351880 3262
rect 351828 3198 351880 3204
rect 352852 480 352880 4014
rect 353220 3398 353248 125598
rect 353208 3392 353260 3398
rect 353208 3334 353260 3340
rect 353956 3058 353984 125666
rect 354508 3738 354536 128166
rect 355428 125662 355456 128166
rect 356348 125730 356376 128166
rect 357268 126274 357296 128166
rect 357256 126268 357308 126274
rect 357256 126210 357308 126216
rect 356336 125724 356388 125730
rect 356336 125666 356388 125672
rect 357348 125724 357400 125730
rect 357348 125666 357400 125672
rect 354588 125656 354640 125662
rect 354588 125598 354640 125604
rect 355416 125656 355468 125662
rect 355416 125598 355468 125604
rect 356704 125656 356756 125662
rect 356704 125598 356756 125604
rect 354600 4078 354628 125598
rect 356716 4146 356744 125598
rect 356704 4140 356756 4146
rect 356704 4082 356756 4088
rect 354588 4072 354640 4078
rect 354588 4014 354640 4020
rect 355232 4004 355284 4010
rect 355232 3946 355284 3952
rect 354036 3732 354088 3738
rect 354036 3674 354088 3680
rect 354496 3732 354548 3738
rect 354496 3674 354548 3680
rect 353944 3052 353996 3058
rect 353944 2994 353996 3000
rect 354048 480 354076 3674
rect 355244 480 355272 3946
rect 356336 3800 356388 3806
rect 356336 3742 356388 3748
rect 356348 480 356376 3742
rect 357360 3330 357388 125666
rect 358188 125662 358216 128166
rect 359108 125662 359136 128166
rect 359464 126336 359516 126342
rect 359464 126278 359516 126284
rect 358176 125656 358228 125662
rect 358176 125598 358228 125604
rect 358728 125656 358780 125662
rect 358728 125598 358780 125604
rect 359096 125656 359148 125662
rect 359096 125598 359148 125604
rect 358740 3874 358768 125598
rect 357532 3868 357584 3874
rect 357532 3810 357584 3816
rect 358728 3868 358780 3874
rect 358728 3810 358780 3816
rect 357348 3324 357400 3330
rect 357348 3266 357400 3272
rect 357544 480 357572 3810
rect 358728 3596 358780 3602
rect 358728 3538 358780 3544
rect 358740 480 358768 3538
rect 359476 2854 359504 126278
rect 359924 3936 359976 3942
rect 359924 3878 359976 3884
rect 359464 2848 359516 2854
rect 359464 2790 359516 2796
rect 359936 480 359964 3878
rect 360028 3602 360056 128166
rect 360856 125662 360884 128166
rect 361776 125662 361804 128166
rect 360108 125656 360160 125662
rect 360108 125598 360160 125604
rect 360844 125656 360896 125662
rect 360844 125598 360896 125604
rect 361488 125656 361540 125662
rect 361488 125598 361540 125604
rect 361764 125656 361816 125662
rect 361764 125598 361816 125604
rect 360120 3942 360148 125598
rect 361500 4010 361528 125598
rect 361488 4004 361540 4010
rect 361488 3946 361540 3952
rect 360108 3936 360160 3942
rect 360108 3878 360160 3884
rect 362788 3670 362816 128166
rect 363616 125662 363644 128166
rect 364536 125662 364564 128166
rect 362868 125656 362920 125662
rect 362868 125598 362920 125604
rect 363604 125656 363656 125662
rect 363604 125598 363656 125604
rect 364248 125656 364300 125662
rect 364248 125598 364300 125604
rect 364524 125656 364576 125662
rect 364524 125598 364576 125604
rect 362880 3806 362908 125598
rect 362868 3800 362920 3806
rect 362868 3742 362920 3748
rect 361120 3664 361172 3670
rect 361120 3606 361172 3612
rect 362776 3664 362828 3670
rect 362776 3606 362828 3612
rect 360016 3596 360068 3602
rect 360016 3538 360068 3544
rect 361132 480 361160 3606
rect 362316 3528 362368 3534
rect 362316 3470 362368 3476
rect 362328 480 362356 3470
rect 363512 3188 363564 3194
rect 363512 3130 363564 3136
rect 363524 480 363552 3130
rect 364260 2922 364288 125598
rect 365548 3534 365576 128166
rect 366376 125662 366404 128166
rect 367204 125662 367232 128166
rect 365628 125656 365680 125662
rect 365628 125598 365680 125604
rect 366364 125656 366416 125662
rect 366364 125598 366416 125604
rect 367008 125656 367060 125662
rect 367008 125598 367060 125604
rect 367192 125656 367244 125662
rect 367192 125598 367244 125604
rect 365536 3528 365588 3534
rect 365536 3470 365588 3476
rect 364616 3052 364668 3058
rect 364616 2994 364668 3000
rect 364248 2916 364300 2922
rect 364248 2858 364300 2864
rect 364628 480 364656 2994
rect 365640 2990 365668 125598
rect 367020 6914 367048 125598
rect 366928 6886 367048 6914
rect 365812 3460 365864 3466
rect 365812 3402 365864 3408
rect 365628 2984 365680 2990
rect 365628 2926 365680 2932
rect 365824 480 365852 3402
rect 366928 3058 366956 6886
rect 368308 3466 368336 128166
rect 369044 125730 369072 128166
rect 369032 125724 369084 125730
rect 369032 125666 369084 125672
rect 369964 125662 369992 128166
rect 368388 125656 368440 125662
rect 368388 125598 368440 125604
rect 369952 125656 370004 125662
rect 369952 125598 370004 125604
rect 368296 3460 368348 3466
rect 368296 3402 368348 3408
rect 368400 3126 368428 125598
rect 371068 3398 371096 128166
rect 371804 125662 371832 128166
rect 371884 125724 371936 125730
rect 371884 125666 371936 125672
rect 371148 125656 371200 125662
rect 371148 125598 371200 125604
rect 371792 125656 371844 125662
rect 371792 125598 371844 125604
rect 370596 3392 370648 3398
rect 370596 3334 370648 3340
rect 371056 3392 371108 3398
rect 371056 3334 371108 3340
rect 369400 3256 369452 3262
rect 369400 3198 369452 3204
rect 367008 3120 367060 3126
rect 367008 3062 367060 3068
rect 368388 3120 368440 3126
rect 368388 3062 368440 3068
rect 366916 3052 366968 3058
rect 366916 2994 366968 3000
rect 367020 480 367048 3062
rect 368204 2848 368256 2854
rect 368204 2790 368256 2796
rect 368216 480 368244 2790
rect 369412 480 369440 3198
rect 370608 480 370636 3334
rect 371160 3194 371188 125598
rect 371896 4826 371924 125666
rect 372724 125662 372752 128166
rect 372528 125656 372580 125662
rect 372528 125598 372580 125604
rect 372712 125656 372764 125662
rect 372712 125598 372764 125604
rect 372540 7614 372568 125598
rect 372528 7608 372580 7614
rect 372528 7550 372580 7556
rect 371884 4820 371936 4826
rect 371884 4762 371936 4768
rect 373828 4078 373856 128166
rect 374472 125662 374500 128166
rect 375300 128166 375374 128194
rect 376266 128194 376294 128452
rect 377186 128194 377214 128452
rect 378106 128194 378134 128452
rect 376266 128166 376708 128194
rect 377186 128166 377260 128194
rect 373908 125656 373960 125662
rect 373908 125598 373960 125604
rect 374460 125656 374512 125662
rect 374460 125598 374512 125604
rect 375196 125656 375248 125662
rect 375196 125598 375248 125604
rect 371700 4072 371752 4078
rect 371700 4014 371752 4020
rect 373816 4072 373868 4078
rect 373816 4014 373868 4020
rect 371148 3188 371200 3194
rect 371148 3130 371200 3136
rect 371712 480 371740 4014
rect 372896 3732 372948 3738
rect 372896 3674 372948 3680
rect 372908 480 372936 3674
rect 373920 3262 373948 125598
rect 375208 4962 375236 125598
rect 375196 4956 375248 4962
rect 375196 4898 375248 4904
rect 375300 4146 375328 128166
rect 375380 126268 375432 126274
rect 375380 126210 375432 126216
rect 375392 16574 375420 126210
rect 375392 16546 376064 16574
rect 374092 4140 374144 4146
rect 374092 4082 374144 4088
rect 375288 4140 375340 4146
rect 375288 4082 375340 4088
rect 373908 3256 373960 3262
rect 373908 3198 373960 3204
rect 374104 480 374132 4082
rect 375288 3324 375340 3330
rect 375288 3266 375340 3272
rect 375300 480 375328 3266
rect 376036 490 376064 16546
rect 376680 3330 376708 128166
rect 377232 126342 377260 128166
rect 378060 128166 378134 128194
rect 379026 128194 379054 128452
rect 379854 128194 379882 128452
rect 380774 128194 380802 128452
rect 381694 128194 381722 128452
rect 382614 128194 382642 128452
rect 383534 128194 383562 128452
rect 384454 128194 384482 128452
rect 385374 128194 385402 128452
rect 386294 128194 386322 128452
rect 387122 128194 387150 128452
rect 388042 128194 388070 128452
rect 388962 128194 388990 128452
rect 389882 128194 389910 128452
rect 390802 128194 390830 128452
rect 391722 128194 391750 128452
rect 392642 128194 392670 128452
rect 393470 128194 393498 128452
rect 394390 128194 394418 128452
rect 395310 128194 395338 128452
rect 396230 128194 396258 128452
rect 397150 128194 397178 128452
rect 398070 128194 398098 128452
rect 398990 128194 399018 128452
rect 399818 128194 399846 128452
rect 400738 128194 400766 128452
rect 401658 128194 401686 128452
rect 402578 128194 402606 128452
rect 403498 128194 403526 128452
rect 404418 128194 404446 128452
rect 405338 128194 405366 128452
rect 406166 128194 406194 128452
rect 407086 128194 407114 128452
rect 379026 128166 379468 128194
rect 379854 128166 379928 128194
rect 380774 128166 380848 128194
rect 381694 128166 381768 128194
rect 382614 128166 382688 128194
rect 383534 128166 383608 128194
rect 384454 128166 384528 128194
rect 385374 128166 385448 128194
rect 386294 128166 386368 128194
rect 387122 128166 387196 128194
rect 388042 128166 388116 128194
rect 388962 128166 389128 128194
rect 389882 128166 389956 128194
rect 390802 128166 390876 128194
rect 391722 128166 391888 128194
rect 392642 128166 392716 128194
rect 393470 128166 393544 128194
rect 394390 128166 394648 128194
rect 395310 128166 395384 128194
rect 396230 128166 396304 128194
rect 397150 128166 397408 128194
rect 398070 128166 398144 128194
rect 398990 128166 399064 128194
rect 399818 128166 400168 128194
rect 400738 128166 400812 128194
rect 401658 128166 401732 128194
rect 402578 128166 402928 128194
rect 403498 128166 403572 128194
rect 404418 128166 404492 128194
rect 405338 128166 405688 128194
rect 406166 128166 406240 128194
rect 377220 126336 377272 126342
rect 377220 126278 377272 126284
rect 378060 3874 378088 128166
rect 379440 3942 379468 128166
rect 379900 126274 379928 128166
rect 379888 126268 379940 126274
rect 379888 126210 379940 126216
rect 378876 3936 378928 3942
rect 378876 3878 378928 3884
rect 379428 3936 379480 3942
rect 379428 3878 379480 3884
rect 377680 3868 377732 3874
rect 377680 3810 377732 3816
rect 378048 3868 378100 3874
rect 378048 3810 378100 3816
rect 376668 3324 376720 3330
rect 376668 3266 376720 3272
rect 376312 598 376524 626
rect 376312 490 376340 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 462 376340 490
rect 376496 480 376524 598
rect 377692 480 377720 3810
rect 378888 480 378916 3878
rect 380820 3738 380848 128166
rect 381740 125662 381768 128166
rect 382660 125662 382688 128166
rect 381728 125656 381780 125662
rect 381728 125598 381780 125604
rect 382188 125656 382240 125662
rect 382188 125598 382240 125604
rect 382648 125656 382700 125662
rect 382648 125598 382700 125604
rect 383476 125656 383528 125662
rect 383476 125598 383528 125604
rect 382200 4010 382228 125598
rect 383488 4894 383516 125598
rect 383476 4888 383528 4894
rect 383476 4830 383528 4836
rect 381176 4004 381228 4010
rect 381176 3946 381228 3952
rect 382188 4004 382240 4010
rect 382188 3946 382240 3952
rect 380808 3732 380860 3738
rect 380808 3674 380860 3680
rect 379980 3596 380032 3602
rect 379980 3538 380032 3544
rect 379992 480 380020 3538
rect 381188 480 381216 3946
rect 383580 3806 383608 128166
rect 384500 125662 384528 128166
rect 385420 125662 385448 128166
rect 384488 125656 384540 125662
rect 384488 125598 384540 125604
rect 384948 125656 385000 125662
rect 384948 125598 385000 125604
rect 385408 125656 385460 125662
rect 385408 125598 385460 125604
rect 386236 125656 386288 125662
rect 386236 125598 386288 125604
rect 382372 3800 382424 3806
rect 382372 3742 382424 3748
rect 383568 3800 383620 3806
rect 383568 3742 383620 3748
rect 382384 480 382412 3742
rect 383568 3664 383620 3670
rect 383568 3606 383620 3612
rect 383580 480 383608 3606
rect 384764 2916 384816 2922
rect 384764 2858 384816 2864
rect 384776 480 384804 2858
rect 384960 2854 384988 125598
rect 386248 11762 386276 125598
rect 386236 11756 386288 11762
rect 386236 11698 386288 11704
rect 386340 3602 386368 128166
rect 387168 125662 387196 128166
rect 388088 126410 388116 128166
rect 388076 126404 388128 126410
rect 388076 126346 388128 126352
rect 387156 125656 387208 125662
rect 387156 125598 387208 125604
rect 387708 125656 387760 125662
rect 387708 125598 387760 125604
rect 387720 3670 387748 125598
rect 387708 3664 387760 3670
rect 387708 3606 387760 3612
rect 386328 3596 386380 3602
rect 386328 3538 386380 3544
rect 389100 3534 389128 128166
rect 389824 126336 389876 126342
rect 389824 126278 389876 126284
rect 389836 5030 389864 126278
rect 389928 125662 389956 128166
rect 390848 125662 390876 128166
rect 389916 125656 389968 125662
rect 389916 125598 389968 125604
rect 390468 125656 390520 125662
rect 390468 125598 390520 125604
rect 390836 125656 390888 125662
rect 390836 125598 390888 125604
rect 389824 5024 389876 5030
rect 389824 4966 389876 4972
rect 387156 3528 387208 3534
rect 387156 3470 387208 3476
rect 389088 3528 389140 3534
rect 389088 3470 389140 3476
rect 385960 2984 386012 2990
rect 385960 2926 386012 2932
rect 384948 2848 385000 2854
rect 384948 2790 385000 2796
rect 385972 480 386000 2926
rect 387168 480 387196 3470
rect 389456 3120 389508 3126
rect 389456 3062 389508 3068
rect 388260 3052 388312 3058
rect 388260 2994 388312 3000
rect 388272 480 388300 2994
rect 389468 480 389496 3062
rect 390480 2922 390508 125598
rect 391756 4820 391808 4826
rect 391756 4762 391808 4768
rect 390652 3460 390704 3466
rect 390652 3402 390704 3408
rect 390468 2916 390520 2922
rect 390468 2858 390520 2864
rect 390664 480 390692 3402
rect 391768 2394 391796 4762
rect 391860 3466 391888 128166
rect 392688 125662 392716 128166
rect 393516 126342 393544 128166
rect 393504 126336 393556 126342
rect 393504 126278 393556 126284
rect 392584 125656 392636 125662
rect 392584 125598 392636 125604
rect 392676 125656 392728 125662
rect 392676 125598 392728 125604
rect 393228 125656 393280 125662
rect 393228 125598 393280 125604
rect 392596 5166 392624 125598
rect 392584 5160 392636 5166
rect 392584 5102 392636 5108
rect 391848 3460 391900 3466
rect 391848 3402 391900 3408
rect 393044 3188 393096 3194
rect 393044 3130 393096 3136
rect 391768 2366 391888 2394
rect 391860 480 391888 2366
rect 393056 480 393084 3130
rect 393240 3058 393268 125598
rect 394240 3392 394292 3398
rect 394240 3334 394292 3340
rect 393228 3052 393280 3058
rect 393228 2994 393280 3000
rect 394252 480 394280 3334
rect 394620 3194 394648 128166
rect 395356 125662 395384 128166
rect 396276 125662 396304 128166
rect 395344 125656 395396 125662
rect 395344 125598 395396 125604
rect 395988 125656 396040 125662
rect 395988 125598 396040 125604
rect 396264 125656 396316 125662
rect 396264 125598 396316 125604
rect 397276 125656 397328 125662
rect 397276 125598 397328 125604
rect 395344 7608 395396 7614
rect 395344 7550 395396 7556
rect 394608 3188 394660 3194
rect 394608 3130 394660 3136
rect 395356 480 395384 7550
rect 396000 2990 396028 125598
rect 397288 4826 397316 125598
rect 397276 4820 397328 4826
rect 397276 4762 397328 4768
rect 397380 3398 397408 128166
rect 398116 125662 398144 128166
rect 399036 126546 399064 128166
rect 399024 126540 399076 126546
rect 399024 126482 399076 126488
rect 398104 125656 398156 125662
rect 398104 125598 398156 125604
rect 398748 125656 398800 125662
rect 398748 125598 398800 125604
rect 397736 4072 397788 4078
rect 397736 4014 397788 4020
rect 397368 3392 397420 3398
rect 397368 3334 397420 3340
rect 396540 3256 396592 3262
rect 396540 3198 396592 3204
rect 395988 2984 396040 2990
rect 395988 2926 396040 2932
rect 396552 480 396580 3198
rect 397748 480 397776 4014
rect 398760 3126 398788 125598
rect 398932 4956 398984 4962
rect 398932 4898 398984 4904
rect 398748 3120 398800 3126
rect 398748 3062 398800 3068
rect 398944 480 398972 4898
rect 400140 4146 400168 128166
rect 400784 125662 400812 128166
rect 401704 126954 401732 128166
rect 401692 126948 401744 126954
rect 401692 126890 401744 126896
rect 400864 126268 400916 126274
rect 400864 126210 400916 126216
rect 400772 125656 400824 125662
rect 400772 125598 400824 125604
rect 400876 4962 400904 126210
rect 401508 125656 401560 125662
rect 401508 125598 401560 125604
rect 400864 4956 400916 4962
rect 400864 4898 400916 4904
rect 400036 4140 400088 4146
rect 400036 4082 400088 4088
rect 400128 4140 400180 4146
rect 400128 4082 400180 4088
rect 400048 2122 400076 4082
rect 401520 3330 401548 125598
rect 402520 5024 402572 5030
rect 402520 4966 402572 4972
rect 401324 3324 401376 3330
rect 401324 3266 401376 3272
rect 401508 3324 401560 3330
rect 401508 3266 401560 3272
rect 400048 2094 400168 2122
rect 400140 480 400168 2094
rect 401336 480 401364 3266
rect 402532 480 402560 4966
rect 402900 4078 402928 128166
rect 403544 125662 403572 128166
rect 403624 126948 403676 126954
rect 403624 126890 403676 126896
rect 403532 125656 403584 125662
rect 403532 125598 403584 125604
rect 403636 5098 403664 126890
rect 404464 126274 404492 128166
rect 404452 126268 404504 126274
rect 404452 126210 404504 126216
rect 404268 125656 404320 125662
rect 404268 125598 404320 125604
rect 403624 5092 403676 5098
rect 403624 5034 403676 5040
rect 402888 4072 402940 4078
rect 402888 4014 402940 4020
rect 403624 3868 403676 3874
rect 403624 3810 403676 3816
rect 403636 480 403664 3810
rect 404280 3262 404308 125598
rect 405660 3942 405688 128166
rect 406212 125662 406240 128166
rect 406948 128166 407114 128194
rect 408006 128194 408034 128452
rect 408926 128194 408954 128452
rect 409846 128194 409874 128452
rect 408006 128166 408448 128194
rect 408926 128166 409000 128194
rect 406200 125656 406252 125662
rect 406200 125598 406252 125604
rect 406948 5030 406976 128166
rect 407764 126404 407816 126410
rect 407764 126346 407816 126352
rect 407028 125656 407080 125662
rect 407028 125598 407080 125604
rect 406936 5024 406988 5030
rect 406936 4966 406988 4972
rect 406016 4956 406068 4962
rect 406016 4898 406068 4904
rect 404820 3936 404872 3942
rect 404820 3878 404872 3884
rect 405648 3936 405700 3942
rect 405648 3878 405700 3884
rect 404268 3256 404320 3262
rect 404268 3198 404320 3204
rect 404832 480 404860 3878
rect 406028 480 406056 4898
rect 407040 4010 407068 125598
rect 407776 5234 407804 126346
rect 408420 6914 408448 128166
rect 408972 125662 409000 128166
rect 409800 128166 409874 128194
rect 410766 128194 410794 128452
rect 411686 128194 411714 128452
rect 412514 128194 412542 128452
rect 410766 128166 411208 128194
rect 411686 128166 411760 128194
rect 409800 126478 409828 128166
rect 409788 126472 409840 126478
rect 409788 126414 409840 126420
rect 408960 125656 409012 125662
rect 408960 125598 409012 125604
rect 409788 125656 409840 125662
rect 409788 125598 409840 125604
rect 408328 6886 408448 6914
rect 407764 5228 407816 5234
rect 407764 5170 407816 5176
rect 407028 4004 407080 4010
rect 407028 3946 407080 3952
rect 408328 3874 408356 6886
rect 409604 4888 409656 4894
rect 409604 4830 409656 4836
rect 408224 3868 408276 3874
rect 408224 3810 408276 3816
rect 408316 3868 408368 3874
rect 408316 3810 408368 3816
rect 407212 3732 407264 3738
rect 407212 3674 407264 3680
rect 407224 480 407252 3674
rect 408236 1986 408264 3810
rect 408236 1958 408448 1986
rect 408420 480 408448 1958
rect 409616 480 409644 4830
rect 409800 3262 409828 125598
rect 411180 3806 411208 128166
rect 411732 125662 411760 128166
rect 412468 128166 412542 128194
rect 413434 128194 413462 128452
rect 414354 128194 414382 128452
rect 415274 128194 415302 128452
rect 416194 128194 416222 128452
rect 417114 128194 417142 128452
rect 418034 128194 418062 128452
rect 413434 128166 413508 128194
rect 414354 128166 414428 128194
rect 415274 128166 415348 128194
rect 416194 128166 416268 128194
rect 417114 128166 417188 128194
rect 411720 125656 411772 125662
rect 411720 125598 411772 125604
rect 412468 4962 412496 128166
rect 413480 125662 413508 128166
rect 414400 125662 414428 128166
rect 415320 126682 415348 128166
rect 415308 126676 415360 126682
rect 415308 126618 415360 126624
rect 416240 125662 416268 128166
rect 417160 125662 417188 128166
rect 417988 128166 418062 128194
rect 418862 128194 418890 128452
rect 419782 128194 419810 128452
rect 420702 128194 420730 128452
rect 421622 128194 421650 128452
rect 422542 128194 422570 128452
rect 423462 128194 423490 128452
rect 424382 128194 424410 128452
rect 425210 128194 425238 128452
rect 426130 128194 426158 128452
rect 427050 128194 427078 128452
rect 427970 128194 427998 128452
rect 428890 128194 428918 128452
rect 429810 128194 429838 128452
rect 430730 128194 430758 128452
rect 431650 128194 431678 128452
rect 432478 128194 432506 128452
rect 433398 128194 433426 128452
rect 434318 128194 434346 128452
rect 435238 128194 435266 128452
rect 436158 128194 436186 128452
rect 437078 128194 437106 128452
rect 437998 128194 438026 128452
rect 438826 128194 438854 128452
rect 418862 128166 418936 128194
rect 419782 128166 419856 128194
rect 420702 128166 420776 128194
rect 421622 128166 421696 128194
rect 422542 128166 422616 128194
rect 423462 128166 423536 128194
rect 424382 128166 424456 128194
rect 425210 128166 425284 128194
rect 426130 128166 426296 128194
rect 427050 128166 427124 128194
rect 427970 128166 428044 128194
rect 428890 128166 428964 128194
rect 429810 128166 429884 128194
rect 430730 128166 430804 128194
rect 431650 128166 431816 128194
rect 432478 128166 432552 128194
rect 433398 128166 433472 128194
rect 434318 128166 434392 128194
rect 435238 128166 435312 128194
rect 436158 128166 436232 128194
rect 437078 128166 437152 128194
rect 437998 128166 438072 128194
rect 412548 125656 412600 125662
rect 412548 125598 412600 125604
rect 413468 125656 413520 125662
rect 413468 125598 413520 125604
rect 413928 125656 413980 125662
rect 413928 125598 413980 125604
rect 414388 125656 414440 125662
rect 414388 125598 414440 125604
rect 415308 125656 415360 125662
rect 415308 125598 415360 125604
rect 416228 125656 416280 125662
rect 416228 125598 416280 125604
rect 416688 125656 416740 125662
rect 416688 125598 416740 125604
rect 417148 125656 417200 125662
rect 417148 125598 417200 125604
rect 412456 4956 412508 4962
rect 412456 4898 412508 4904
rect 410800 3800 410852 3806
rect 410800 3742 410852 3748
rect 411168 3800 411220 3806
rect 412560 3777 412588 125598
rect 412640 11756 412692 11762
rect 412640 11698 412692 11704
rect 411168 3742 411220 3748
rect 412546 3768 412602 3777
rect 409788 3256 409840 3262
rect 409788 3198 409840 3204
rect 410812 480 410840 3742
rect 412546 3703 412602 3712
rect 411904 2848 411956 2854
rect 411904 2790 411956 2796
rect 411916 480 411944 2790
rect 412652 490 412680 11698
rect 413940 3738 413968 125598
rect 413928 3732 413980 3738
rect 413928 3674 413980 3680
rect 415320 3602 415348 125598
rect 416700 6914 416728 125598
rect 416608 6886 416728 6914
rect 416608 3670 416636 6886
rect 416688 5228 416740 5234
rect 416688 5170 416740 5176
rect 415492 3664 415544 3670
rect 415492 3606 415544 3612
rect 416596 3664 416648 3670
rect 416596 3606 416648 3612
rect 414296 3596 414348 3602
rect 414296 3538 414348 3544
rect 415308 3596 415360 3602
rect 415308 3538 415360 3544
rect 412928 598 413140 626
rect 412928 490 412956 598
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 462 412956 490
rect 413112 480 413140 598
rect 414308 480 414336 3538
rect 415504 480 415532 3606
rect 416700 480 416728 5170
rect 417988 4894 418016 128166
rect 418804 126540 418856 126546
rect 418804 126482 418856 126488
rect 418068 125656 418120 125662
rect 418068 125598 418120 125604
rect 417976 4888 418028 4894
rect 417976 4830 418028 4836
rect 418080 3738 418108 125598
rect 418816 5234 418844 126482
rect 418908 125662 418936 128166
rect 419828 126546 419856 128166
rect 420748 126614 420776 128166
rect 420736 126608 420788 126614
rect 420736 126550 420788 126556
rect 419816 126540 419868 126546
rect 419816 126482 419868 126488
rect 421564 126336 421616 126342
rect 421564 126278 421616 126284
rect 418896 125656 418948 125662
rect 418896 125598 418948 125604
rect 419448 125656 419500 125662
rect 419448 125598 419500 125604
rect 418804 5228 418856 5234
rect 418804 5170 418856 5176
rect 418068 3732 418120 3738
rect 418068 3674 418120 3680
rect 419460 3670 419488 125598
rect 420184 5160 420236 5166
rect 420184 5102 420236 5108
rect 419448 3664 419500 3670
rect 419448 3606 419500 3612
rect 417884 3528 417936 3534
rect 417884 3470 417936 3476
rect 417896 480 417924 3470
rect 418988 2916 419040 2922
rect 418988 2858 419040 2864
rect 419000 480 419028 2858
rect 420196 480 420224 5102
rect 421576 4486 421604 126278
rect 421668 125662 421696 128166
rect 422588 125662 422616 128166
rect 423508 126342 423536 128166
rect 423496 126336 423548 126342
rect 423496 126278 423548 126284
rect 424428 125662 424456 128166
rect 425256 125662 425284 128166
rect 421656 125656 421708 125662
rect 421656 125598 421708 125604
rect 422208 125656 422260 125662
rect 422208 125598 422260 125604
rect 422576 125656 422628 125662
rect 422576 125598 422628 125604
rect 423588 125656 423640 125662
rect 423588 125598 423640 125604
rect 424416 125656 424468 125662
rect 424416 125598 424468 125604
rect 424968 125656 425020 125662
rect 424968 125598 425020 125604
rect 425244 125656 425296 125662
rect 425244 125598 425296 125604
rect 421564 4480 421616 4486
rect 421564 4422 421616 4428
rect 421380 3596 421432 3602
rect 421380 3538 421432 3544
rect 421392 480 421420 3538
rect 422220 3534 422248 125598
rect 422208 3528 422260 3534
rect 422208 3470 422260 3476
rect 423600 3194 423628 125598
rect 424980 6914 425008 125598
rect 426268 10334 426296 128166
rect 427096 125662 427124 128166
rect 428016 125662 428044 128166
rect 428936 126410 428964 128166
rect 429752 126472 429804 126478
rect 429752 126414 429804 126420
rect 428924 126404 428976 126410
rect 428924 126346 428976 126352
rect 426348 125656 426400 125662
rect 426348 125598 426400 125604
rect 427084 125656 427136 125662
rect 427084 125598 427136 125604
rect 427728 125656 427780 125662
rect 427728 125598 427780 125604
rect 428004 125656 428056 125662
rect 428004 125598 428056 125604
rect 429108 125656 429160 125662
rect 429108 125598 429160 125604
rect 426256 10328 426308 10334
rect 426256 10270 426308 10276
rect 424888 6886 425008 6914
rect 423772 4480 423824 4486
rect 423772 4422 423824 4428
rect 422576 3188 422628 3194
rect 422576 3130 422628 3136
rect 423588 3188 423640 3194
rect 423588 3130 423640 3136
rect 422588 480 422616 3130
rect 423784 480 423812 4422
rect 424888 3194 424916 6886
rect 426360 3641 426388 125598
rect 427268 4820 427320 4826
rect 427268 4762 427320 4768
rect 426346 3632 426402 3641
rect 426346 3567 426402 3576
rect 424968 3460 425020 3466
rect 424968 3402 425020 3408
rect 424876 3188 424928 3194
rect 424876 3130 424928 3136
rect 424980 480 425008 3402
rect 426164 2984 426216 2990
rect 426164 2926 426216 2932
rect 426176 480 426204 2926
rect 427280 480 427308 4762
rect 427740 3194 427768 125598
rect 428464 3392 428516 3398
rect 428464 3334 428516 3340
rect 427728 3188 427780 3194
rect 427728 3130 427780 3136
rect 428476 480 428504 3334
rect 429120 3058 429148 125598
rect 429764 122834 429792 126414
rect 429856 125662 429884 128166
rect 430776 125662 430804 128166
rect 429844 125656 429896 125662
rect 429844 125598 429896 125604
rect 430488 125656 430540 125662
rect 430488 125598 430540 125604
rect 430764 125656 430816 125662
rect 430764 125598 430816 125604
rect 429764 122806 429884 122834
rect 429856 5166 429884 122806
rect 429844 5160 429896 5166
rect 429844 5102 429896 5108
rect 430500 3126 430528 125598
rect 430856 5228 430908 5234
rect 430856 5170 430908 5176
rect 429660 3120 429712 3126
rect 429660 3062 429712 3068
rect 430488 3120 430540 3126
rect 430488 3062 430540 3068
rect 429108 3052 429160 3058
rect 429108 2994 429160 3000
rect 429672 480 429700 3062
rect 430868 480 430896 5170
rect 431788 4826 431816 128166
rect 432524 125662 432552 128166
rect 432604 126608 432656 126614
rect 432604 126550 432656 126556
rect 431868 125656 431920 125662
rect 431868 125598 431920 125604
rect 432512 125656 432564 125662
rect 432512 125598 432564 125604
rect 431776 4820 431828 4826
rect 431776 4762 431828 4768
rect 431880 3505 431908 125598
rect 432616 7614 432644 126550
rect 433444 125662 433472 128166
rect 434364 126478 434392 128166
rect 434352 126472 434404 126478
rect 434352 126414 434404 126420
rect 435284 125662 435312 128166
rect 436204 125662 436232 128166
rect 437124 126614 437152 128166
rect 437112 126608 437164 126614
rect 437112 126550 437164 126556
rect 436744 126268 436796 126274
rect 436744 126210 436796 126216
rect 433248 125656 433300 125662
rect 433248 125598 433300 125604
rect 433432 125656 433484 125662
rect 433432 125598 433484 125604
rect 434628 125656 434680 125662
rect 434628 125598 434680 125604
rect 435272 125656 435324 125662
rect 435272 125598 435324 125604
rect 436008 125656 436060 125662
rect 436008 125598 436060 125604
rect 436192 125656 436244 125662
rect 436192 125598 436244 125604
rect 432604 7608 432656 7614
rect 432604 7550 432656 7556
rect 433260 6914 433288 125598
rect 433168 6886 433288 6914
rect 432052 4140 432104 4146
rect 432052 4082 432104 4088
rect 431866 3496 431922 3505
rect 431866 3431 431922 3440
rect 432064 480 432092 4082
rect 433168 4010 433196 6886
rect 434444 5092 434496 5098
rect 434444 5034 434496 5040
rect 433156 4004 433208 4010
rect 433156 3946 433208 3952
rect 433248 3324 433300 3330
rect 433248 3266 433300 3272
rect 433260 480 433288 3266
rect 434456 480 434484 5034
rect 434640 3330 434668 125598
rect 436020 4078 436048 125598
rect 436756 4214 436784 126210
rect 438044 125662 438072 128166
rect 438780 128166 438854 128194
rect 439746 128194 439774 128452
rect 440666 128194 440694 128452
rect 441586 128194 441614 128452
rect 439746 128166 440188 128194
rect 440666 128166 440740 128194
rect 437388 125656 437440 125662
rect 437388 125598 437440 125604
rect 438032 125656 438084 125662
rect 438032 125598 438084 125604
rect 436744 4208 436796 4214
rect 436744 4150 436796 4156
rect 437400 4146 437428 125598
rect 437940 4208 437992 4214
rect 437940 4150 437992 4156
rect 437388 4140 437440 4146
rect 437388 4082 437440 4088
rect 435548 4072 435600 4078
rect 435548 4014 435600 4020
rect 436008 4072 436060 4078
rect 436008 4014 436060 4020
rect 434628 3324 434680 3330
rect 434628 3266 434680 3272
rect 435560 480 435588 4014
rect 436468 3256 436520 3262
rect 436468 3198 436520 3204
rect 436480 1714 436508 3198
rect 436480 1686 436784 1714
rect 436756 480 436784 1686
rect 437952 480 437980 4150
rect 438780 3369 438808 128166
rect 439504 125656 439556 125662
rect 439504 125598 439556 125604
rect 439516 15910 439544 125598
rect 439504 15904 439556 15910
rect 439504 15846 439556 15852
rect 440160 5370 440188 128166
rect 440712 126818 440740 128166
rect 441540 128166 441614 128194
rect 442506 128194 442534 128452
rect 443426 128194 443454 128452
rect 444346 128194 444374 128452
rect 442506 128166 442580 128194
rect 443426 128166 443500 128194
rect 440700 126812 440752 126818
rect 440700 126754 440752 126760
rect 440148 5364 440200 5370
rect 440148 5306 440200 5312
rect 441436 5024 441488 5030
rect 441436 4966 441488 4972
rect 440332 4004 440384 4010
rect 440332 3946 440384 3952
rect 439136 3936 439188 3942
rect 439136 3878 439188 3884
rect 438766 3360 438822 3369
rect 438766 3295 438822 3304
rect 439148 480 439176 3878
rect 440344 480 440372 3946
rect 441448 2530 441476 4966
rect 441540 4010 441568 128166
rect 442264 126676 442316 126682
rect 442264 126618 442316 126624
rect 442276 5030 442304 126618
rect 442552 126274 442580 128166
rect 442540 126268 442592 126274
rect 442540 126210 442592 126216
rect 443472 125662 443500 128166
rect 444300 128166 444374 128194
rect 445174 128194 445202 128452
rect 446094 128194 446122 128452
rect 447014 128194 447042 128452
rect 447934 128194 447962 128452
rect 448854 128194 448882 128452
rect 449774 128194 449802 128452
rect 450694 128194 450722 128452
rect 451522 128194 451550 128452
rect 452442 128194 452470 128452
rect 453362 128194 453390 128452
rect 454282 128194 454310 128452
rect 455202 128194 455230 128452
rect 456122 128194 456150 128452
rect 457042 128194 457070 128452
rect 457870 128194 457898 128452
rect 458790 128194 458818 128452
rect 459710 128194 459738 128452
rect 460630 128194 460658 128452
rect 461550 128194 461578 128452
rect 462470 128194 462498 128452
rect 463390 128194 463418 128452
rect 464218 128194 464246 128452
rect 465138 128194 465166 128452
rect 466058 128194 466086 128452
rect 466978 128194 467006 128452
rect 467898 128194 467926 128452
rect 468818 128194 468846 128452
rect 469738 128194 469766 128452
rect 470566 128194 470594 128452
rect 445174 128166 445248 128194
rect 446094 128166 446168 128194
rect 447014 128166 447088 128194
rect 447934 128166 448008 128194
rect 448854 128166 448928 128194
rect 449774 128166 449848 128194
rect 450694 128166 450768 128194
rect 451522 128166 451596 128194
rect 452442 128166 452608 128194
rect 453362 128166 453436 128194
rect 454282 128166 454356 128194
rect 455202 128166 455368 128194
rect 456122 128166 456196 128194
rect 457042 128166 457116 128194
rect 457870 128166 458128 128194
rect 458790 128166 458864 128194
rect 459710 128166 459784 128194
rect 460630 128166 460888 128194
rect 461550 128166 461624 128194
rect 462470 128166 462544 128194
rect 463390 128166 463648 128194
rect 464218 128166 464292 128194
rect 465138 128166 465212 128194
rect 466058 128166 466132 128194
rect 466978 128166 467052 128194
rect 467898 128166 467972 128194
rect 468818 128166 469168 128194
rect 469738 128166 469812 128194
rect 443460 125656 443512 125662
rect 443460 125598 443512 125604
rect 444196 125656 444248 125662
rect 444196 125598 444248 125604
rect 444208 9042 444236 125598
rect 444196 9036 444248 9042
rect 444196 8978 444248 8984
rect 442264 5024 442316 5030
rect 442264 4966 442316 4972
rect 441528 4004 441580 4010
rect 441528 3946 441580 3952
rect 444300 3942 444328 128166
rect 445220 125730 445248 128166
rect 445208 125724 445260 125730
rect 445208 125666 445260 125672
rect 446140 125662 446168 128166
rect 446128 125656 446180 125662
rect 446128 125598 446180 125604
rect 446956 125656 447008 125662
rect 446956 125598 447008 125604
rect 446968 5302 446996 125598
rect 446956 5296 447008 5302
rect 446956 5238 447008 5244
rect 445024 5160 445076 5166
rect 445024 5102 445076 5108
rect 444288 3936 444340 3942
rect 444288 3878 444340 3884
rect 442632 3868 442684 3874
rect 442632 3810 442684 3816
rect 441448 2502 441568 2530
rect 441540 480 441568 2502
rect 442644 480 442672 3810
rect 443828 2848 443880 2854
rect 443828 2790 443880 2796
rect 443840 480 443868 2790
rect 445036 480 445064 5102
rect 447060 3874 447088 128166
rect 447784 125724 447836 125730
rect 447784 125666 447836 125672
rect 447796 89010 447824 125666
rect 447980 125662 448008 128166
rect 448900 126750 448928 128166
rect 448888 126744 448940 126750
rect 448888 126686 448940 126692
rect 447968 125656 448020 125662
rect 447968 125598 448020 125604
rect 448428 125656 448480 125662
rect 448428 125598 448480 125604
rect 447784 89004 447836 89010
rect 447784 88946 447836 88952
rect 448440 5234 448468 125598
rect 449820 6914 449848 128166
rect 450544 126812 450596 126818
rect 450544 126754 450596 126760
rect 450556 11762 450584 126754
rect 450740 125662 450768 128166
rect 451568 126002 451596 128166
rect 451556 125996 451608 126002
rect 451556 125938 451608 125944
rect 450728 125656 450780 125662
rect 450728 125598 450780 125604
rect 451188 125656 451240 125662
rect 451188 125598 451240 125604
rect 450544 11756 450596 11762
rect 450544 11698 450596 11704
rect 449728 6886 449848 6914
rect 448428 5228 448480 5234
rect 448428 5170 448480 5176
rect 448612 4956 448664 4962
rect 448612 4898 448664 4904
rect 447048 3868 447100 3874
rect 447048 3810 447100 3816
rect 446220 3800 446272 3806
rect 446220 3742 446272 3748
rect 447414 3768 447470 3777
rect 446232 480 446260 3742
rect 447414 3703 447470 3712
rect 447428 480 447456 3703
rect 448624 480 448652 4898
rect 449728 3806 449756 6886
rect 451200 5098 451228 125598
rect 451188 5092 451240 5098
rect 451188 5034 451240 5040
rect 452108 5024 452160 5030
rect 452108 4966 452160 4972
rect 449716 3800 449768 3806
rect 449716 3742 449768 3748
rect 449808 3732 449860 3738
rect 449808 3674 449860 3680
rect 449820 480 449848 3674
rect 450912 2916 450964 2922
rect 450912 2858 450964 2864
rect 450924 480 450952 2858
rect 452120 480 452148 4966
rect 452580 3738 452608 128166
rect 453408 125662 453436 128166
rect 454328 125662 454356 128166
rect 453396 125656 453448 125662
rect 453396 125598 453448 125604
rect 453948 125656 454000 125662
rect 453948 125598 454000 125604
rect 454316 125656 454368 125662
rect 454316 125598 454368 125604
rect 455236 125656 455288 125662
rect 455236 125598 455288 125604
rect 453960 5166 453988 125598
rect 455248 90370 455276 125598
rect 455236 90364 455288 90370
rect 455236 90306 455288 90312
rect 453948 5160 454000 5166
rect 453948 5102 454000 5108
rect 452568 3732 452620 3738
rect 452568 3674 452620 3680
rect 454500 3664 454552 3670
rect 454500 3606 454552 3612
rect 453304 3596 453356 3602
rect 453304 3538 453356 3544
rect 453316 480 453344 3538
rect 454512 480 454540 3606
rect 455340 3602 455368 128166
rect 456168 126206 456196 128166
rect 457088 126682 457116 128166
rect 457076 126676 457128 126682
rect 457076 126618 457128 126624
rect 456892 126540 456944 126546
rect 456892 126482 456944 126488
rect 456156 126200 456208 126206
rect 456156 126142 456208 126148
rect 456904 16574 456932 126482
rect 456904 16546 458036 16574
rect 455696 4888 455748 4894
rect 455696 4830 455748 4836
rect 455328 3596 455380 3602
rect 455328 3538 455380 3544
rect 455708 480 455736 4830
rect 456892 3528 456944 3534
rect 456892 3470 456944 3476
rect 458008 3482 458036 16546
rect 458100 3670 458128 128166
rect 458836 125662 458864 128166
rect 459756 126546 459784 128166
rect 459744 126540 459796 126546
rect 459744 126482 459796 126488
rect 458824 125656 458876 125662
rect 458824 125598 458876 125604
rect 459468 125656 459520 125662
rect 459468 125598 459520 125604
rect 459480 26926 459508 125598
rect 459468 26920 459520 26926
rect 459468 26862 459520 26868
rect 459192 7608 459244 7614
rect 459192 7550 459244 7556
rect 458088 3664 458140 3670
rect 458088 3606 458140 3612
rect 456904 480 456932 3470
rect 458008 3454 458128 3482
rect 458100 480 458128 3454
rect 459204 480 459232 7550
rect 460860 3534 460888 128166
rect 461492 126336 461544 126342
rect 461492 126278 461544 126284
rect 461504 122834 461532 126278
rect 461596 125662 461624 128166
rect 462516 126070 462544 128166
rect 462504 126064 462556 126070
rect 462504 126006 462556 126012
rect 461584 125656 461636 125662
rect 461584 125598 461636 125604
rect 462228 125656 462280 125662
rect 462228 125598 462280 125604
rect 461504 122806 461624 122834
rect 461596 4214 461624 122806
rect 462240 4894 462268 125598
rect 462228 4888 462280 4894
rect 462228 4830 462280 4836
rect 461584 4208 461636 4214
rect 461584 4150 461636 4156
rect 462780 4208 462832 4214
rect 462780 4150 462832 4156
rect 460848 3528 460900 3534
rect 460848 3470 460900 3476
rect 460388 3460 460440 3466
rect 460388 3402 460440 3408
rect 460400 480 460428 3402
rect 461584 2984 461636 2990
rect 461584 2926 461636 2932
rect 461596 480 461624 2926
rect 462792 480 462820 4150
rect 463620 3466 463648 128166
rect 464264 125662 464292 128166
rect 464344 126676 464396 126682
rect 464344 126618 464396 126624
rect 464252 125656 464304 125662
rect 464252 125598 464304 125604
rect 464356 7682 464384 126618
rect 465184 125662 465212 128166
rect 466104 126818 466132 128166
rect 466092 126812 466144 126818
rect 466092 126754 466144 126760
rect 467024 125662 467052 128166
rect 467104 126404 467156 126410
rect 467104 126346 467156 126352
rect 464988 125656 465040 125662
rect 464988 125598 465040 125604
rect 465172 125656 465224 125662
rect 465172 125598 465224 125604
rect 466368 125656 466420 125662
rect 466368 125598 466420 125604
rect 467012 125656 467064 125662
rect 467012 125598 467064 125604
rect 464344 7676 464396 7682
rect 464344 7618 464396 7624
rect 465000 4962 465028 125598
rect 465816 10328 465868 10334
rect 465816 10270 465868 10276
rect 464988 4956 465040 4962
rect 464988 4898 465040 4904
rect 465170 3632 465226 3641
rect 465170 3567 465226 3576
rect 463608 3460 463660 3466
rect 463608 3402 463660 3408
rect 463976 3188 464028 3194
rect 463976 3130 464028 3136
rect 463988 480 464016 3130
rect 465184 480 465212 3567
rect 465828 490 465856 10270
rect 466380 6254 466408 125598
rect 466368 6248 466420 6254
rect 466368 6190 466420 6196
rect 467116 4214 467144 126346
rect 467944 125662 467972 128166
rect 467748 125656 467800 125662
rect 467748 125598 467800 125604
rect 467932 125656 467984 125662
rect 467932 125598 467984 125604
rect 469036 125656 469088 125662
rect 469036 125598 469088 125604
rect 467760 8974 467788 125598
rect 469048 10334 469076 125598
rect 469036 10328 469088 10334
rect 469036 10270 469088 10276
rect 467748 8968 467800 8974
rect 467748 8910 467800 8916
rect 467104 4208 467156 4214
rect 467104 4150 467156 4156
rect 468668 3120 468720 3126
rect 468668 3062 468720 3068
rect 467472 3052 467524 3058
rect 467472 2994 467524 3000
rect 466104 598 466316 626
rect 466104 490 466132 598
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 462 466132 490
rect 466288 480 466316 598
rect 467484 480 467512 2994
rect 468680 480 468708 3062
rect 469140 2854 469168 128166
rect 469784 126886 469812 128166
rect 470520 128166 470594 128194
rect 471486 128194 471514 128452
rect 472406 128194 472434 128452
rect 473326 128194 473354 128452
rect 471486 128166 471560 128194
rect 472406 128166 472480 128194
rect 469772 126880 469824 126886
rect 469772 126822 469824 126828
rect 470520 126342 470548 128166
rect 471532 126682 471560 128166
rect 472452 126954 472480 128166
rect 473280 128166 473354 128194
rect 474246 128194 474274 128452
rect 475166 128194 475194 128452
rect 476086 128194 476114 128452
rect 474246 128166 474688 128194
rect 475166 128166 475240 128194
rect 472440 126948 472492 126954
rect 472440 126890 472492 126896
rect 471520 126676 471572 126682
rect 471520 126618 471572 126624
rect 471336 126608 471388 126614
rect 471336 126550 471388 126556
rect 471244 126540 471296 126546
rect 471244 126482 471296 126488
rect 470508 126336 470560 126342
rect 470508 126278 470560 126284
rect 471256 5438 471284 126482
rect 471244 5432 471296 5438
rect 471244 5374 471296 5380
rect 471348 4690 471376 126550
rect 472624 126132 472676 126138
rect 472624 126074 472676 126080
rect 471336 4684 471388 4690
rect 471336 4626 471388 4632
rect 472636 4214 472664 126074
rect 473280 6186 473308 128166
rect 473268 6180 473320 6186
rect 473268 6122 473320 6128
rect 473452 4820 473504 4826
rect 473452 4762 473504 4768
rect 469864 4208 469916 4214
rect 469864 4150 469916 4156
rect 472624 4208 472676 4214
rect 472624 4150 472676 4156
rect 469128 2848 469180 2854
rect 469128 2790 469180 2796
rect 469876 480 469904 4150
rect 472254 3496 472310 3505
rect 472254 3431 472310 3440
rect 471060 3324 471112 3330
rect 471060 3266 471112 3272
rect 471072 480 471100 3266
rect 472268 480 472296 3431
rect 473464 480 473492 4762
rect 474556 3392 474608 3398
rect 474556 3334 474608 3340
rect 474568 480 474596 3334
rect 474660 2922 474688 128166
rect 475212 125322 475240 128166
rect 475948 128166 476114 128194
rect 477006 128194 477034 128452
rect 477834 128194 477862 128452
rect 478754 128194 478782 128452
rect 479674 128194 479702 128452
rect 480594 128194 480622 128452
rect 481514 128194 481542 128452
rect 482434 128194 482462 128452
rect 483354 128194 483382 128452
rect 484182 128194 484210 128452
rect 485102 128194 485130 128452
rect 486022 128194 486050 128452
rect 486942 128194 486970 128452
rect 487862 128194 487890 128452
rect 488782 128194 488810 128452
rect 489702 128194 489730 128452
rect 490530 128194 490558 128452
rect 491450 128194 491478 128452
rect 492370 128194 492398 128452
rect 493290 128194 493318 128452
rect 494210 128194 494238 128452
rect 495130 128194 495158 128452
rect 496050 128194 496078 128452
rect 496878 128194 496906 128452
rect 497798 128194 497826 128452
rect 498718 128194 498746 128452
rect 499638 128194 499666 128452
rect 500558 128194 500586 128452
rect 501478 128194 501506 128452
rect 502398 128194 502426 128452
rect 503226 128194 503254 128452
rect 504146 128194 504174 128452
rect 505066 128194 505094 128452
rect 477006 128166 477080 128194
rect 477834 128166 477908 128194
rect 478754 128166 478828 128194
rect 479674 128166 479748 128194
rect 480594 128166 480668 128194
rect 481514 128166 481588 128194
rect 482434 128166 482508 128194
rect 483354 128166 483428 128194
rect 484182 128166 484256 128194
rect 485102 128166 485176 128194
rect 486022 128166 486096 128194
rect 486942 128166 487016 128194
rect 487862 128166 487936 128194
rect 488782 128166 488856 128194
rect 489702 128166 489776 128194
rect 490530 128166 490604 128194
rect 491450 128166 491524 128194
rect 492370 128166 492444 128194
rect 493290 128166 493364 128194
rect 494210 128166 494284 128194
rect 495130 128166 495296 128194
rect 496050 128166 496124 128194
rect 496878 128166 496952 128194
rect 497798 128166 498056 128194
rect 498718 128166 498792 128194
rect 499638 128166 499712 128194
rect 500558 128166 500816 128194
rect 501478 128166 501552 128194
rect 502398 128166 502472 128194
rect 503226 128166 503576 128194
rect 504146 128166 504220 128194
rect 475384 126336 475436 126342
rect 475384 126278 475436 126284
rect 475200 125316 475252 125322
rect 475200 125258 475252 125264
rect 475396 5030 475424 126278
rect 475384 5024 475436 5030
rect 475384 4966 475436 4972
rect 475948 4826 475976 128166
rect 477052 126750 477080 128166
rect 477040 126744 477092 126750
rect 477040 126686 477092 126692
rect 476764 126200 476816 126206
rect 476764 126142 476816 126148
rect 476776 5506 476804 126142
rect 477880 126138 477908 128166
rect 478800 126546 478828 128166
rect 479524 126608 479576 126614
rect 479524 126550 479576 126556
rect 478788 126540 478840 126546
rect 478788 126482 478840 126488
rect 477868 126132 477920 126138
rect 477868 126074 477920 126080
rect 476764 5500 476816 5506
rect 476764 5442 476816 5448
rect 475936 4820 475988 4826
rect 475936 4762 475988 4768
rect 479536 4758 479564 126550
rect 479720 125662 479748 128166
rect 480640 125662 480668 128166
rect 479708 125656 479760 125662
rect 479708 125598 479760 125604
rect 480168 125656 480220 125662
rect 480168 125598 480220 125604
rect 480628 125656 480680 125662
rect 480628 125598 480680 125604
rect 481560 125610 481588 128166
rect 482480 126342 482508 128166
rect 482468 126336 482520 126342
rect 482468 126278 482520 126284
rect 482284 126268 482336 126274
rect 482284 126210 482336 126216
rect 479524 4752 479576 4758
rect 479524 4694 479576 4700
rect 476948 4208 477000 4214
rect 476948 4150 477000 4156
rect 475752 3256 475804 3262
rect 475752 3198 475804 3204
rect 474648 2916 474700 2922
rect 474648 2858 474700 2864
rect 475764 480 475792 3198
rect 476960 480 476988 4150
rect 479340 4140 479392 4146
rect 479340 4082 479392 4088
rect 478144 4072 478196 4078
rect 478144 4014 478196 4020
rect 478156 480 478184 4014
rect 479352 480 479380 4082
rect 480180 2990 480208 125598
rect 481560 125582 481680 125610
rect 481652 125254 481680 125582
rect 481640 125248 481692 125254
rect 481640 125190 481692 125196
rect 481732 15904 481784 15910
rect 481732 15846 481784 15852
rect 480536 4684 480588 4690
rect 480536 4626 480588 4632
rect 480168 2984 480220 2990
rect 480168 2926 480220 2932
rect 480548 480 480576 4626
rect 481744 480 481772 15846
rect 482296 4214 482324 126210
rect 483400 126206 483428 128166
rect 484228 126478 484256 128166
rect 484216 126472 484268 126478
rect 484216 126414 484268 126420
rect 483388 126200 483440 126206
rect 483388 126142 483440 126148
rect 483664 125996 483716 126002
rect 483664 125938 483716 125944
rect 483676 5370 483704 125938
rect 485148 125662 485176 128166
rect 486068 126002 486096 128166
rect 486988 126410 487016 128166
rect 486976 126404 487028 126410
rect 486976 126346 487028 126352
rect 486056 125996 486108 126002
rect 486056 125938 486108 125944
rect 487908 125662 487936 128166
rect 485136 125656 485188 125662
rect 485136 125598 485188 125604
rect 485688 125656 485740 125662
rect 485688 125598 485740 125604
rect 487896 125656 487948 125662
rect 487896 125598 487948 125604
rect 488448 125656 488500 125662
rect 488448 125598 488500 125604
rect 484768 11756 484820 11762
rect 484768 11698 484820 11704
rect 483020 5364 483072 5370
rect 483020 5306 483072 5312
rect 483664 5364 483716 5370
rect 483664 5306 483716 5312
rect 483032 4282 483060 5306
rect 483020 4276 483072 4282
rect 483020 4218 483072 4224
rect 484032 4276 484084 4282
rect 484032 4218 484084 4224
rect 482284 4208 482336 4214
rect 482284 4150 482336 4156
rect 482834 3360 482890 3369
rect 482834 3295 482890 3304
rect 482848 480 482876 3295
rect 484044 480 484072 4218
rect 484780 490 484808 11698
rect 485700 3058 485728 125598
rect 487620 4208 487672 4214
rect 487620 4150 487672 4156
rect 486424 4004 486476 4010
rect 486424 3946 486476 3952
rect 485688 3052 485740 3058
rect 485688 2994 485740 3000
rect 485056 598 485268 626
rect 485056 490 485084 598
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 462 485084 490
rect 485240 480 485268 598
rect 486436 480 486464 3946
rect 487632 480 487660 4150
rect 488460 3126 488488 125598
rect 488828 125186 488856 128166
rect 488816 125180 488868 125186
rect 488816 125122 488868 125128
rect 488816 9036 488868 9042
rect 488816 8978 488868 8984
rect 488448 3120 488500 3126
rect 488448 3062 488500 3068
rect 488828 480 488856 8978
rect 489748 7614 489776 128166
rect 490576 125662 490604 128166
rect 491496 125934 491524 128166
rect 492416 126274 492444 128166
rect 492404 126268 492456 126274
rect 492404 126210 492456 126216
rect 491484 125928 491536 125934
rect 491484 125870 491536 125876
rect 493336 125662 493364 128166
rect 490564 125656 490616 125662
rect 490564 125598 490616 125604
rect 491208 125656 491260 125662
rect 491208 125598 491260 125604
rect 493324 125656 493376 125662
rect 493324 125598 493376 125604
rect 493968 125656 494020 125662
rect 493968 125598 494020 125604
rect 490012 89004 490064 89010
rect 490012 88946 490064 88952
rect 490024 16574 490052 88946
rect 490024 16546 490696 16574
rect 489736 7608 489788 7614
rect 489736 7550 489788 7556
rect 489920 3936 489972 3942
rect 489920 3878 489972 3884
rect 489932 480 489960 3878
rect 490668 490 490696 16546
rect 491220 3194 491248 125598
rect 492312 4616 492364 4622
rect 492312 4558 492364 4564
rect 491208 3188 491260 3194
rect 491208 3130 491260 3136
rect 490944 598 491156 626
rect 490944 490 490972 598
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 462 490972 490
rect 491128 480 491156 598
rect 492324 480 492352 4558
rect 493508 3868 493560 3874
rect 493508 3810 493560 3816
rect 493520 480 493548 3810
rect 493980 3262 494008 125598
rect 494256 125118 494284 128166
rect 494244 125112 494296 125118
rect 494244 125054 494296 125060
rect 494704 5228 494756 5234
rect 494704 5170 494756 5176
rect 493968 3256 494020 3262
rect 493968 3198 494020 3204
rect 494716 480 494744 5170
rect 495268 4078 495296 128166
rect 496096 125662 496124 128166
rect 496084 125656 496136 125662
rect 496084 125598 496136 125604
rect 496728 125656 496780 125662
rect 496728 125598 496780 125604
rect 495900 4752 495952 4758
rect 495900 4694 495952 4700
rect 495256 4072 495308 4078
rect 495256 4014 495308 4020
rect 495912 480 495940 4694
rect 496740 3330 496768 125598
rect 496924 125050 496952 128166
rect 496912 125044 496964 125050
rect 496912 124986 496964 124992
rect 498028 4146 498056 128166
rect 498764 125662 498792 128166
rect 498752 125656 498804 125662
rect 498752 125598 498804 125604
rect 499488 125656 499540 125662
rect 499488 125598 499540 125604
rect 499396 5364 499448 5370
rect 499396 5306 499448 5312
rect 498200 5092 498252 5098
rect 498200 5034 498252 5040
rect 498016 4140 498068 4146
rect 498016 4082 498068 4088
rect 497096 3800 497148 3806
rect 497096 3742 497148 3748
rect 496728 3324 496780 3330
rect 496728 3266 496780 3272
rect 497108 480 497136 3742
rect 498212 480 498240 5034
rect 499408 480 499436 5306
rect 499500 3398 499528 125598
rect 499684 124982 499712 128166
rect 499672 124976 499724 124982
rect 499672 124918 499724 124924
rect 500788 3874 500816 128166
rect 501524 125662 501552 128166
rect 501512 125656 501564 125662
rect 501512 125598 501564 125604
rect 502248 125656 502300 125662
rect 502248 125598 502300 125604
rect 501788 5160 501840 5166
rect 501788 5102 501840 5108
rect 500776 3868 500828 3874
rect 500776 3810 500828 3816
rect 500592 3732 500644 3738
rect 500592 3674 500644 3680
rect 499488 3392 499540 3398
rect 499488 3334 499540 3340
rect 500604 480 500632 3674
rect 501800 480 501828 5102
rect 502260 4010 502288 125598
rect 502444 124914 502472 128166
rect 502432 124908 502484 124914
rect 502432 124850 502484 124856
rect 502340 90364 502392 90370
rect 502340 90306 502392 90312
rect 502352 16574 502380 90306
rect 502352 16546 503024 16574
rect 502248 4004 502300 4010
rect 502248 3946 502300 3952
rect 502996 480 503024 16546
rect 503548 3806 503576 128166
rect 504192 125662 504220 128166
rect 505020 128166 505094 128194
rect 505986 128194 506014 128452
rect 506906 128194 506934 128452
rect 507826 128194 507854 128452
rect 505986 128166 506428 128194
rect 506906 128166 506980 128194
rect 504364 126064 504416 126070
rect 504364 126006 504416 126012
rect 504180 125656 504232 125662
rect 504180 125598 504232 125604
rect 504376 5098 504404 126006
rect 505020 125866 505048 128166
rect 505008 125860 505060 125866
rect 505008 125802 505060 125808
rect 505008 125656 505060 125662
rect 505008 125598 505060 125604
rect 504364 5092 504416 5098
rect 504364 5034 504416 5040
rect 505020 3942 505048 125598
rect 505376 5500 505428 5506
rect 505376 5442 505428 5448
rect 505008 3936 505060 3942
rect 505008 3878 505060 3884
rect 503536 3800 503588 3806
rect 503536 3742 503588 3748
rect 504180 3596 504232 3602
rect 504180 3538 504232 3544
rect 504192 480 504220 3538
rect 505388 480 505416 5442
rect 506400 3602 506428 128166
rect 506952 125662 506980 128166
rect 507688 128166 507854 128194
rect 508746 128194 508774 128452
rect 509574 128194 509602 128452
rect 510494 128194 510522 128452
rect 511414 128194 511442 128452
rect 512334 128194 512362 128452
rect 513254 128194 513282 128452
rect 508746 128166 509188 128194
rect 509574 128166 509648 128194
rect 510494 128166 510568 128194
rect 511414 128166 511488 128194
rect 512334 128166 512408 128194
rect 506940 125656 506992 125662
rect 506940 125598 506992 125604
rect 507688 123486 507716 128166
rect 507860 125928 507912 125934
rect 507860 125870 507912 125876
rect 507768 125656 507820 125662
rect 507768 125598 507820 125604
rect 507676 123480 507728 123486
rect 507676 123422 507728 123428
rect 506480 7676 506532 7682
rect 506480 7618 506532 7624
rect 506388 3596 506440 3602
rect 506388 3538 506440 3544
rect 506492 480 506520 7618
rect 507780 3738 507808 125598
rect 507872 125458 507900 125870
rect 507860 125452 507912 125458
rect 507860 125394 507912 125400
rect 507860 26920 507912 26926
rect 507860 26862 507912 26868
rect 507872 16574 507900 26862
rect 507872 16546 508912 16574
rect 507768 3732 507820 3738
rect 507768 3674 507820 3680
rect 507676 3664 507728 3670
rect 507676 3606 507728 3612
rect 507688 480 507716 3606
rect 508884 480 508912 16546
rect 509160 3670 509188 128166
rect 509620 125662 509648 128166
rect 510540 126070 510568 128166
rect 510528 126064 510580 126070
rect 510528 126006 510580 126012
rect 511460 125662 511488 128166
rect 512380 125662 512408 128166
rect 513208 128166 513282 128194
rect 514174 128194 514202 128452
rect 515108 128438 515444 128466
rect 514174 128166 514248 128194
rect 509608 125656 509660 125662
rect 509608 125598 509660 125604
rect 510528 125656 510580 125662
rect 510528 125598 510580 125604
rect 511448 125656 511500 125662
rect 511448 125598 511500 125604
rect 511908 125656 511960 125662
rect 511908 125598 511960 125604
rect 512368 125656 512420 125662
rect 512368 125598 512420 125604
rect 510068 5432 510120 5438
rect 510068 5374 510120 5380
rect 509148 3664 509200 3670
rect 509148 3606 509200 3612
rect 510080 480 510108 5374
rect 510540 3777 510568 125598
rect 510526 3768 510582 3777
rect 510526 3703 510582 3712
rect 511920 3534 511948 125598
rect 512460 4888 512512 4894
rect 512460 4830 512512 4836
rect 511264 3528 511316 3534
rect 511264 3470 511316 3476
rect 511908 3528 511960 3534
rect 511908 3470 511960 3476
rect 511276 480 511304 3470
rect 512472 480 512500 4830
rect 513208 3369 513236 128166
rect 514220 125662 514248 128166
rect 515416 125662 515444 128438
rect 519544 126880 519596 126886
rect 519544 126822 519596 126828
rect 517520 126812 517572 126818
rect 517520 126754 517572 126760
rect 513288 125656 513340 125662
rect 513288 125598 513340 125604
rect 514208 125656 514260 125662
rect 514208 125598 514260 125604
rect 514668 125656 514720 125662
rect 514668 125598 514720 125604
rect 515404 125656 515456 125662
rect 515404 125598 515456 125604
rect 516048 125656 516100 125662
rect 516048 125598 516100 125604
rect 513300 3641 513328 125598
rect 513564 5092 513616 5098
rect 513564 5034 513616 5040
rect 513286 3632 513342 3641
rect 513286 3567 513342 3576
rect 513194 3360 513250 3369
rect 513194 3295 513250 3304
rect 513576 480 513604 5034
rect 514680 3505 514708 125598
rect 515956 4956 516008 4962
rect 515956 4898 516008 4904
rect 514666 3496 514722 3505
rect 514666 3431 514722 3440
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 514772 480 514800 3402
rect 515968 480 515996 4898
rect 516060 3466 516088 125598
rect 517532 16574 517560 126754
rect 517532 16546 517928 16574
rect 517152 6248 517204 6254
rect 517152 6190 517204 6196
rect 516048 3460 516100 3466
rect 516048 3402 516100 3408
rect 517164 480 517192 6190
rect 517900 490 517928 16546
rect 519556 9654 519584 126822
rect 536104 126744 536156 126750
rect 536104 126686 536156 126692
rect 524420 126676 524472 126682
rect 524420 126618 524472 126624
rect 522304 126132 522356 126138
rect 522304 126074 522356 126080
rect 520924 125928 520976 125934
rect 520924 125870 520976 125876
rect 520280 10328 520332 10334
rect 520280 10270 520332 10276
rect 519544 9648 519596 9654
rect 519544 9590 519596 9596
rect 519544 8968 519596 8974
rect 519544 8910 519596 8916
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 8910
rect 520292 490 520320 10270
rect 520936 4214 520964 125870
rect 522316 4962 522344 126074
rect 524432 16574 524460 126618
rect 531320 126608 531372 126614
rect 531320 126550 531372 126556
rect 529204 126200 529256 126206
rect 529204 126142 529256 126148
rect 526444 125996 526496 126002
rect 526444 125938 526496 125944
rect 524432 16546 525472 16574
rect 524236 5024 524288 5030
rect 524236 4966 524288 4972
rect 522304 4956 522356 4962
rect 522304 4898 522356 4904
rect 520924 4208 520976 4214
rect 520924 4150 520976 4156
rect 523040 4208 523092 4214
rect 523040 4150 523092 4156
rect 521844 2848 521896 2854
rect 521844 2790 521896 2796
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 2790
rect 523052 480 523080 4150
rect 524248 480 524276 4966
rect 525444 480 525472 16546
rect 526456 8974 526484 125938
rect 526628 9648 526680 9654
rect 526628 9590 526680 9596
rect 526444 8968 526496 8974
rect 526444 8910 526496 8916
rect 526640 480 526668 9590
rect 527824 6180 527876 6186
rect 527824 6122 527876 6128
rect 527836 480 527864 6122
rect 529216 4894 529244 126142
rect 529940 125316 529992 125322
rect 529940 125258 529992 125264
rect 529952 16574 529980 125258
rect 531332 16574 531360 126550
rect 533344 126540 533396 126546
rect 533344 126482 533396 126488
rect 529952 16546 530164 16574
rect 531332 16546 532096 16574
rect 529204 4888 529256 4894
rect 529204 4830 529256 4836
rect 529020 2916 529072 2922
rect 529020 2858 529072 2864
rect 529032 480 529060 2858
rect 530136 480 530164 16546
rect 531320 4820 531372 4826
rect 531320 4762 531372 4768
rect 531332 480 531360 4762
rect 532068 490 532096 16546
rect 533356 4214 533384 126482
rect 533436 126064 533488 126070
rect 533436 126006 533488 126012
rect 533448 50386 533476 126006
rect 533436 50380 533488 50386
rect 533436 50322 533488 50328
rect 533712 4956 533764 4962
rect 533712 4898 533764 4904
rect 533344 4208 533396 4214
rect 533344 4150 533396 4156
rect 532344 598 532556 626
rect 532344 490 532372 598
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 462 532372 490
rect 532528 480 532556 598
rect 533724 480 533752 4898
rect 536116 4826 536144 126686
rect 547144 126472 547196 126478
rect 547144 126414 547196 126420
rect 543004 126404 543056 126410
rect 543004 126346 543056 126352
rect 539600 126336 539652 126342
rect 539600 126278 539652 126284
rect 536840 125384 536892 125390
rect 536840 125326 536892 125332
rect 536852 16574 536880 125326
rect 538220 125248 538272 125254
rect 538220 125190 538272 125196
rect 538232 16574 538260 125190
rect 536852 16546 537248 16574
rect 538232 16546 538444 16574
rect 536104 4820 536156 4826
rect 536104 4762 536156 4768
rect 534908 4208 534960 4214
rect 534908 4150 534960 4156
rect 534920 480 534948 4150
rect 536104 2984 536156 2990
rect 536104 2926 536156 2932
rect 536116 480 536144 2926
rect 537220 480 537248 16546
rect 538416 480 538444 16546
rect 539612 480 539640 126278
rect 540796 4888 540848 4894
rect 540796 4830 540848 4836
rect 540808 480 540836 4830
rect 541992 4820 542044 4826
rect 541992 4762 542044 4768
rect 542004 480 542032 4762
rect 543016 4214 543044 126346
rect 544384 8968 544436 8974
rect 544384 8910 544436 8916
rect 543004 4208 543056 4214
rect 543004 4150 543056 4156
rect 543188 3052 543240 3058
rect 543188 2994 543240 3000
rect 543200 480 543228 2994
rect 544396 480 544424 8910
rect 547156 4826 547184 126414
rect 568580 126268 568632 126274
rect 568580 126210 568632 126216
rect 550640 125452 550692 125458
rect 550640 125394 550692 125400
rect 547880 125180 547932 125186
rect 547880 125122 547932 125128
rect 547144 4820 547196 4826
rect 547144 4762 547196 4768
rect 545488 4208 545540 4214
rect 545488 4150 545540 4156
rect 545500 480 545528 4150
rect 546684 3120 546736 3126
rect 546684 3062 546736 3068
rect 546696 480 546724 3062
rect 547892 480 547920 125122
rect 550652 16574 550680 125394
rect 554780 125112 554832 125118
rect 554780 125054 554832 125060
rect 554792 16574 554820 125054
rect 557540 125044 557592 125050
rect 557540 124986 557592 124992
rect 557552 16574 557580 124986
rect 561680 124976 561732 124982
rect 561680 124918 561732 124924
rect 561692 16574 561720 124918
rect 564532 124908 564584 124914
rect 564532 124850 564584 124856
rect 564544 16574 564572 124850
rect 568592 16574 568620 126210
rect 572812 123480 572864 123486
rect 572812 123422 572864 123428
rect 550652 16546 551048 16574
rect 554792 16546 555004 16574
rect 557552 16546 558592 16574
rect 561692 16546 562088 16574
rect 564544 16546 565216 16574
rect 568592 16546 568712 16574
rect 549076 7608 549128 7614
rect 549076 7550 549128 7556
rect 549088 480 549116 7550
rect 550272 3188 550324 3194
rect 550272 3130 550324 3136
rect 550284 480 550312 3130
rect 551020 490 551048 16546
rect 552664 4820 552716 4826
rect 552664 4762 552716 4768
rect 551296 598 551508 626
rect 551296 490 551324 598
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 462 551324 490
rect 551480 480 551508 598
rect 552676 480 552704 4762
rect 553768 3256 553820 3262
rect 553768 3198 553820 3204
rect 553780 480 553808 3198
rect 554976 480 555004 16546
rect 556160 4072 556212 4078
rect 556160 4014 556212 4020
rect 556172 480 556200 4014
rect 557356 3324 557408 3330
rect 557356 3266 557408 3272
rect 557368 480 557396 3266
rect 558564 480 558592 16546
rect 559748 4140 559800 4146
rect 559748 4082 559800 4088
rect 559760 480 559788 4082
rect 560852 3392 560904 3398
rect 560852 3334 560904 3340
rect 560864 480 560892 3334
rect 562060 480 562088 16546
rect 564440 4004 564492 4010
rect 564440 3946 564492 3952
rect 563244 3868 563296 3874
rect 563244 3810 563296 3816
rect 563256 480 563284 3810
rect 564452 480 564480 3946
rect 565188 490 565216 16546
rect 568028 3936 568080 3942
rect 568028 3878 568080 3884
rect 566832 3800 566884 3806
rect 566832 3742 566884 3748
rect 565464 598 565676 626
rect 565464 490 565492 598
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 462 565492 490
rect 565648 480 565676 598
rect 566844 480 566872 3742
rect 568040 480 568068 3878
rect 568684 490 568712 16546
rect 572824 6914 572852 123422
rect 575480 50380 575532 50386
rect 575480 50322 575532 50328
rect 575492 16574 575520 50322
rect 575492 16546 575888 16574
rect 572732 6886 572852 6914
rect 571524 3732 571576 3738
rect 571524 3674 571576 3680
rect 570328 3596 570380 3602
rect 570328 3538 570380 3544
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 3538
rect 571536 480 571564 3674
rect 572732 480 572760 6886
rect 575110 3768 575166 3777
rect 575110 3703 575166 3712
rect 573916 3664 573968 3670
rect 573916 3606 573968 3612
rect 573928 480 573956 3606
rect 575124 480 575152 3703
rect 575860 490 575888 16546
rect 578606 3632 578662 3641
rect 578606 3567 578662 3576
rect 577412 3528 577464 3534
rect 577412 3470 577464 3476
rect 576136 598 576348 626
rect 576136 490 576164 598
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 462 576164 490
rect 576320 480 576348 598
rect 577424 480 577452 3470
rect 578620 480 578648 3567
rect 582194 3496 582250 3505
rect 582194 3431 582250 3440
rect 583392 3460 583444 3466
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582208 480 582236 3431
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3238 527856 3294 527912
rect 3330 514800 3386 514856
rect 3330 475632 3386 475688
rect 3330 462576 3386 462632
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 3330 371320 3386 371376
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3146 254088 3202 254144
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3974 566888 4030 566944
rect 3882 553832 3938 553888
rect 3790 501744 3846 501800
rect 3698 449520 3754 449576
rect 3606 397432 3662 397488
rect 21362 577088 21418 577144
rect 3514 293120 3570 293176
rect 3514 267144 3570 267200
rect 3514 241032 3570 241088
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 113822 576952 113878 577008
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 477958 577088 478014 577144
rect 526442 576952 526498 577008
rect 70214 574912 70270 574968
rect 73894 574912 73950 574968
rect 78402 574912 78458 574968
rect 82358 574912 82414 574968
rect 86314 574912 86370 574968
rect 90270 574912 90326 574968
rect 93674 574912 93730 574968
rect 97630 574912 97686 574968
rect 101954 574912 102010 574968
rect 105910 574912 105966 574968
rect 481914 574912 481970 574968
rect 485870 574912 485926 574968
rect 489918 574912 489974 574968
rect 493690 574912 493746 574968
rect 497554 574912 497610 574968
rect 501510 574912 501566 574968
rect 505466 574912 505522 574968
rect 509330 574912 509386 574968
rect 513930 574912 513986 574968
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 511264 580226 511320
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 579710 418240 579766 418296
rect 580170 378392 580226 378448
rect 579986 365064 580042 365120
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 579618 298696 579674 298752
rect 579894 272176 579950 272232
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 579894 219000 579950 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 579986 179152 580042 179208
rect 580906 537784 580962 537840
rect 580814 524456 580870 524512
rect 580722 484608 580778 484664
rect 580630 471416 580686 471472
rect 580538 431568 580594 431624
rect 580446 404912 580502 404968
rect 580354 351872 580410 351928
rect 580262 165824 580318 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 3238 136720 3294 136776
rect 3422 111696 3478 111752
rect 3422 110608 3478 110664
rect 3422 85448 3478 85504
rect 3422 84632 3478 84688
rect 3238 59200 3294 59256
rect 3238 58520 3294 58576
rect 3514 33088 3570 33144
rect 3514 32408 3570 32464
rect 3514 20576 3570 20632
rect 3514 19352 3570 19408
rect 13542 3304 13598 3360
rect 15934 3440 15990 3496
rect 71502 3576 71558 3632
rect 73802 3712 73858 3768
rect 78770 3168 78826 3224
rect 80886 3440 80942 3496
rect 80058 3304 80114 3360
rect 82082 3304 82138 3360
rect 122930 3576 122986 3632
rect 123298 3576 123354 3632
rect 124218 3712 124274 3768
rect 127070 3576 127126 3632
rect 129830 3440 129886 3496
rect 131210 3304 131266 3360
rect 412546 3712 412602 3768
rect 426346 3576 426402 3632
rect 431866 3440 431922 3496
rect 438766 3304 438822 3360
rect 447414 3712 447470 3768
rect 465170 3576 465226 3632
rect 472254 3440 472310 3496
rect 482834 3304 482890 3360
rect 510526 3712 510582 3768
rect 513286 3576 513342 3632
rect 513194 3304 513250 3360
rect 514666 3440 514722 3496
rect 575110 3712 575166 3768
rect 578606 3576 578662 3632
rect 582194 3440 582250 3496
rect 580998 3304 581054 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 21357 577146 21423 577149
rect 477953 577146 478019 577149
rect 21357 577144 478019 577146
rect 21357 577088 21362 577144
rect 21418 577088 477958 577144
rect 478014 577088 478019 577144
rect 21357 577086 478019 577088
rect 21357 577083 21423 577086
rect 477953 577083 478019 577086
rect 113817 577010 113883 577013
rect 526437 577010 526503 577013
rect 113817 577008 526503 577010
rect 113817 576952 113822 577008
rect 113878 576952 526442 577008
rect 526498 576952 526503 577008
rect 113817 576950 526503 576952
rect 113817 576947 113883 576950
rect 526437 576947 526503 576950
rect 70209 574972 70275 574973
rect 70158 574970 70164 574972
rect 70118 574910 70164 574970
rect 70228 574968 70275 574972
rect 70270 574912 70275 574968
rect 70158 574908 70164 574910
rect 70228 574908 70275 574912
rect 73470 574908 73476 574972
rect 73540 574970 73546 574972
rect 73889 574970 73955 574973
rect 73540 574968 73955 574970
rect 73540 574912 73894 574968
rect 73950 574912 73955 574968
rect 73540 574910 73955 574912
rect 73540 574908 73546 574910
rect 70209 574907 70275 574908
rect 73889 574907 73955 574910
rect 78397 574972 78463 574973
rect 78397 574968 78444 574972
rect 78508 574970 78514 574972
rect 82353 574970 82419 574973
rect 82670 574970 82676 574972
rect 78397 574912 78402 574968
rect 78397 574908 78444 574912
rect 78508 574910 78554 574970
rect 82353 574968 82676 574970
rect 82353 574912 82358 574968
rect 82414 574912 82676 574968
rect 82353 574910 82676 574912
rect 78508 574908 78514 574910
rect 78397 574907 78463 574908
rect 82353 574907 82419 574910
rect 82670 574908 82676 574910
rect 82740 574908 82746 574972
rect 86309 574970 86375 574973
rect 86718 574970 86724 574972
rect 86309 574968 86724 574970
rect 86309 574912 86314 574968
rect 86370 574912 86724 574968
rect 86309 574910 86724 574912
rect 86309 574907 86375 574910
rect 86718 574908 86724 574910
rect 86788 574908 86794 574972
rect 90265 574970 90331 574973
rect 93669 574972 93735 574973
rect 90950 574970 90956 574972
rect 90265 574968 90956 574970
rect 90265 574912 90270 574968
rect 90326 574912 90956 574968
rect 90265 574910 90956 574912
rect 90265 574907 90331 574910
rect 90950 574908 90956 574910
rect 91020 574908 91026 574972
rect 93669 574968 93716 574972
rect 93780 574970 93786 574972
rect 97625 574970 97691 574973
rect 101949 574972 102015 574973
rect 97758 574970 97764 574972
rect 93669 574912 93674 574968
rect 93669 574908 93716 574912
rect 93780 574910 93826 574970
rect 97625 574968 97764 574970
rect 97625 574912 97630 574968
rect 97686 574912 97764 574968
rect 97625 574910 97764 574912
rect 93780 574908 93786 574910
rect 93669 574907 93735 574908
rect 97625 574907 97691 574910
rect 97758 574908 97764 574910
rect 97828 574908 97834 574972
rect 101949 574968 101996 574972
rect 102060 574970 102066 574972
rect 105905 574970 105971 574973
rect 106038 574970 106044 574972
rect 101949 574912 101954 574968
rect 101949 574908 101996 574912
rect 102060 574910 102106 574970
rect 105905 574968 106044 574970
rect 105905 574912 105910 574968
rect 105966 574912 106044 574968
rect 105905 574910 106044 574912
rect 102060 574908 102066 574910
rect 101949 574907 102015 574908
rect 105905 574907 105971 574910
rect 106038 574908 106044 574910
rect 106108 574908 106114 574972
rect 481766 574908 481772 574972
rect 481836 574970 481842 574972
rect 481909 574970 481975 574973
rect 485865 574972 485931 574973
rect 489913 574972 489979 574973
rect 485814 574970 485820 574972
rect 481836 574968 481975 574970
rect 481836 574912 481914 574968
rect 481970 574912 481975 574968
rect 481836 574910 481975 574912
rect 485774 574910 485820 574970
rect 485884 574968 485931 574972
rect 485926 574912 485931 574968
rect 481836 574908 481842 574910
rect 481909 574907 481975 574910
rect 485814 574908 485820 574910
rect 485884 574908 485931 574912
rect 489862 574908 489868 574972
rect 489932 574970 489979 574972
rect 489932 574968 490024 574970
rect 489974 574912 490024 574968
rect 489932 574910 490024 574912
rect 489932 574908 489979 574910
rect 492806 574908 492812 574972
rect 492876 574970 492882 574972
rect 493685 574970 493751 574973
rect 492876 574968 493751 574970
rect 492876 574912 493690 574968
rect 493746 574912 493751 574968
rect 492876 574910 493751 574912
rect 492876 574908 492882 574910
rect 485865 574907 485931 574908
rect 489913 574907 489979 574908
rect 493685 574907 493751 574910
rect 496854 574908 496860 574972
rect 496924 574970 496930 574972
rect 497549 574970 497615 574973
rect 496924 574968 497615 574970
rect 496924 574912 497554 574968
rect 497610 574912 497615 574968
rect 496924 574910 497615 574912
rect 496924 574908 496930 574910
rect 497549 574907 497615 574910
rect 500902 574908 500908 574972
rect 500972 574970 500978 574972
rect 501505 574970 501571 574973
rect 500972 574968 501571 574970
rect 500972 574912 501510 574968
rect 501566 574912 501571 574968
rect 500972 574910 501571 574912
rect 500972 574908 500978 574910
rect 501505 574907 501571 574910
rect 505134 574908 505140 574972
rect 505204 574970 505210 574972
rect 505461 574970 505527 574973
rect 505204 574968 505527 574970
rect 505204 574912 505466 574968
rect 505522 574912 505527 574968
rect 505204 574910 505527 574912
rect 505204 574908 505210 574910
rect 505461 574907 505527 574910
rect 509182 574908 509188 574972
rect 509252 574970 509258 574972
rect 509325 574970 509391 574973
rect 509252 574968 509391 574970
rect 509252 574912 509330 574968
rect 509386 574912 509391 574968
rect 509252 574910 509391 574912
rect 509252 574908 509258 574910
rect 509325 574907 509391 574910
rect 513925 574972 513991 574973
rect 513925 574968 513972 574972
rect 514036 574970 514042 574972
rect 513925 574912 513930 574968
rect 513925 574908 513972 574912
rect 514036 574910 514082 574970
rect 514036 574908 514042 574910
rect 513925 574907 513991 574908
rect -960 566946 480 567036
rect 3969 566946 4035 566949
rect -960 566944 4035 566946
rect -960 566888 3974 566944
rect 4030 566888 4035 566944
rect -960 566886 4035 566888
rect -960 566796 480 566886
rect 3969 566883 4035 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3877 553890 3943 553893
rect -960 553888 3943 553890
rect -960 553832 3882 553888
rect 3938 553832 3943 553888
rect -960 553830 3943 553832
rect -960 553740 480 553830
rect 3877 553827 3943 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3233 527914 3299 527917
rect -960 527912 3299 527914
rect -960 527856 3238 527912
rect 3294 527856 3299 527912
rect -960 527854 3299 527856
rect -960 527764 480 527854
rect 3233 527851 3299 527854
rect 580809 524514 580875 524517
rect 583520 524514 584960 524604
rect 580809 524512 584960 524514
rect 580809 524456 580814 524512
rect 580870 524456 584960 524512
rect 580809 524454 584960 524456
rect 580809 524451 580875 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580717 484666 580783 484669
rect 583520 484666 584960 484756
rect 580717 484664 584960 484666
rect 580717 484608 580722 484664
rect 580778 484608 584960 484664
rect 580717 484606 584960 484608
rect 580717 484603 580783 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 580625 471474 580691 471477
rect 583520 471474 584960 471564
rect 580625 471472 584960 471474
rect 580625 471416 580630 471472
rect 580686 471416 584960 471472
rect 580625 471414 584960 471416
rect 580625 471411 580691 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3693 449578 3759 449581
rect -960 449576 3759 449578
rect -960 449520 3698 449576
rect 3754 449520 3759 449576
rect -960 449518 3759 449520
rect -960 449428 480 449518
rect 3693 449515 3759 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580533 431626 580599 431629
rect 583520 431626 584960 431716
rect 580533 431624 584960 431626
rect 580533 431568 580538 431624
rect 580594 431568 584960 431624
rect 580533 431566 584960 431568
rect 580533 431563 580599 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580441 404970 580507 404973
rect 583520 404970 584960 405060
rect 580441 404968 584960 404970
rect 580441 404912 580446 404968
rect 580502 404912 584960 404968
rect 580441 404910 584960 404912
rect 580441 404907 580507 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3601 397490 3667 397493
rect -960 397488 3667 397490
rect -960 397432 3606 397488
rect 3662 397432 3667 397488
rect -960 397430 3667 397432
rect -960 397340 480 397430
rect 3601 397427 3667 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 579981 365122 580047 365125
rect 583520 365122 584960 365212
rect 579981 365120 584960 365122
rect 579981 365064 579986 365120
rect 580042 365064 584960 365120
rect 579981 365062 584960 365064
rect 579981 365059 580047 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580257 165882 580323 165885
rect 583520 165882 584960 165972
rect 580257 165880 584960 165882
rect 580257 165824 580262 165880
rect 580318 165824 584960 165880
rect 580257 165822 584960 165824
rect 580257 165819 580323 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 106038 125564 106044 125628
rect 106108 125626 106114 125628
rect 583526 125626 583586 125838
rect 106108 125566 583586 125626
rect 106108 125564 106114 125566
rect -960 123572 480 123812
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 97758 111828 97764 111892
rect 97828 111890 97834 111892
rect 583526 111890 583586 112646
rect 97828 111830 583586 111890
rect 97828 111828 97834 111830
rect 3417 111754 3483 111757
rect 481766 111754 481772 111756
rect 3417 111752 481772 111754
rect 3417 111696 3422 111752
rect 3478 111696 481772 111752
rect 3417 111694 481772 111696
rect 3417 111691 3483 111694
rect 481766 111692 481772 111694
rect 481836 111692 481842 111756
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 101990 99452 101996 99516
rect 102060 99514 102066 99516
rect 583520 99514 584960 99604
rect 102060 99454 584960 99514
rect 102060 99452 102066 99454
rect 583520 99364 584960 99454
rect 489678 97882 489684 97884
rect 6870 97822 489684 97882
rect -960 97610 480 97700
rect 6870 97610 6930 97822
rect 489678 97820 489684 97822
rect 489748 97820 489754 97884
rect -960 97550 6930 97610
rect -960 97460 480 97550
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 93710 85580 93716 85644
rect 93780 85642 93786 85644
rect 583526 85642 583586 85990
rect 93780 85582 583586 85642
rect 93780 85580 93786 85582
rect 3417 85506 3483 85509
rect 485814 85506 485820 85508
rect 3417 85504 485820 85506
rect 3417 85448 3422 85504
rect 3478 85448 485820 85504
rect 3417 85446 485820 85448
rect 3417 85443 3483 85446
rect 485814 85444 485820 85446
rect 485884 85444 485890 85508
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 86718 71844 86724 71908
rect 86788 71906 86794 71908
rect 583526 71906 583586 72798
rect 86788 71846 583586 71906
rect 86788 71844 86794 71846
rect 492806 71770 492812 71772
rect -960 71634 480 71724
rect 6870 71710 492812 71770
rect 6870 71634 6930 71710
rect 492806 71708 492812 71710
rect 492876 71708 492882 71772
rect -960 71574 6930 71634
rect -960 71484 480 71574
rect 583520 59666 584960 59756
rect 567150 59606 584960 59666
rect 90950 59332 90956 59396
rect 91020 59394 91026 59396
rect 567150 59394 567210 59606
rect 583520 59516 584960 59606
rect 91020 59334 567210 59394
rect 91020 59332 91026 59334
rect 3233 59258 3299 59261
rect 500902 59258 500908 59260
rect 3233 59256 500908 59258
rect 3233 59200 3238 59256
rect 3294 59200 500908 59256
rect 3233 59198 500908 59200
rect 3233 59195 3299 59198
rect 500902 59196 500908 59198
rect 500972 59196 500978 59260
rect -960 58578 480 58668
rect 3233 58578 3299 58581
rect -960 58576 3299 58578
rect -960 58520 3238 58576
rect 3294 58520 3299 58576
rect -960 58518 3299 58520
rect -960 58428 480 58518
rect 3233 58515 3299 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 82670 45596 82676 45660
rect 82740 45658 82746 45660
rect 583526 45658 583586 46142
rect 82740 45598 583586 45658
rect 82740 45596 82746 45598
rect 496854 45522 496860 45524
rect -960 45462 496860 45522
rect -960 45372 480 45462
rect 496854 45460 496860 45462
rect 496924 45460 496930 45524
rect 3509 33146 3575 33149
rect 505134 33146 505140 33148
rect 3509 33144 505140 33146
rect 3509 33088 3514 33144
rect 3570 33088 505140 33144
rect 3509 33086 505140 33088
rect 3509 33083 3575 33086
rect 505134 33084 505140 33086
rect 505204 33084 505210 33148
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 73470 31724 73476 31788
rect 73540 31786 73546 31788
rect 583526 31786 583586 32950
rect 73540 31726 583586 31786
rect 73540 31724 73546 31726
rect 3509 20634 3575 20637
rect 513966 20634 513972 20636
rect 3509 20632 513972 20634
rect 3509 20576 3514 20632
rect 3570 20576 513972 20632
rect 3509 20574 513972 20576
rect 3509 20571 3575 20574
rect 513966 20572 513972 20574
rect 514036 20572 514042 20636
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 78438 19348 78444 19412
rect 78508 19410 78514 19412
rect 583526 19410 583586 19622
rect 78508 19350 583586 19410
rect 78508 19348 78514 19350
rect 509182 6898 509188 6900
rect 6870 6838 509188 6898
rect -960 6490 480 6580
rect 6870 6490 6930 6838
rect 509182 6836 509188 6838
rect 509252 6836 509258 6900
rect 583520 6626 584960 6716
rect -960 6430 6930 6490
rect 583342 6566 584960 6626
rect 583342 6490 583402 6566
rect 583520 6490 584960 6566
rect 583342 6476 584960 6490
rect 583342 6430 583586 6476
rect -960 6340 480 6430
rect 70158 5612 70164 5676
rect 70228 5674 70234 5676
rect 583526 5674 583586 6430
rect 70228 5614 583586 5674
rect 70228 5612 70234 5614
rect 73797 3770 73863 3773
rect 124213 3770 124279 3773
rect 73797 3768 124279 3770
rect 73797 3712 73802 3768
rect 73858 3712 124218 3768
rect 124274 3712 124279 3768
rect 73797 3710 124279 3712
rect 73797 3707 73863 3710
rect 124213 3707 124279 3710
rect 412541 3770 412607 3773
rect 447409 3770 447475 3773
rect 412541 3768 447475 3770
rect 412541 3712 412546 3768
rect 412602 3712 447414 3768
rect 447470 3712 447475 3768
rect 412541 3710 447475 3712
rect 412541 3707 412607 3710
rect 447409 3707 447475 3710
rect 510521 3770 510587 3773
rect 575105 3770 575171 3773
rect 510521 3768 575171 3770
rect 510521 3712 510526 3768
rect 510582 3712 575110 3768
rect 575166 3712 575171 3768
rect 510521 3710 575171 3712
rect 510521 3707 510587 3710
rect 575105 3707 575171 3710
rect 71497 3634 71563 3637
rect 122925 3634 122991 3637
rect 71497 3632 122991 3634
rect 71497 3576 71502 3632
rect 71558 3576 122930 3632
rect 122986 3576 122991 3632
rect 71497 3574 122991 3576
rect 71497 3571 71563 3574
rect 122925 3571 122991 3574
rect 123293 3634 123359 3637
rect 127065 3634 127131 3637
rect 123293 3632 127131 3634
rect 123293 3576 123298 3632
rect 123354 3576 127070 3632
rect 127126 3576 127131 3632
rect 123293 3574 127131 3576
rect 123293 3571 123359 3574
rect 127065 3571 127131 3574
rect 426341 3634 426407 3637
rect 465165 3634 465231 3637
rect 426341 3632 465231 3634
rect 426341 3576 426346 3632
rect 426402 3576 465170 3632
rect 465226 3576 465231 3632
rect 426341 3574 465231 3576
rect 426341 3571 426407 3574
rect 465165 3571 465231 3574
rect 513281 3634 513347 3637
rect 578601 3634 578667 3637
rect 513281 3632 578667 3634
rect 513281 3576 513286 3632
rect 513342 3576 578606 3632
rect 578662 3576 578667 3632
rect 513281 3574 578667 3576
rect 513281 3571 513347 3574
rect 578601 3571 578667 3574
rect 15929 3498 15995 3501
rect 80881 3498 80947 3501
rect 129825 3498 129891 3501
rect 15929 3496 74826 3498
rect 15929 3440 15934 3496
rect 15990 3440 74826 3496
rect 15929 3438 74826 3440
rect 15929 3435 15995 3438
rect 13537 3362 13603 3365
rect 74766 3362 74826 3438
rect 80881 3496 129891 3498
rect 80881 3440 80886 3496
rect 80942 3440 129830 3496
rect 129886 3440 129891 3496
rect 80881 3438 129891 3440
rect 80881 3435 80947 3438
rect 129825 3435 129891 3438
rect 431861 3498 431927 3501
rect 472249 3498 472315 3501
rect 431861 3496 472315 3498
rect 431861 3440 431866 3496
rect 431922 3440 472254 3496
rect 472310 3440 472315 3496
rect 431861 3438 472315 3440
rect 431861 3435 431927 3438
rect 472249 3435 472315 3438
rect 514661 3498 514727 3501
rect 582189 3498 582255 3501
rect 514661 3496 582255 3498
rect 514661 3440 514666 3496
rect 514722 3440 582194 3496
rect 582250 3440 582255 3496
rect 514661 3438 582255 3440
rect 514661 3435 514727 3438
rect 582189 3435 582255 3438
rect 80053 3362 80119 3365
rect 13537 3360 74642 3362
rect 13537 3304 13542 3360
rect 13598 3304 74642 3360
rect 13537 3302 74642 3304
rect 74766 3360 80119 3362
rect 74766 3304 80058 3360
rect 80114 3304 80119 3360
rect 74766 3302 80119 3304
rect 13537 3299 13603 3302
rect 74582 3226 74642 3302
rect 80053 3299 80119 3302
rect 82077 3362 82143 3365
rect 131205 3362 131271 3365
rect 82077 3360 131271 3362
rect 82077 3304 82082 3360
rect 82138 3304 131210 3360
rect 131266 3304 131271 3360
rect 82077 3302 131271 3304
rect 82077 3299 82143 3302
rect 131205 3299 131271 3302
rect 438761 3362 438827 3365
rect 482829 3362 482895 3365
rect 438761 3360 482895 3362
rect 438761 3304 438766 3360
rect 438822 3304 482834 3360
rect 482890 3304 482895 3360
rect 438761 3302 482895 3304
rect 438761 3299 438827 3302
rect 482829 3299 482895 3302
rect 513189 3362 513255 3365
rect 580993 3362 581059 3365
rect 513189 3360 581059 3362
rect 513189 3304 513194 3360
rect 513250 3304 580998 3360
rect 581054 3304 581059 3360
rect 513189 3302 581059 3304
rect 513189 3299 513255 3302
rect 580993 3299 581059 3302
rect 78765 3226 78831 3229
rect 74582 3224 78831 3226
rect 74582 3168 78770 3224
rect 78826 3168 78831 3224
rect 74582 3166 78831 3168
rect 78765 3163 78831 3166
<< via3 >>
rect 70164 574968 70228 574972
rect 70164 574912 70214 574968
rect 70214 574912 70228 574968
rect 70164 574908 70228 574912
rect 73476 574908 73540 574972
rect 78444 574968 78508 574972
rect 78444 574912 78458 574968
rect 78458 574912 78508 574968
rect 78444 574908 78508 574912
rect 82676 574908 82740 574972
rect 86724 574908 86788 574972
rect 90956 574908 91020 574972
rect 93716 574968 93780 574972
rect 93716 574912 93730 574968
rect 93730 574912 93780 574968
rect 93716 574908 93780 574912
rect 97764 574908 97828 574972
rect 101996 574968 102060 574972
rect 101996 574912 102010 574968
rect 102010 574912 102060 574968
rect 101996 574908 102060 574912
rect 106044 574908 106108 574972
rect 481772 574908 481836 574972
rect 485820 574968 485884 574972
rect 485820 574912 485870 574968
rect 485870 574912 485884 574968
rect 485820 574908 485884 574912
rect 489868 574968 489932 574972
rect 489868 574912 489918 574968
rect 489918 574912 489932 574968
rect 489868 574908 489932 574912
rect 492812 574908 492876 574972
rect 496860 574908 496924 574972
rect 500908 574908 500972 574972
rect 505140 574908 505204 574972
rect 509188 574908 509252 574972
rect 513972 574968 514036 574972
rect 513972 574912 513986 574968
rect 513986 574912 514036 574968
rect 513972 574908 514036 574912
rect 106044 125564 106108 125628
rect 97764 111828 97828 111892
rect 481772 111692 481836 111756
rect 101996 99452 102060 99516
rect 489684 97820 489748 97884
rect 93716 85580 93780 85644
rect 485820 85444 485884 85508
rect 86724 71844 86788 71908
rect 492812 71708 492876 71772
rect 90956 59332 91020 59396
rect 500908 59196 500972 59260
rect 82676 45596 82740 45660
rect 496860 45460 496924 45524
rect 505140 33084 505204 33148
rect 73476 31724 73540 31788
rect 513972 20572 514036 20636
rect 78444 19348 78508 19412
rect 509188 6836 509252 6900
rect 70164 5612 70228 5676
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 577600 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 577600 74414 578898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 577600 78134 582618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 577600 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 577600 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 577600 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 577600 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 577600 99854 604338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 577600 103574 608058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 577600 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 577600 114134 582618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 577600 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 577600 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 577600 128414 596898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 577600 132134 600618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 577600 135854 604338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 577600 139574 608058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 577600 146414 578898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 577600 150134 582618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 577600 153854 586338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 577600 157574 590058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 577600 164414 596898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 577600 168134 600618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 577600 171854 604338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 577600 175574 608058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 577600 182414 578898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 577600 186134 582618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 577600 189854 586338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 577600 193574 590058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 577600 200414 596898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 577600 204134 600618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 577600 207854 604338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 577600 211574 608058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 577600 218414 578898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 577600 222134 582618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 577600 225854 586338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 577600 229574 590058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 577600 236414 596898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 577600 240134 600618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 577600 243854 604338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 577600 247574 608058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 577600 254414 578898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 577600 258134 582618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 577600 261854 586338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 577600 265574 590058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 577600 272414 596898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 577600 276134 600618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 577600 279854 604338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 577600 283574 608058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 577600 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 577600 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 577600 297854 586338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 577600 301574 590058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 577600 308414 596898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 577600 312134 600618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 577600 315854 604338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 577600 319574 608058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 577600 326414 578898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 577600 330134 582618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 577600 333854 586338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 577600 337574 590058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 577600 344414 596898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 577600 348134 600618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 577600 351854 604338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 577600 355574 608058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 577600 362414 578898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 577600 366134 582618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 577600 369854 586338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 577600 373574 590058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 577600 380414 596898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 577600 384134 600618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 577600 387854 604338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 577600 391574 608058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 577600 398414 578898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 577600 402134 582618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 577600 405854 586338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 577600 409574 590058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 577600 416414 596898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 577600 420134 600618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 577600 423854 604338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 577600 427574 608058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 577600 434414 578898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 577600 438134 582618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 577600 441854 586338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 577600 445574 590058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 577600 452414 596898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 577600 456134 600618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 577600 459854 604338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 577600 463574 608058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 577600 470414 578898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 577600 474134 582618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 577600 477854 586338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 577600 481574 590058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 577600 488414 596898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 577600 492134 600618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 577600 495854 604338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 577600 499574 608058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 577600 506414 578898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 577600 510134 582618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 577600 513854 586338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 577600 517574 590058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 70163 574972 70229 574973
rect 70163 574908 70164 574972
rect 70228 574908 70229 574972
rect 70163 574907 70229 574908
rect 73475 574972 73541 574973
rect 73475 574908 73476 574972
rect 73540 574908 73541 574972
rect 73475 574907 73541 574908
rect 78443 574972 78509 574973
rect 78443 574908 78444 574972
rect 78508 574908 78509 574972
rect 78443 574907 78509 574908
rect 82675 574972 82741 574973
rect 82675 574908 82676 574972
rect 82740 574908 82741 574972
rect 82675 574907 82741 574908
rect 86723 574972 86789 574973
rect 86723 574908 86724 574972
rect 86788 574908 86789 574972
rect 86723 574907 86789 574908
rect 90955 574972 91021 574973
rect 90955 574908 90956 574972
rect 91020 574908 91021 574972
rect 90955 574907 91021 574908
rect 93715 574972 93781 574973
rect 93715 574908 93716 574972
rect 93780 574908 93781 574972
rect 93715 574907 93781 574908
rect 97763 574972 97829 574973
rect 97763 574908 97764 574972
rect 97828 574908 97829 574972
rect 97763 574907 97829 574908
rect 101995 574972 102061 574973
rect 101995 574908 101996 574972
rect 102060 574908 102061 574972
rect 101995 574907 102061 574908
rect 106043 574972 106109 574973
rect 106043 574908 106044 574972
rect 106108 574908 106109 574972
rect 106043 574907 106109 574908
rect 481771 574972 481837 574973
rect 481771 574908 481772 574972
rect 481836 574908 481837 574972
rect 481771 574907 481837 574908
rect 485819 574972 485885 574973
rect 485819 574908 485820 574972
rect 485884 574908 485885 574972
rect 489867 574972 489933 574973
rect 489867 574970 489868 574972
rect 485819 574907 485885 574908
rect 489686 574910 489868 574970
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 104614 67574 126400
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 70166 5677 70226 574907
rect 72608 543454 72928 543486
rect 72608 543218 72650 543454
rect 72886 543218 72928 543454
rect 72608 543134 72928 543218
rect 72608 542898 72650 543134
rect 72886 542898 72928 543134
rect 72608 542866 72928 542898
rect 72608 507454 72928 507486
rect 72608 507218 72650 507454
rect 72886 507218 72928 507454
rect 72608 507134 72928 507218
rect 72608 506898 72650 507134
rect 72886 506898 72928 507134
rect 72608 506866 72928 506898
rect 72608 471454 72928 471486
rect 72608 471218 72650 471454
rect 72886 471218 72928 471454
rect 72608 471134 72928 471218
rect 72608 470898 72650 471134
rect 72886 470898 72928 471134
rect 72608 470866 72928 470898
rect 72608 435454 72928 435486
rect 72608 435218 72650 435454
rect 72886 435218 72928 435454
rect 72608 435134 72928 435218
rect 72608 434898 72650 435134
rect 72886 434898 72928 435134
rect 72608 434866 72928 434898
rect 72608 399454 72928 399486
rect 72608 399218 72650 399454
rect 72886 399218 72928 399454
rect 72608 399134 72928 399218
rect 72608 398898 72650 399134
rect 72886 398898 72928 399134
rect 72608 398866 72928 398898
rect 72608 363454 72928 363486
rect 72608 363218 72650 363454
rect 72886 363218 72928 363454
rect 72608 363134 72928 363218
rect 72608 362898 72650 363134
rect 72886 362898 72928 363134
rect 72608 362866 72928 362898
rect 72608 327454 72928 327486
rect 72608 327218 72650 327454
rect 72886 327218 72928 327454
rect 72608 327134 72928 327218
rect 72608 326898 72650 327134
rect 72886 326898 72928 327134
rect 72608 326866 72928 326898
rect 72608 291454 72928 291486
rect 72608 291218 72650 291454
rect 72886 291218 72928 291454
rect 72608 291134 72928 291218
rect 72608 290898 72650 291134
rect 72886 290898 72928 291134
rect 72608 290866 72928 290898
rect 72608 255454 72928 255486
rect 72608 255218 72650 255454
rect 72886 255218 72928 255454
rect 72608 255134 72928 255218
rect 72608 254898 72650 255134
rect 72886 254898 72928 255134
rect 72608 254866 72928 254898
rect 72608 219454 72928 219486
rect 72608 219218 72650 219454
rect 72886 219218 72928 219454
rect 72608 219134 72928 219218
rect 72608 218898 72650 219134
rect 72886 218898 72928 219134
rect 72608 218866 72928 218898
rect 72608 183454 72928 183486
rect 72608 183218 72650 183454
rect 72886 183218 72928 183454
rect 72608 183134 72928 183218
rect 72608 182898 72650 183134
rect 72886 182898 72928 183134
rect 72608 182866 72928 182898
rect 72608 147454 72928 147486
rect 72608 147218 72650 147454
rect 72886 147218 72928 147454
rect 72608 147134 72928 147218
rect 72608 146898 72650 147134
rect 72886 146898 72928 147134
rect 72608 146866 72928 146898
rect 73478 31789 73538 574907
rect 73794 111454 74414 126400
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73475 31788 73541 31789
rect 73475 31724 73476 31788
rect 73540 31724 73541 31788
rect 73475 31723 73541 31724
rect 70163 5676 70229 5677
rect 70163 5612 70164 5676
rect 70228 5612 70229 5676
rect 70163 5611 70229 5612
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 115174 78134 126400
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 78446 19413 78506 574907
rect 81234 118894 81854 126400
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 78443 19412 78509 19413
rect 78443 19348 78444 19412
rect 78508 19348 78509 19412
rect 78443 19347 78509 19348
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 46338
rect 82678 45661 82738 574907
rect 84954 122614 85574 126400
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 86726 71909 86786 574907
rect 87968 561454 88288 561486
rect 87968 561218 88010 561454
rect 88246 561218 88288 561454
rect 87968 561134 88288 561218
rect 87968 560898 88010 561134
rect 88246 560898 88288 561134
rect 87968 560866 88288 560898
rect 87968 525454 88288 525486
rect 87968 525218 88010 525454
rect 88246 525218 88288 525454
rect 87968 525134 88288 525218
rect 87968 524898 88010 525134
rect 88246 524898 88288 525134
rect 87968 524866 88288 524898
rect 87968 489454 88288 489486
rect 87968 489218 88010 489454
rect 88246 489218 88288 489454
rect 87968 489134 88288 489218
rect 87968 488898 88010 489134
rect 88246 488898 88288 489134
rect 87968 488866 88288 488898
rect 87968 453454 88288 453486
rect 87968 453218 88010 453454
rect 88246 453218 88288 453454
rect 87968 453134 88288 453218
rect 87968 452898 88010 453134
rect 88246 452898 88288 453134
rect 87968 452866 88288 452898
rect 87968 417454 88288 417486
rect 87968 417218 88010 417454
rect 88246 417218 88288 417454
rect 87968 417134 88288 417218
rect 87968 416898 88010 417134
rect 88246 416898 88288 417134
rect 87968 416866 88288 416898
rect 87968 381454 88288 381486
rect 87968 381218 88010 381454
rect 88246 381218 88288 381454
rect 87968 381134 88288 381218
rect 87968 380898 88010 381134
rect 88246 380898 88288 381134
rect 87968 380866 88288 380898
rect 87968 345454 88288 345486
rect 87968 345218 88010 345454
rect 88246 345218 88288 345454
rect 87968 345134 88288 345218
rect 87968 344898 88010 345134
rect 88246 344898 88288 345134
rect 87968 344866 88288 344898
rect 87968 309454 88288 309486
rect 87968 309218 88010 309454
rect 88246 309218 88288 309454
rect 87968 309134 88288 309218
rect 87968 308898 88010 309134
rect 88246 308898 88288 309134
rect 87968 308866 88288 308898
rect 87968 273454 88288 273486
rect 87968 273218 88010 273454
rect 88246 273218 88288 273454
rect 87968 273134 88288 273218
rect 87968 272898 88010 273134
rect 88246 272898 88288 273134
rect 87968 272866 88288 272898
rect 87968 237454 88288 237486
rect 87968 237218 88010 237454
rect 88246 237218 88288 237454
rect 87968 237134 88288 237218
rect 87968 236898 88010 237134
rect 88246 236898 88288 237134
rect 87968 236866 88288 236898
rect 87968 201454 88288 201486
rect 87968 201218 88010 201454
rect 88246 201218 88288 201454
rect 87968 201134 88288 201218
rect 87968 200898 88010 201134
rect 88246 200898 88288 201134
rect 87968 200866 88288 200898
rect 87968 165454 88288 165486
rect 87968 165218 88010 165454
rect 88246 165218 88288 165454
rect 87968 165134 88288 165218
rect 87968 164898 88010 165134
rect 88246 164898 88288 165134
rect 87968 164866 88288 164898
rect 86723 71908 86789 71909
rect 86723 71844 86724 71908
rect 86788 71844 86789 71908
rect 86723 71843 86789 71844
rect 90958 59397 91018 574907
rect 91794 93454 92414 126400
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 90955 59396 91021 59397
rect 90955 59332 90956 59396
rect 91020 59332 91021 59396
rect 90955 59331 91021 59332
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 82675 45660 82741 45661
rect 82675 45596 82676 45660
rect 82740 45596 82741 45660
rect 82675 45595 82741 45596
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 92898
rect 93718 85645 93778 574907
rect 95514 97174 96134 126400
rect 97766 111893 97826 574907
rect 97763 111892 97829 111893
rect 97763 111828 97764 111892
rect 97828 111828 97829 111892
rect 97763 111827 97829 111828
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 93715 85644 93781 85645
rect 93715 85580 93716 85644
rect 93780 85580 93781 85644
rect 93715 85579 93781 85580
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 100894 99854 126400
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 101998 99517 102058 574907
rect 103328 543454 103648 543486
rect 103328 543218 103370 543454
rect 103606 543218 103648 543454
rect 103328 543134 103648 543218
rect 103328 542898 103370 543134
rect 103606 542898 103648 543134
rect 103328 542866 103648 542898
rect 103328 507454 103648 507486
rect 103328 507218 103370 507454
rect 103606 507218 103648 507454
rect 103328 507134 103648 507218
rect 103328 506898 103370 507134
rect 103606 506898 103648 507134
rect 103328 506866 103648 506898
rect 103328 471454 103648 471486
rect 103328 471218 103370 471454
rect 103606 471218 103648 471454
rect 103328 471134 103648 471218
rect 103328 470898 103370 471134
rect 103606 470898 103648 471134
rect 103328 470866 103648 470898
rect 103328 435454 103648 435486
rect 103328 435218 103370 435454
rect 103606 435218 103648 435454
rect 103328 435134 103648 435218
rect 103328 434898 103370 435134
rect 103606 434898 103648 435134
rect 103328 434866 103648 434898
rect 103328 399454 103648 399486
rect 103328 399218 103370 399454
rect 103606 399218 103648 399454
rect 103328 399134 103648 399218
rect 103328 398898 103370 399134
rect 103606 398898 103648 399134
rect 103328 398866 103648 398898
rect 103328 363454 103648 363486
rect 103328 363218 103370 363454
rect 103606 363218 103648 363454
rect 103328 363134 103648 363218
rect 103328 362898 103370 363134
rect 103606 362898 103648 363134
rect 103328 362866 103648 362898
rect 103328 327454 103648 327486
rect 103328 327218 103370 327454
rect 103606 327218 103648 327454
rect 103328 327134 103648 327218
rect 103328 326898 103370 327134
rect 103606 326898 103648 327134
rect 103328 326866 103648 326898
rect 103328 291454 103648 291486
rect 103328 291218 103370 291454
rect 103606 291218 103648 291454
rect 103328 291134 103648 291218
rect 103328 290898 103370 291134
rect 103606 290898 103648 291134
rect 103328 290866 103648 290898
rect 103328 255454 103648 255486
rect 103328 255218 103370 255454
rect 103606 255218 103648 255454
rect 103328 255134 103648 255218
rect 103328 254898 103370 255134
rect 103606 254898 103648 255134
rect 103328 254866 103648 254898
rect 103328 219454 103648 219486
rect 103328 219218 103370 219454
rect 103606 219218 103648 219454
rect 103328 219134 103648 219218
rect 103328 218898 103370 219134
rect 103606 218898 103648 219134
rect 103328 218866 103648 218898
rect 103328 183454 103648 183486
rect 103328 183218 103370 183454
rect 103606 183218 103648 183454
rect 103328 183134 103648 183218
rect 103328 182898 103370 183134
rect 103606 182898 103648 183134
rect 103328 182866 103648 182898
rect 103328 147454 103648 147486
rect 103328 147218 103370 147454
rect 103606 147218 103648 147454
rect 103328 147134 103648 147218
rect 103328 146898 103370 147134
rect 103606 146898 103648 147134
rect 103328 146866 103648 146898
rect 102954 104614 103574 126400
rect 106046 125629 106106 574907
rect 118688 561454 119008 561486
rect 118688 561218 118730 561454
rect 118966 561218 119008 561454
rect 118688 561134 119008 561218
rect 118688 560898 118730 561134
rect 118966 560898 119008 561134
rect 118688 560866 119008 560898
rect 149408 561454 149728 561486
rect 149408 561218 149450 561454
rect 149686 561218 149728 561454
rect 149408 561134 149728 561218
rect 149408 560898 149450 561134
rect 149686 560898 149728 561134
rect 149408 560866 149728 560898
rect 180128 561454 180448 561486
rect 180128 561218 180170 561454
rect 180406 561218 180448 561454
rect 180128 561134 180448 561218
rect 180128 560898 180170 561134
rect 180406 560898 180448 561134
rect 180128 560866 180448 560898
rect 210848 561454 211168 561486
rect 210848 561218 210890 561454
rect 211126 561218 211168 561454
rect 210848 561134 211168 561218
rect 210848 560898 210890 561134
rect 211126 560898 211168 561134
rect 210848 560866 211168 560898
rect 241568 561454 241888 561486
rect 241568 561218 241610 561454
rect 241846 561218 241888 561454
rect 241568 561134 241888 561218
rect 241568 560898 241610 561134
rect 241846 560898 241888 561134
rect 241568 560866 241888 560898
rect 272288 561454 272608 561486
rect 272288 561218 272330 561454
rect 272566 561218 272608 561454
rect 272288 561134 272608 561218
rect 272288 560898 272330 561134
rect 272566 560898 272608 561134
rect 272288 560866 272608 560898
rect 303008 561454 303328 561486
rect 303008 561218 303050 561454
rect 303286 561218 303328 561454
rect 303008 561134 303328 561218
rect 303008 560898 303050 561134
rect 303286 560898 303328 561134
rect 303008 560866 303328 560898
rect 333728 561454 334048 561486
rect 333728 561218 333770 561454
rect 334006 561218 334048 561454
rect 333728 561134 334048 561218
rect 333728 560898 333770 561134
rect 334006 560898 334048 561134
rect 333728 560866 334048 560898
rect 364448 561454 364768 561486
rect 364448 561218 364490 561454
rect 364726 561218 364768 561454
rect 364448 561134 364768 561218
rect 364448 560898 364490 561134
rect 364726 560898 364768 561134
rect 364448 560866 364768 560898
rect 395168 561454 395488 561486
rect 395168 561218 395210 561454
rect 395446 561218 395488 561454
rect 395168 561134 395488 561218
rect 395168 560898 395210 561134
rect 395446 560898 395488 561134
rect 395168 560866 395488 560898
rect 425888 561454 426208 561486
rect 425888 561218 425930 561454
rect 426166 561218 426208 561454
rect 425888 561134 426208 561218
rect 425888 560898 425930 561134
rect 426166 560898 426208 561134
rect 425888 560866 426208 560898
rect 456608 561454 456928 561486
rect 456608 561218 456650 561454
rect 456886 561218 456928 561454
rect 456608 561134 456928 561218
rect 456608 560898 456650 561134
rect 456886 560898 456928 561134
rect 456608 560866 456928 560898
rect 134048 543454 134368 543486
rect 134048 543218 134090 543454
rect 134326 543218 134368 543454
rect 134048 543134 134368 543218
rect 134048 542898 134090 543134
rect 134326 542898 134368 543134
rect 134048 542866 134368 542898
rect 164768 543454 165088 543486
rect 164768 543218 164810 543454
rect 165046 543218 165088 543454
rect 164768 543134 165088 543218
rect 164768 542898 164810 543134
rect 165046 542898 165088 543134
rect 164768 542866 165088 542898
rect 195488 543454 195808 543486
rect 195488 543218 195530 543454
rect 195766 543218 195808 543454
rect 195488 543134 195808 543218
rect 195488 542898 195530 543134
rect 195766 542898 195808 543134
rect 195488 542866 195808 542898
rect 226208 543454 226528 543486
rect 226208 543218 226250 543454
rect 226486 543218 226528 543454
rect 226208 543134 226528 543218
rect 226208 542898 226250 543134
rect 226486 542898 226528 543134
rect 226208 542866 226528 542898
rect 256928 543454 257248 543486
rect 256928 543218 256970 543454
rect 257206 543218 257248 543454
rect 256928 543134 257248 543218
rect 256928 542898 256970 543134
rect 257206 542898 257248 543134
rect 256928 542866 257248 542898
rect 287648 543454 287968 543486
rect 287648 543218 287690 543454
rect 287926 543218 287968 543454
rect 287648 543134 287968 543218
rect 287648 542898 287690 543134
rect 287926 542898 287968 543134
rect 287648 542866 287968 542898
rect 318368 543454 318688 543486
rect 318368 543218 318410 543454
rect 318646 543218 318688 543454
rect 318368 543134 318688 543218
rect 318368 542898 318410 543134
rect 318646 542898 318688 543134
rect 318368 542866 318688 542898
rect 349088 543454 349408 543486
rect 349088 543218 349130 543454
rect 349366 543218 349408 543454
rect 349088 543134 349408 543218
rect 349088 542898 349130 543134
rect 349366 542898 349408 543134
rect 349088 542866 349408 542898
rect 379808 543454 380128 543486
rect 379808 543218 379850 543454
rect 380086 543218 380128 543454
rect 379808 543134 380128 543218
rect 379808 542898 379850 543134
rect 380086 542898 380128 543134
rect 379808 542866 380128 542898
rect 410528 543454 410848 543486
rect 410528 543218 410570 543454
rect 410806 543218 410848 543454
rect 410528 543134 410848 543218
rect 410528 542898 410570 543134
rect 410806 542898 410848 543134
rect 410528 542866 410848 542898
rect 441248 543454 441568 543486
rect 441248 543218 441290 543454
rect 441526 543218 441568 543454
rect 441248 543134 441568 543218
rect 441248 542898 441290 543134
rect 441526 542898 441568 543134
rect 441248 542866 441568 542898
rect 471968 543454 472288 543486
rect 471968 543218 472010 543454
rect 472246 543218 472288 543454
rect 471968 543134 472288 543218
rect 471968 542898 472010 543134
rect 472246 542898 472288 543134
rect 471968 542866 472288 542898
rect 118688 525454 119008 525486
rect 118688 525218 118730 525454
rect 118966 525218 119008 525454
rect 118688 525134 119008 525218
rect 118688 524898 118730 525134
rect 118966 524898 119008 525134
rect 118688 524866 119008 524898
rect 149408 525454 149728 525486
rect 149408 525218 149450 525454
rect 149686 525218 149728 525454
rect 149408 525134 149728 525218
rect 149408 524898 149450 525134
rect 149686 524898 149728 525134
rect 149408 524866 149728 524898
rect 180128 525454 180448 525486
rect 180128 525218 180170 525454
rect 180406 525218 180448 525454
rect 180128 525134 180448 525218
rect 180128 524898 180170 525134
rect 180406 524898 180448 525134
rect 180128 524866 180448 524898
rect 210848 525454 211168 525486
rect 210848 525218 210890 525454
rect 211126 525218 211168 525454
rect 210848 525134 211168 525218
rect 210848 524898 210890 525134
rect 211126 524898 211168 525134
rect 210848 524866 211168 524898
rect 241568 525454 241888 525486
rect 241568 525218 241610 525454
rect 241846 525218 241888 525454
rect 241568 525134 241888 525218
rect 241568 524898 241610 525134
rect 241846 524898 241888 525134
rect 241568 524866 241888 524898
rect 272288 525454 272608 525486
rect 272288 525218 272330 525454
rect 272566 525218 272608 525454
rect 272288 525134 272608 525218
rect 272288 524898 272330 525134
rect 272566 524898 272608 525134
rect 272288 524866 272608 524898
rect 303008 525454 303328 525486
rect 303008 525218 303050 525454
rect 303286 525218 303328 525454
rect 303008 525134 303328 525218
rect 303008 524898 303050 525134
rect 303286 524898 303328 525134
rect 303008 524866 303328 524898
rect 333728 525454 334048 525486
rect 333728 525218 333770 525454
rect 334006 525218 334048 525454
rect 333728 525134 334048 525218
rect 333728 524898 333770 525134
rect 334006 524898 334048 525134
rect 333728 524866 334048 524898
rect 364448 525454 364768 525486
rect 364448 525218 364490 525454
rect 364726 525218 364768 525454
rect 364448 525134 364768 525218
rect 364448 524898 364490 525134
rect 364726 524898 364768 525134
rect 364448 524866 364768 524898
rect 395168 525454 395488 525486
rect 395168 525218 395210 525454
rect 395446 525218 395488 525454
rect 395168 525134 395488 525218
rect 395168 524898 395210 525134
rect 395446 524898 395488 525134
rect 395168 524866 395488 524898
rect 425888 525454 426208 525486
rect 425888 525218 425930 525454
rect 426166 525218 426208 525454
rect 425888 525134 426208 525218
rect 425888 524898 425930 525134
rect 426166 524898 426208 525134
rect 425888 524866 426208 524898
rect 456608 525454 456928 525486
rect 456608 525218 456650 525454
rect 456886 525218 456928 525454
rect 456608 525134 456928 525218
rect 456608 524898 456650 525134
rect 456886 524898 456928 525134
rect 456608 524866 456928 524898
rect 134048 507454 134368 507486
rect 134048 507218 134090 507454
rect 134326 507218 134368 507454
rect 134048 507134 134368 507218
rect 134048 506898 134090 507134
rect 134326 506898 134368 507134
rect 134048 506866 134368 506898
rect 164768 507454 165088 507486
rect 164768 507218 164810 507454
rect 165046 507218 165088 507454
rect 164768 507134 165088 507218
rect 164768 506898 164810 507134
rect 165046 506898 165088 507134
rect 164768 506866 165088 506898
rect 195488 507454 195808 507486
rect 195488 507218 195530 507454
rect 195766 507218 195808 507454
rect 195488 507134 195808 507218
rect 195488 506898 195530 507134
rect 195766 506898 195808 507134
rect 195488 506866 195808 506898
rect 226208 507454 226528 507486
rect 226208 507218 226250 507454
rect 226486 507218 226528 507454
rect 226208 507134 226528 507218
rect 226208 506898 226250 507134
rect 226486 506898 226528 507134
rect 226208 506866 226528 506898
rect 256928 507454 257248 507486
rect 256928 507218 256970 507454
rect 257206 507218 257248 507454
rect 256928 507134 257248 507218
rect 256928 506898 256970 507134
rect 257206 506898 257248 507134
rect 256928 506866 257248 506898
rect 287648 507454 287968 507486
rect 287648 507218 287690 507454
rect 287926 507218 287968 507454
rect 287648 507134 287968 507218
rect 287648 506898 287690 507134
rect 287926 506898 287968 507134
rect 287648 506866 287968 506898
rect 318368 507454 318688 507486
rect 318368 507218 318410 507454
rect 318646 507218 318688 507454
rect 318368 507134 318688 507218
rect 318368 506898 318410 507134
rect 318646 506898 318688 507134
rect 318368 506866 318688 506898
rect 349088 507454 349408 507486
rect 349088 507218 349130 507454
rect 349366 507218 349408 507454
rect 349088 507134 349408 507218
rect 349088 506898 349130 507134
rect 349366 506898 349408 507134
rect 349088 506866 349408 506898
rect 379808 507454 380128 507486
rect 379808 507218 379850 507454
rect 380086 507218 380128 507454
rect 379808 507134 380128 507218
rect 379808 506898 379850 507134
rect 380086 506898 380128 507134
rect 379808 506866 380128 506898
rect 410528 507454 410848 507486
rect 410528 507218 410570 507454
rect 410806 507218 410848 507454
rect 410528 507134 410848 507218
rect 410528 506898 410570 507134
rect 410806 506898 410848 507134
rect 410528 506866 410848 506898
rect 441248 507454 441568 507486
rect 441248 507218 441290 507454
rect 441526 507218 441568 507454
rect 441248 507134 441568 507218
rect 441248 506898 441290 507134
rect 441526 506898 441568 507134
rect 441248 506866 441568 506898
rect 471968 507454 472288 507486
rect 471968 507218 472010 507454
rect 472246 507218 472288 507454
rect 471968 507134 472288 507218
rect 471968 506898 472010 507134
rect 472246 506898 472288 507134
rect 471968 506866 472288 506898
rect 118688 489454 119008 489486
rect 118688 489218 118730 489454
rect 118966 489218 119008 489454
rect 118688 489134 119008 489218
rect 118688 488898 118730 489134
rect 118966 488898 119008 489134
rect 118688 488866 119008 488898
rect 149408 489454 149728 489486
rect 149408 489218 149450 489454
rect 149686 489218 149728 489454
rect 149408 489134 149728 489218
rect 149408 488898 149450 489134
rect 149686 488898 149728 489134
rect 149408 488866 149728 488898
rect 180128 489454 180448 489486
rect 180128 489218 180170 489454
rect 180406 489218 180448 489454
rect 180128 489134 180448 489218
rect 180128 488898 180170 489134
rect 180406 488898 180448 489134
rect 180128 488866 180448 488898
rect 210848 489454 211168 489486
rect 210848 489218 210890 489454
rect 211126 489218 211168 489454
rect 210848 489134 211168 489218
rect 210848 488898 210890 489134
rect 211126 488898 211168 489134
rect 210848 488866 211168 488898
rect 241568 489454 241888 489486
rect 241568 489218 241610 489454
rect 241846 489218 241888 489454
rect 241568 489134 241888 489218
rect 241568 488898 241610 489134
rect 241846 488898 241888 489134
rect 241568 488866 241888 488898
rect 272288 489454 272608 489486
rect 272288 489218 272330 489454
rect 272566 489218 272608 489454
rect 272288 489134 272608 489218
rect 272288 488898 272330 489134
rect 272566 488898 272608 489134
rect 272288 488866 272608 488898
rect 303008 489454 303328 489486
rect 303008 489218 303050 489454
rect 303286 489218 303328 489454
rect 303008 489134 303328 489218
rect 303008 488898 303050 489134
rect 303286 488898 303328 489134
rect 303008 488866 303328 488898
rect 333728 489454 334048 489486
rect 333728 489218 333770 489454
rect 334006 489218 334048 489454
rect 333728 489134 334048 489218
rect 333728 488898 333770 489134
rect 334006 488898 334048 489134
rect 333728 488866 334048 488898
rect 364448 489454 364768 489486
rect 364448 489218 364490 489454
rect 364726 489218 364768 489454
rect 364448 489134 364768 489218
rect 364448 488898 364490 489134
rect 364726 488898 364768 489134
rect 364448 488866 364768 488898
rect 395168 489454 395488 489486
rect 395168 489218 395210 489454
rect 395446 489218 395488 489454
rect 395168 489134 395488 489218
rect 395168 488898 395210 489134
rect 395446 488898 395488 489134
rect 395168 488866 395488 488898
rect 425888 489454 426208 489486
rect 425888 489218 425930 489454
rect 426166 489218 426208 489454
rect 425888 489134 426208 489218
rect 425888 488898 425930 489134
rect 426166 488898 426208 489134
rect 425888 488866 426208 488898
rect 456608 489454 456928 489486
rect 456608 489218 456650 489454
rect 456886 489218 456928 489454
rect 456608 489134 456928 489218
rect 456608 488898 456650 489134
rect 456886 488898 456928 489134
rect 456608 488866 456928 488898
rect 134048 471454 134368 471486
rect 134048 471218 134090 471454
rect 134326 471218 134368 471454
rect 134048 471134 134368 471218
rect 134048 470898 134090 471134
rect 134326 470898 134368 471134
rect 134048 470866 134368 470898
rect 164768 471454 165088 471486
rect 164768 471218 164810 471454
rect 165046 471218 165088 471454
rect 164768 471134 165088 471218
rect 164768 470898 164810 471134
rect 165046 470898 165088 471134
rect 164768 470866 165088 470898
rect 195488 471454 195808 471486
rect 195488 471218 195530 471454
rect 195766 471218 195808 471454
rect 195488 471134 195808 471218
rect 195488 470898 195530 471134
rect 195766 470898 195808 471134
rect 195488 470866 195808 470898
rect 226208 471454 226528 471486
rect 226208 471218 226250 471454
rect 226486 471218 226528 471454
rect 226208 471134 226528 471218
rect 226208 470898 226250 471134
rect 226486 470898 226528 471134
rect 226208 470866 226528 470898
rect 256928 471454 257248 471486
rect 256928 471218 256970 471454
rect 257206 471218 257248 471454
rect 256928 471134 257248 471218
rect 256928 470898 256970 471134
rect 257206 470898 257248 471134
rect 256928 470866 257248 470898
rect 287648 471454 287968 471486
rect 287648 471218 287690 471454
rect 287926 471218 287968 471454
rect 287648 471134 287968 471218
rect 287648 470898 287690 471134
rect 287926 470898 287968 471134
rect 287648 470866 287968 470898
rect 318368 471454 318688 471486
rect 318368 471218 318410 471454
rect 318646 471218 318688 471454
rect 318368 471134 318688 471218
rect 318368 470898 318410 471134
rect 318646 470898 318688 471134
rect 318368 470866 318688 470898
rect 349088 471454 349408 471486
rect 349088 471218 349130 471454
rect 349366 471218 349408 471454
rect 349088 471134 349408 471218
rect 349088 470898 349130 471134
rect 349366 470898 349408 471134
rect 349088 470866 349408 470898
rect 379808 471454 380128 471486
rect 379808 471218 379850 471454
rect 380086 471218 380128 471454
rect 379808 471134 380128 471218
rect 379808 470898 379850 471134
rect 380086 470898 380128 471134
rect 379808 470866 380128 470898
rect 410528 471454 410848 471486
rect 410528 471218 410570 471454
rect 410806 471218 410848 471454
rect 410528 471134 410848 471218
rect 410528 470898 410570 471134
rect 410806 470898 410848 471134
rect 410528 470866 410848 470898
rect 441248 471454 441568 471486
rect 441248 471218 441290 471454
rect 441526 471218 441568 471454
rect 441248 471134 441568 471218
rect 441248 470898 441290 471134
rect 441526 470898 441568 471134
rect 441248 470866 441568 470898
rect 471968 471454 472288 471486
rect 471968 471218 472010 471454
rect 472246 471218 472288 471454
rect 471968 471134 472288 471218
rect 471968 470898 472010 471134
rect 472246 470898 472288 471134
rect 471968 470866 472288 470898
rect 118688 453454 119008 453486
rect 118688 453218 118730 453454
rect 118966 453218 119008 453454
rect 118688 453134 119008 453218
rect 118688 452898 118730 453134
rect 118966 452898 119008 453134
rect 118688 452866 119008 452898
rect 149408 453454 149728 453486
rect 149408 453218 149450 453454
rect 149686 453218 149728 453454
rect 149408 453134 149728 453218
rect 149408 452898 149450 453134
rect 149686 452898 149728 453134
rect 149408 452866 149728 452898
rect 180128 453454 180448 453486
rect 180128 453218 180170 453454
rect 180406 453218 180448 453454
rect 180128 453134 180448 453218
rect 180128 452898 180170 453134
rect 180406 452898 180448 453134
rect 180128 452866 180448 452898
rect 210848 453454 211168 453486
rect 210848 453218 210890 453454
rect 211126 453218 211168 453454
rect 210848 453134 211168 453218
rect 210848 452898 210890 453134
rect 211126 452898 211168 453134
rect 210848 452866 211168 452898
rect 241568 453454 241888 453486
rect 241568 453218 241610 453454
rect 241846 453218 241888 453454
rect 241568 453134 241888 453218
rect 241568 452898 241610 453134
rect 241846 452898 241888 453134
rect 241568 452866 241888 452898
rect 272288 453454 272608 453486
rect 272288 453218 272330 453454
rect 272566 453218 272608 453454
rect 272288 453134 272608 453218
rect 272288 452898 272330 453134
rect 272566 452898 272608 453134
rect 272288 452866 272608 452898
rect 303008 453454 303328 453486
rect 303008 453218 303050 453454
rect 303286 453218 303328 453454
rect 303008 453134 303328 453218
rect 303008 452898 303050 453134
rect 303286 452898 303328 453134
rect 303008 452866 303328 452898
rect 333728 453454 334048 453486
rect 333728 453218 333770 453454
rect 334006 453218 334048 453454
rect 333728 453134 334048 453218
rect 333728 452898 333770 453134
rect 334006 452898 334048 453134
rect 333728 452866 334048 452898
rect 364448 453454 364768 453486
rect 364448 453218 364490 453454
rect 364726 453218 364768 453454
rect 364448 453134 364768 453218
rect 364448 452898 364490 453134
rect 364726 452898 364768 453134
rect 364448 452866 364768 452898
rect 395168 453454 395488 453486
rect 395168 453218 395210 453454
rect 395446 453218 395488 453454
rect 395168 453134 395488 453218
rect 395168 452898 395210 453134
rect 395446 452898 395488 453134
rect 395168 452866 395488 452898
rect 425888 453454 426208 453486
rect 425888 453218 425930 453454
rect 426166 453218 426208 453454
rect 425888 453134 426208 453218
rect 425888 452898 425930 453134
rect 426166 452898 426208 453134
rect 425888 452866 426208 452898
rect 456608 453454 456928 453486
rect 456608 453218 456650 453454
rect 456886 453218 456928 453454
rect 456608 453134 456928 453218
rect 456608 452898 456650 453134
rect 456886 452898 456928 453134
rect 456608 452866 456928 452898
rect 134048 435454 134368 435486
rect 134048 435218 134090 435454
rect 134326 435218 134368 435454
rect 134048 435134 134368 435218
rect 134048 434898 134090 435134
rect 134326 434898 134368 435134
rect 134048 434866 134368 434898
rect 164768 435454 165088 435486
rect 164768 435218 164810 435454
rect 165046 435218 165088 435454
rect 164768 435134 165088 435218
rect 164768 434898 164810 435134
rect 165046 434898 165088 435134
rect 164768 434866 165088 434898
rect 195488 435454 195808 435486
rect 195488 435218 195530 435454
rect 195766 435218 195808 435454
rect 195488 435134 195808 435218
rect 195488 434898 195530 435134
rect 195766 434898 195808 435134
rect 195488 434866 195808 434898
rect 226208 435454 226528 435486
rect 226208 435218 226250 435454
rect 226486 435218 226528 435454
rect 226208 435134 226528 435218
rect 226208 434898 226250 435134
rect 226486 434898 226528 435134
rect 226208 434866 226528 434898
rect 256928 435454 257248 435486
rect 256928 435218 256970 435454
rect 257206 435218 257248 435454
rect 256928 435134 257248 435218
rect 256928 434898 256970 435134
rect 257206 434898 257248 435134
rect 256928 434866 257248 434898
rect 287648 435454 287968 435486
rect 287648 435218 287690 435454
rect 287926 435218 287968 435454
rect 287648 435134 287968 435218
rect 287648 434898 287690 435134
rect 287926 434898 287968 435134
rect 287648 434866 287968 434898
rect 318368 435454 318688 435486
rect 318368 435218 318410 435454
rect 318646 435218 318688 435454
rect 318368 435134 318688 435218
rect 318368 434898 318410 435134
rect 318646 434898 318688 435134
rect 318368 434866 318688 434898
rect 349088 435454 349408 435486
rect 349088 435218 349130 435454
rect 349366 435218 349408 435454
rect 349088 435134 349408 435218
rect 349088 434898 349130 435134
rect 349366 434898 349408 435134
rect 349088 434866 349408 434898
rect 379808 435454 380128 435486
rect 379808 435218 379850 435454
rect 380086 435218 380128 435454
rect 379808 435134 380128 435218
rect 379808 434898 379850 435134
rect 380086 434898 380128 435134
rect 379808 434866 380128 434898
rect 410528 435454 410848 435486
rect 410528 435218 410570 435454
rect 410806 435218 410848 435454
rect 410528 435134 410848 435218
rect 410528 434898 410570 435134
rect 410806 434898 410848 435134
rect 410528 434866 410848 434898
rect 441248 435454 441568 435486
rect 441248 435218 441290 435454
rect 441526 435218 441568 435454
rect 441248 435134 441568 435218
rect 441248 434898 441290 435134
rect 441526 434898 441568 435134
rect 441248 434866 441568 434898
rect 471968 435454 472288 435486
rect 471968 435218 472010 435454
rect 472246 435218 472288 435454
rect 471968 435134 472288 435218
rect 471968 434898 472010 435134
rect 472246 434898 472288 435134
rect 471968 434866 472288 434898
rect 118688 417454 119008 417486
rect 118688 417218 118730 417454
rect 118966 417218 119008 417454
rect 118688 417134 119008 417218
rect 118688 416898 118730 417134
rect 118966 416898 119008 417134
rect 118688 416866 119008 416898
rect 149408 417454 149728 417486
rect 149408 417218 149450 417454
rect 149686 417218 149728 417454
rect 149408 417134 149728 417218
rect 149408 416898 149450 417134
rect 149686 416898 149728 417134
rect 149408 416866 149728 416898
rect 180128 417454 180448 417486
rect 180128 417218 180170 417454
rect 180406 417218 180448 417454
rect 180128 417134 180448 417218
rect 180128 416898 180170 417134
rect 180406 416898 180448 417134
rect 180128 416866 180448 416898
rect 210848 417454 211168 417486
rect 210848 417218 210890 417454
rect 211126 417218 211168 417454
rect 210848 417134 211168 417218
rect 210848 416898 210890 417134
rect 211126 416898 211168 417134
rect 210848 416866 211168 416898
rect 241568 417454 241888 417486
rect 241568 417218 241610 417454
rect 241846 417218 241888 417454
rect 241568 417134 241888 417218
rect 241568 416898 241610 417134
rect 241846 416898 241888 417134
rect 241568 416866 241888 416898
rect 272288 417454 272608 417486
rect 272288 417218 272330 417454
rect 272566 417218 272608 417454
rect 272288 417134 272608 417218
rect 272288 416898 272330 417134
rect 272566 416898 272608 417134
rect 272288 416866 272608 416898
rect 303008 417454 303328 417486
rect 303008 417218 303050 417454
rect 303286 417218 303328 417454
rect 303008 417134 303328 417218
rect 303008 416898 303050 417134
rect 303286 416898 303328 417134
rect 303008 416866 303328 416898
rect 333728 417454 334048 417486
rect 333728 417218 333770 417454
rect 334006 417218 334048 417454
rect 333728 417134 334048 417218
rect 333728 416898 333770 417134
rect 334006 416898 334048 417134
rect 333728 416866 334048 416898
rect 364448 417454 364768 417486
rect 364448 417218 364490 417454
rect 364726 417218 364768 417454
rect 364448 417134 364768 417218
rect 364448 416898 364490 417134
rect 364726 416898 364768 417134
rect 364448 416866 364768 416898
rect 395168 417454 395488 417486
rect 395168 417218 395210 417454
rect 395446 417218 395488 417454
rect 395168 417134 395488 417218
rect 395168 416898 395210 417134
rect 395446 416898 395488 417134
rect 395168 416866 395488 416898
rect 425888 417454 426208 417486
rect 425888 417218 425930 417454
rect 426166 417218 426208 417454
rect 425888 417134 426208 417218
rect 425888 416898 425930 417134
rect 426166 416898 426208 417134
rect 425888 416866 426208 416898
rect 456608 417454 456928 417486
rect 456608 417218 456650 417454
rect 456886 417218 456928 417454
rect 456608 417134 456928 417218
rect 456608 416898 456650 417134
rect 456886 416898 456928 417134
rect 456608 416866 456928 416898
rect 134048 399454 134368 399486
rect 134048 399218 134090 399454
rect 134326 399218 134368 399454
rect 134048 399134 134368 399218
rect 134048 398898 134090 399134
rect 134326 398898 134368 399134
rect 134048 398866 134368 398898
rect 164768 399454 165088 399486
rect 164768 399218 164810 399454
rect 165046 399218 165088 399454
rect 164768 399134 165088 399218
rect 164768 398898 164810 399134
rect 165046 398898 165088 399134
rect 164768 398866 165088 398898
rect 195488 399454 195808 399486
rect 195488 399218 195530 399454
rect 195766 399218 195808 399454
rect 195488 399134 195808 399218
rect 195488 398898 195530 399134
rect 195766 398898 195808 399134
rect 195488 398866 195808 398898
rect 226208 399454 226528 399486
rect 226208 399218 226250 399454
rect 226486 399218 226528 399454
rect 226208 399134 226528 399218
rect 226208 398898 226250 399134
rect 226486 398898 226528 399134
rect 226208 398866 226528 398898
rect 256928 399454 257248 399486
rect 256928 399218 256970 399454
rect 257206 399218 257248 399454
rect 256928 399134 257248 399218
rect 256928 398898 256970 399134
rect 257206 398898 257248 399134
rect 256928 398866 257248 398898
rect 287648 399454 287968 399486
rect 287648 399218 287690 399454
rect 287926 399218 287968 399454
rect 287648 399134 287968 399218
rect 287648 398898 287690 399134
rect 287926 398898 287968 399134
rect 287648 398866 287968 398898
rect 318368 399454 318688 399486
rect 318368 399218 318410 399454
rect 318646 399218 318688 399454
rect 318368 399134 318688 399218
rect 318368 398898 318410 399134
rect 318646 398898 318688 399134
rect 318368 398866 318688 398898
rect 349088 399454 349408 399486
rect 349088 399218 349130 399454
rect 349366 399218 349408 399454
rect 349088 399134 349408 399218
rect 349088 398898 349130 399134
rect 349366 398898 349408 399134
rect 349088 398866 349408 398898
rect 379808 399454 380128 399486
rect 379808 399218 379850 399454
rect 380086 399218 380128 399454
rect 379808 399134 380128 399218
rect 379808 398898 379850 399134
rect 380086 398898 380128 399134
rect 379808 398866 380128 398898
rect 410528 399454 410848 399486
rect 410528 399218 410570 399454
rect 410806 399218 410848 399454
rect 410528 399134 410848 399218
rect 410528 398898 410570 399134
rect 410806 398898 410848 399134
rect 410528 398866 410848 398898
rect 441248 399454 441568 399486
rect 441248 399218 441290 399454
rect 441526 399218 441568 399454
rect 441248 399134 441568 399218
rect 441248 398898 441290 399134
rect 441526 398898 441568 399134
rect 441248 398866 441568 398898
rect 471968 399454 472288 399486
rect 471968 399218 472010 399454
rect 472246 399218 472288 399454
rect 471968 399134 472288 399218
rect 471968 398898 472010 399134
rect 472246 398898 472288 399134
rect 471968 398866 472288 398898
rect 118688 381454 119008 381486
rect 118688 381218 118730 381454
rect 118966 381218 119008 381454
rect 118688 381134 119008 381218
rect 118688 380898 118730 381134
rect 118966 380898 119008 381134
rect 118688 380866 119008 380898
rect 149408 381454 149728 381486
rect 149408 381218 149450 381454
rect 149686 381218 149728 381454
rect 149408 381134 149728 381218
rect 149408 380898 149450 381134
rect 149686 380898 149728 381134
rect 149408 380866 149728 380898
rect 180128 381454 180448 381486
rect 180128 381218 180170 381454
rect 180406 381218 180448 381454
rect 180128 381134 180448 381218
rect 180128 380898 180170 381134
rect 180406 380898 180448 381134
rect 180128 380866 180448 380898
rect 210848 381454 211168 381486
rect 210848 381218 210890 381454
rect 211126 381218 211168 381454
rect 210848 381134 211168 381218
rect 210848 380898 210890 381134
rect 211126 380898 211168 381134
rect 210848 380866 211168 380898
rect 241568 381454 241888 381486
rect 241568 381218 241610 381454
rect 241846 381218 241888 381454
rect 241568 381134 241888 381218
rect 241568 380898 241610 381134
rect 241846 380898 241888 381134
rect 241568 380866 241888 380898
rect 272288 381454 272608 381486
rect 272288 381218 272330 381454
rect 272566 381218 272608 381454
rect 272288 381134 272608 381218
rect 272288 380898 272330 381134
rect 272566 380898 272608 381134
rect 272288 380866 272608 380898
rect 303008 381454 303328 381486
rect 303008 381218 303050 381454
rect 303286 381218 303328 381454
rect 303008 381134 303328 381218
rect 303008 380898 303050 381134
rect 303286 380898 303328 381134
rect 303008 380866 303328 380898
rect 333728 381454 334048 381486
rect 333728 381218 333770 381454
rect 334006 381218 334048 381454
rect 333728 381134 334048 381218
rect 333728 380898 333770 381134
rect 334006 380898 334048 381134
rect 333728 380866 334048 380898
rect 364448 381454 364768 381486
rect 364448 381218 364490 381454
rect 364726 381218 364768 381454
rect 364448 381134 364768 381218
rect 364448 380898 364490 381134
rect 364726 380898 364768 381134
rect 364448 380866 364768 380898
rect 395168 381454 395488 381486
rect 395168 381218 395210 381454
rect 395446 381218 395488 381454
rect 395168 381134 395488 381218
rect 395168 380898 395210 381134
rect 395446 380898 395488 381134
rect 395168 380866 395488 380898
rect 425888 381454 426208 381486
rect 425888 381218 425930 381454
rect 426166 381218 426208 381454
rect 425888 381134 426208 381218
rect 425888 380898 425930 381134
rect 426166 380898 426208 381134
rect 425888 380866 426208 380898
rect 456608 381454 456928 381486
rect 456608 381218 456650 381454
rect 456886 381218 456928 381454
rect 456608 381134 456928 381218
rect 456608 380898 456650 381134
rect 456886 380898 456928 381134
rect 456608 380866 456928 380898
rect 134048 363454 134368 363486
rect 134048 363218 134090 363454
rect 134326 363218 134368 363454
rect 134048 363134 134368 363218
rect 134048 362898 134090 363134
rect 134326 362898 134368 363134
rect 134048 362866 134368 362898
rect 164768 363454 165088 363486
rect 164768 363218 164810 363454
rect 165046 363218 165088 363454
rect 164768 363134 165088 363218
rect 164768 362898 164810 363134
rect 165046 362898 165088 363134
rect 164768 362866 165088 362898
rect 195488 363454 195808 363486
rect 195488 363218 195530 363454
rect 195766 363218 195808 363454
rect 195488 363134 195808 363218
rect 195488 362898 195530 363134
rect 195766 362898 195808 363134
rect 195488 362866 195808 362898
rect 226208 363454 226528 363486
rect 226208 363218 226250 363454
rect 226486 363218 226528 363454
rect 226208 363134 226528 363218
rect 226208 362898 226250 363134
rect 226486 362898 226528 363134
rect 226208 362866 226528 362898
rect 256928 363454 257248 363486
rect 256928 363218 256970 363454
rect 257206 363218 257248 363454
rect 256928 363134 257248 363218
rect 256928 362898 256970 363134
rect 257206 362898 257248 363134
rect 256928 362866 257248 362898
rect 287648 363454 287968 363486
rect 287648 363218 287690 363454
rect 287926 363218 287968 363454
rect 287648 363134 287968 363218
rect 287648 362898 287690 363134
rect 287926 362898 287968 363134
rect 287648 362866 287968 362898
rect 318368 363454 318688 363486
rect 318368 363218 318410 363454
rect 318646 363218 318688 363454
rect 318368 363134 318688 363218
rect 318368 362898 318410 363134
rect 318646 362898 318688 363134
rect 318368 362866 318688 362898
rect 349088 363454 349408 363486
rect 349088 363218 349130 363454
rect 349366 363218 349408 363454
rect 349088 363134 349408 363218
rect 349088 362898 349130 363134
rect 349366 362898 349408 363134
rect 349088 362866 349408 362898
rect 379808 363454 380128 363486
rect 379808 363218 379850 363454
rect 380086 363218 380128 363454
rect 379808 363134 380128 363218
rect 379808 362898 379850 363134
rect 380086 362898 380128 363134
rect 379808 362866 380128 362898
rect 410528 363454 410848 363486
rect 410528 363218 410570 363454
rect 410806 363218 410848 363454
rect 410528 363134 410848 363218
rect 410528 362898 410570 363134
rect 410806 362898 410848 363134
rect 410528 362866 410848 362898
rect 441248 363454 441568 363486
rect 441248 363218 441290 363454
rect 441526 363218 441568 363454
rect 441248 363134 441568 363218
rect 441248 362898 441290 363134
rect 441526 362898 441568 363134
rect 441248 362866 441568 362898
rect 471968 363454 472288 363486
rect 471968 363218 472010 363454
rect 472246 363218 472288 363454
rect 471968 363134 472288 363218
rect 471968 362898 472010 363134
rect 472246 362898 472288 363134
rect 471968 362866 472288 362898
rect 118688 345454 119008 345486
rect 118688 345218 118730 345454
rect 118966 345218 119008 345454
rect 118688 345134 119008 345218
rect 118688 344898 118730 345134
rect 118966 344898 119008 345134
rect 118688 344866 119008 344898
rect 149408 345454 149728 345486
rect 149408 345218 149450 345454
rect 149686 345218 149728 345454
rect 149408 345134 149728 345218
rect 149408 344898 149450 345134
rect 149686 344898 149728 345134
rect 149408 344866 149728 344898
rect 180128 345454 180448 345486
rect 180128 345218 180170 345454
rect 180406 345218 180448 345454
rect 180128 345134 180448 345218
rect 180128 344898 180170 345134
rect 180406 344898 180448 345134
rect 180128 344866 180448 344898
rect 210848 345454 211168 345486
rect 210848 345218 210890 345454
rect 211126 345218 211168 345454
rect 210848 345134 211168 345218
rect 210848 344898 210890 345134
rect 211126 344898 211168 345134
rect 210848 344866 211168 344898
rect 241568 345454 241888 345486
rect 241568 345218 241610 345454
rect 241846 345218 241888 345454
rect 241568 345134 241888 345218
rect 241568 344898 241610 345134
rect 241846 344898 241888 345134
rect 241568 344866 241888 344898
rect 272288 345454 272608 345486
rect 272288 345218 272330 345454
rect 272566 345218 272608 345454
rect 272288 345134 272608 345218
rect 272288 344898 272330 345134
rect 272566 344898 272608 345134
rect 272288 344866 272608 344898
rect 303008 345454 303328 345486
rect 303008 345218 303050 345454
rect 303286 345218 303328 345454
rect 303008 345134 303328 345218
rect 303008 344898 303050 345134
rect 303286 344898 303328 345134
rect 303008 344866 303328 344898
rect 333728 345454 334048 345486
rect 333728 345218 333770 345454
rect 334006 345218 334048 345454
rect 333728 345134 334048 345218
rect 333728 344898 333770 345134
rect 334006 344898 334048 345134
rect 333728 344866 334048 344898
rect 364448 345454 364768 345486
rect 364448 345218 364490 345454
rect 364726 345218 364768 345454
rect 364448 345134 364768 345218
rect 364448 344898 364490 345134
rect 364726 344898 364768 345134
rect 364448 344866 364768 344898
rect 395168 345454 395488 345486
rect 395168 345218 395210 345454
rect 395446 345218 395488 345454
rect 395168 345134 395488 345218
rect 395168 344898 395210 345134
rect 395446 344898 395488 345134
rect 395168 344866 395488 344898
rect 425888 345454 426208 345486
rect 425888 345218 425930 345454
rect 426166 345218 426208 345454
rect 425888 345134 426208 345218
rect 425888 344898 425930 345134
rect 426166 344898 426208 345134
rect 425888 344866 426208 344898
rect 456608 345454 456928 345486
rect 456608 345218 456650 345454
rect 456886 345218 456928 345454
rect 456608 345134 456928 345218
rect 456608 344898 456650 345134
rect 456886 344898 456928 345134
rect 456608 344866 456928 344898
rect 134048 327454 134368 327486
rect 134048 327218 134090 327454
rect 134326 327218 134368 327454
rect 134048 327134 134368 327218
rect 134048 326898 134090 327134
rect 134326 326898 134368 327134
rect 134048 326866 134368 326898
rect 164768 327454 165088 327486
rect 164768 327218 164810 327454
rect 165046 327218 165088 327454
rect 164768 327134 165088 327218
rect 164768 326898 164810 327134
rect 165046 326898 165088 327134
rect 164768 326866 165088 326898
rect 195488 327454 195808 327486
rect 195488 327218 195530 327454
rect 195766 327218 195808 327454
rect 195488 327134 195808 327218
rect 195488 326898 195530 327134
rect 195766 326898 195808 327134
rect 195488 326866 195808 326898
rect 226208 327454 226528 327486
rect 226208 327218 226250 327454
rect 226486 327218 226528 327454
rect 226208 327134 226528 327218
rect 226208 326898 226250 327134
rect 226486 326898 226528 327134
rect 226208 326866 226528 326898
rect 256928 327454 257248 327486
rect 256928 327218 256970 327454
rect 257206 327218 257248 327454
rect 256928 327134 257248 327218
rect 256928 326898 256970 327134
rect 257206 326898 257248 327134
rect 256928 326866 257248 326898
rect 287648 327454 287968 327486
rect 287648 327218 287690 327454
rect 287926 327218 287968 327454
rect 287648 327134 287968 327218
rect 287648 326898 287690 327134
rect 287926 326898 287968 327134
rect 287648 326866 287968 326898
rect 318368 327454 318688 327486
rect 318368 327218 318410 327454
rect 318646 327218 318688 327454
rect 318368 327134 318688 327218
rect 318368 326898 318410 327134
rect 318646 326898 318688 327134
rect 318368 326866 318688 326898
rect 349088 327454 349408 327486
rect 349088 327218 349130 327454
rect 349366 327218 349408 327454
rect 349088 327134 349408 327218
rect 349088 326898 349130 327134
rect 349366 326898 349408 327134
rect 349088 326866 349408 326898
rect 379808 327454 380128 327486
rect 379808 327218 379850 327454
rect 380086 327218 380128 327454
rect 379808 327134 380128 327218
rect 379808 326898 379850 327134
rect 380086 326898 380128 327134
rect 379808 326866 380128 326898
rect 410528 327454 410848 327486
rect 410528 327218 410570 327454
rect 410806 327218 410848 327454
rect 410528 327134 410848 327218
rect 410528 326898 410570 327134
rect 410806 326898 410848 327134
rect 410528 326866 410848 326898
rect 441248 327454 441568 327486
rect 441248 327218 441290 327454
rect 441526 327218 441568 327454
rect 441248 327134 441568 327218
rect 441248 326898 441290 327134
rect 441526 326898 441568 327134
rect 441248 326866 441568 326898
rect 471968 327454 472288 327486
rect 471968 327218 472010 327454
rect 472246 327218 472288 327454
rect 471968 327134 472288 327218
rect 471968 326898 472010 327134
rect 472246 326898 472288 327134
rect 471968 326866 472288 326898
rect 118688 309454 119008 309486
rect 118688 309218 118730 309454
rect 118966 309218 119008 309454
rect 118688 309134 119008 309218
rect 118688 308898 118730 309134
rect 118966 308898 119008 309134
rect 118688 308866 119008 308898
rect 149408 309454 149728 309486
rect 149408 309218 149450 309454
rect 149686 309218 149728 309454
rect 149408 309134 149728 309218
rect 149408 308898 149450 309134
rect 149686 308898 149728 309134
rect 149408 308866 149728 308898
rect 180128 309454 180448 309486
rect 180128 309218 180170 309454
rect 180406 309218 180448 309454
rect 180128 309134 180448 309218
rect 180128 308898 180170 309134
rect 180406 308898 180448 309134
rect 180128 308866 180448 308898
rect 210848 309454 211168 309486
rect 210848 309218 210890 309454
rect 211126 309218 211168 309454
rect 210848 309134 211168 309218
rect 210848 308898 210890 309134
rect 211126 308898 211168 309134
rect 210848 308866 211168 308898
rect 241568 309454 241888 309486
rect 241568 309218 241610 309454
rect 241846 309218 241888 309454
rect 241568 309134 241888 309218
rect 241568 308898 241610 309134
rect 241846 308898 241888 309134
rect 241568 308866 241888 308898
rect 272288 309454 272608 309486
rect 272288 309218 272330 309454
rect 272566 309218 272608 309454
rect 272288 309134 272608 309218
rect 272288 308898 272330 309134
rect 272566 308898 272608 309134
rect 272288 308866 272608 308898
rect 303008 309454 303328 309486
rect 303008 309218 303050 309454
rect 303286 309218 303328 309454
rect 303008 309134 303328 309218
rect 303008 308898 303050 309134
rect 303286 308898 303328 309134
rect 303008 308866 303328 308898
rect 333728 309454 334048 309486
rect 333728 309218 333770 309454
rect 334006 309218 334048 309454
rect 333728 309134 334048 309218
rect 333728 308898 333770 309134
rect 334006 308898 334048 309134
rect 333728 308866 334048 308898
rect 364448 309454 364768 309486
rect 364448 309218 364490 309454
rect 364726 309218 364768 309454
rect 364448 309134 364768 309218
rect 364448 308898 364490 309134
rect 364726 308898 364768 309134
rect 364448 308866 364768 308898
rect 395168 309454 395488 309486
rect 395168 309218 395210 309454
rect 395446 309218 395488 309454
rect 395168 309134 395488 309218
rect 395168 308898 395210 309134
rect 395446 308898 395488 309134
rect 395168 308866 395488 308898
rect 425888 309454 426208 309486
rect 425888 309218 425930 309454
rect 426166 309218 426208 309454
rect 425888 309134 426208 309218
rect 425888 308898 425930 309134
rect 426166 308898 426208 309134
rect 425888 308866 426208 308898
rect 456608 309454 456928 309486
rect 456608 309218 456650 309454
rect 456886 309218 456928 309454
rect 456608 309134 456928 309218
rect 456608 308898 456650 309134
rect 456886 308898 456928 309134
rect 456608 308866 456928 308898
rect 134048 291454 134368 291486
rect 134048 291218 134090 291454
rect 134326 291218 134368 291454
rect 134048 291134 134368 291218
rect 134048 290898 134090 291134
rect 134326 290898 134368 291134
rect 134048 290866 134368 290898
rect 164768 291454 165088 291486
rect 164768 291218 164810 291454
rect 165046 291218 165088 291454
rect 164768 291134 165088 291218
rect 164768 290898 164810 291134
rect 165046 290898 165088 291134
rect 164768 290866 165088 290898
rect 195488 291454 195808 291486
rect 195488 291218 195530 291454
rect 195766 291218 195808 291454
rect 195488 291134 195808 291218
rect 195488 290898 195530 291134
rect 195766 290898 195808 291134
rect 195488 290866 195808 290898
rect 226208 291454 226528 291486
rect 226208 291218 226250 291454
rect 226486 291218 226528 291454
rect 226208 291134 226528 291218
rect 226208 290898 226250 291134
rect 226486 290898 226528 291134
rect 226208 290866 226528 290898
rect 256928 291454 257248 291486
rect 256928 291218 256970 291454
rect 257206 291218 257248 291454
rect 256928 291134 257248 291218
rect 256928 290898 256970 291134
rect 257206 290898 257248 291134
rect 256928 290866 257248 290898
rect 287648 291454 287968 291486
rect 287648 291218 287690 291454
rect 287926 291218 287968 291454
rect 287648 291134 287968 291218
rect 287648 290898 287690 291134
rect 287926 290898 287968 291134
rect 287648 290866 287968 290898
rect 318368 291454 318688 291486
rect 318368 291218 318410 291454
rect 318646 291218 318688 291454
rect 318368 291134 318688 291218
rect 318368 290898 318410 291134
rect 318646 290898 318688 291134
rect 318368 290866 318688 290898
rect 349088 291454 349408 291486
rect 349088 291218 349130 291454
rect 349366 291218 349408 291454
rect 349088 291134 349408 291218
rect 349088 290898 349130 291134
rect 349366 290898 349408 291134
rect 349088 290866 349408 290898
rect 379808 291454 380128 291486
rect 379808 291218 379850 291454
rect 380086 291218 380128 291454
rect 379808 291134 380128 291218
rect 379808 290898 379850 291134
rect 380086 290898 380128 291134
rect 379808 290866 380128 290898
rect 410528 291454 410848 291486
rect 410528 291218 410570 291454
rect 410806 291218 410848 291454
rect 410528 291134 410848 291218
rect 410528 290898 410570 291134
rect 410806 290898 410848 291134
rect 410528 290866 410848 290898
rect 441248 291454 441568 291486
rect 441248 291218 441290 291454
rect 441526 291218 441568 291454
rect 441248 291134 441568 291218
rect 441248 290898 441290 291134
rect 441526 290898 441568 291134
rect 441248 290866 441568 290898
rect 471968 291454 472288 291486
rect 471968 291218 472010 291454
rect 472246 291218 472288 291454
rect 471968 291134 472288 291218
rect 471968 290898 472010 291134
rect 472246 290898 472288 291134
rect 471968 290866 472288 290898
rect 118688 273454 119008 273486
rect 118688 273218 118730 273454
rect 118966 273218 119008 273454
rect 118688 273134 119008 273218
rect 118688 272898 118730 273134
rect 118966 272898 119008 273134
rect 118688 272866 119008 272898
rect 149408 273454 149728 273486
rect 149408 273218 149450 273454
rect 149686 273218 149728 273454
rect 149408 273134 149728 273218
rect 149408 272898 149450 273134
rect 149686 272898 149728 273134
rect 149408 272866 149728 272898
rect 180128 273454 180448 273486
rect 180128 273218 180170 273454
rect 180406 273218 180448 273454
rect 180128 273134 180448 273218
rect 180128 272898 180170 273134
rect 180406 272898 180448 273134
rect 180128 272866 180448 272898
rect 210848 273454 211168 273486
rect 210848 273218 210890 273454
rect 211126 273218 211168 273454
rect 210848 273134 211168 273218
rect 210848 272898 210890 273134
rect 211126 272898 211168 273134
rect 210848 272866 211168 272898
rect 241568 273454 241888 273486
rect 241568 273218 241610 273454
rect 241846 273218 241888 273454
rect 241568 273134 241888 273218
rect 241568 272898 241610 273134
rect 241846 272898 241888 273134
rect 241568 272866 241888 272898
rect 272288 273454 272608 273486
rect 272288 273218 272330 273454
rect 272566 273218 272608 273454
rect 272288 273134 272608 273218
rect 272288 272898 272330 273134
rect 272566 272898 272608 273134
rect 272288 272866 272608 272898
rect 303008 273454 303328 273486
rect 303008 273218 303050 273454
rect 303286 273218 303328 273454
rect 303008 273134 303328 273218
rect 303008 272898 303050 273134
rect 303286 272898 303328 273134
rect 303008 272866 303328 272898
rect 333728 273454 334048 273486
rect 333728 273218 333770 273454
rect 334006 273218 334048 273454
rect 333728 273134 334048 273218
rect 333728 272898 333770 273134
rect 334006 272898 334048 273134
rect 333728 272866 334048 272898
rect 364448 273454 364768 273486
rect 364448 273218 364490 273454
rect 364726 273218 364768 273454
rect 364448 273134 364768 273218
rect 364448 272898 364490 273134
rect 364726 272898 364768 273134
rect 364448 272866 364768 272898
rect 395168 273454 395488 273486
rect 395168 273218 395210 273454
rect 395446 273218 395488 273454
rect 395168 273134 395488 273218
rect 395168 272898 395210 273134
rect 395446 272898 395488 273134
rect 395168 272866 395488 272898
rect 425888 273454 426208 273486
rect 425888 273218 425930 273454
rect 426166 273218 426208 273454
rect 425888 273134 426208 273218
rect 425888 272898 425930 273134
rect 426166 272898 426208 273134
rect 425888 272866 426208 272898
rect 456608 273454 456928 273486
rect 456608 273218 456650 273454
rect 456886 273218 456928 273454
rect 456608 273134 456928 273218
rect 456608 272898 456650 273134
rect 456886 272898 456928 273134
rect 456608 272866 456928 272898
rect 134048 255454 134368 255486
rect 134048 255218 134090 255454
rect 134326 255218 134368 255454
rect 134048 255134 134368 255218
rect 134048 254898 134090 255134
rect 134326 254898 134368 255134
rect 134048 254866 134368 254898
rect 164768 255454 165088 255486
rect 164768 255218 164810 255454
rect 165046 255218 165088 255454
rect 164768 255134 165088 255218
rect 164768 254898 164810 255134
rect 165046 254898 165088 255134
rect 164768 254866 165088 254898
rect 195488 255454 195808 255486
rect 195488 255218 195530 255454
rect 195766 255218 195808 255454
rect 195488 255134 195808 255218
rect 195488 254898 195530 255134
rect 195766 254898 195808 255134
rect 195488 254866 195808 254898
rect 226208 255454 226528 255486
rect 226208 255218 226250 255454
rect 226486 255218 226528 255454
rect 226208 255134 226528 255218
rect 226208 254898 226250 255134
rect 226486 254898 226528 255134
rect 226208 254866 226528 254898
rect 256928 255454 257248 255486
rect 256928 255218 256970 255454
rect 257206 255218 257248 255454
rect 256928 255134 257248 255218
rect 256928 254898 256970 255134
rect 257206 254898 257248 255134
rect 256928 254866 257248 254898
rect 287648 255454 287968 255486
rect 287648 255218 287690 255454
rect 287926 255218 287968 255454
rect 287648 255134 287968 255218
rect 287648 254898 287690 255134
rect 287926 254898 287968 255134
rect 287648 254866 287968 254898
rect 318368 255454 318688 255486
rect 318368 255218 318410 255454
rect 318646 255218 318688 255454
rect 318368 255134 318688 255218
rect 318368 254898 318410 255134
rect 318646 254898 318688 255134
rect 318368 254866 318688 254898
rect 349088 255454 349408 255486
rect 349088 255218 349130 255454
rect 349366 255218 349408 255454
rect 349088 255134 349408 255218
rect 349088 254898 349130 255134
rect 349366 254898 349408 255134
rect 349088 254866 349408 254898
rect 379808 255454 380128 255486
rect 379808 255218 379850 255454
rect 380086 255218 380128 255454
rect 379808 255134 380128 255218
rect 379808 254898 379850 255134
rect 380086 254898 380128 255134
rect 379808 254866 380128 254898
rect 410528 255454 410848 255486
rect 410528 255218 410570 255454
rect 410806 255218 410848 255454
rect 410528 255134 410848 255218
rect 410528 254898 410570 255134
rect 410806 254898 410848 255134
rect 410528 254866 410848 254898
rect 441248 255454 441568 255486
rect 441248 255218 441290 255454
rect 441526 255218 441568 255454
rect 441248 255134 441568 255218
rect 441248 254898 441290 255134
rect 441526 254898 441568 255134
rect 441248 254866 441568 254898
rect 471968 255454 472288 255486
rect 471968 255218 472010 255454
rect 472246 255218 472288 255454
rect 471968 255134 472288 255218
rect 471968 254898 472010 255134
rect 472246 254898 472288 255134
rect 471968 254866 472288 254898
rect 118688 237454 119008 237486
rect 118688 237218 118730 237454
rect 118966 237218 119008 237454
rect 118688 237134 119008 237218
rect 118688 236898 118730 237134
rect 118966 236898 119008 237134
rect 118688 236866 119008 236898
rect 149408 237454 149728 237486
rect 149408 237218 149450 237454
rect 149686 237218 149728 237454
rect 149408 237134 149728 237218
rect 149408 236898 149450 237134
rect 149686 236898 149728 237134
rect 149408 236866 149728 236898
rect 180128 237454 180448 237486
rect 180128 237218 180170 237454
rect 180406 237218 180448 237454
rect 180128 237134 180448 237218
rect 180128 236898 180170 237134
rect 180406 236898 180448 237134
rect 180128 236866 180448 236898
rect 210848 237454 211168 237486
rect 210848 237218 210890 237454
rect 211126 237218 211168 237454
rect 210848 237134 211168 237218
rect 210848 236898 210890 237134
rect 211126 236898 211168 237134
rect 210848 236866 211168 236898
rect 241568 237454 241888 237486
rect 241568 237218 241610 237454
rect 241846 237218 241888 237454
rect 241568 237134 241888 237218
rect 241568 236898 241610 237134
rect 241846 236898 241888 237134
rect 241568 236866 241888 236898
rect 272288 237454 272608 237486
rect 272288 237218 272330 237454
rect 272566 237218 272608 237454
rect 272288 237134 272608 237218
rect 272288 236898 272330 237134
rect 272566 236898 272608 237134
rect 272288 236866 272608 236898
rect 303008 237454 303328 237486
rect 303008 237218 303050 237454
rect 303286 237218 303328 237454
rect 303008 237134 303328 237218
rect 303008 236898 303050 237134
rect 303286 236898 303328 237134
rect 303008 236866 303328 236898
rect 333728 237454 334048 237486
rect 333728 237218 333770 237454
rect 334006 237218 334048 237454
rect 333728 237134 334048 237218
rect 333728 236898 333770 237134
rect 334006 236898 334048 237134
rect 333728 236866 334048 236898
rect 364448 237454 364768 237486
rect 364448 237218 364490 237454
rect 364726 237218 364768 237454
rect 364448 237134 364768 237218
rect 364448 236898 364490 237134
rect 364726 236898 364768 237134
rect 364448 236866 364768 236898
rect 395168 237454 395488 237486
rect 395168 237218 395210 237454
rect 395446 237218 395488 237454
rect 395168 237134 395488 237218
rect 395168 236898 395210 237134
rect 395446 236898 395488 237134
rect 395168 236866 395488 236898
rect 425888 237454 426208 237486
rect 425888 237218 425930 237454
rect 426166 237218 426208 237454
rect 425888 237134 426208 237218
rect 425888 236898 425930 237134
rect 426166 236898 426208 237134
rect 425888 236866 426208 236898
rect 456608 237454 456928 237486
rect 456608 237218 456650 237454
rect 456886 237218 456928 237454
rect 456608 237134 456928 237218
rect 456608 236898 456650 237134
rect 456886 236898 456928 237134
rect 456608 236866 456928 236898
rect 134048 219454 134368 219486
rect 134048 219218 134090 219454
rect 134326 219218 134368 219454
rect 134048 219134 134368 219218
rect 134048 218898 134090 219134
rect 134326 218898 134368 219134
rect 134048 218866 134368 218898
rect 164768 219454 165088 219486
rect 164768 219218 164810 219454
rect 165046 219218 165088 219454
rect 164768 219134 165088 219218
rect 164768 218898 164810 219134
rect 165046 218898 165088 219134
rect 164768 218866 165088 218898
rect 195488 219454 195808 219486
rect 195488 219218 195530 219454
rect 195766 219218 195808 219454
rect 195488 219134 195808 219218
rect 195488 218898 195530 219134
rect 195766 218898 195808 219134
rect 195488 218866 195808 218898
rect 226208 219454 226528 219486
rect 226208 219218 226250 219454
rect 226486 219218 226528 219454
rect 226208 219134 226528 219218
rect 226208 218898 226250 219134
rect 226486 218898 226528 219134
rect 226208 218866 226528 218898
rect 256928 219454 257248 219486
rect 256928 219218 256970 219454
rect 257206 219218 257248 219454
rect 256928 219134 257248 219218
rect 256928 218898 256970 219134
rect 257206 218898 257248 219134
rect 256928 218866 257248 218898
rect 287648 219454 287968 219486
rect 287648 219218 287690 219454
rect 287926 219218 287968 219454
rect 287648 219134 287968 219218
rect 287648 218898 287690 219134
rect 287926 218898 287968 219134
rect 287648 218866 287968 218898
rect 318368 219454 318688 219486
rect 318368 219218 318410 219454
rect 318646 219218 318688 219454
rect 318368 219134 318688 219218
rect 318368 218898 318410 219134
rect 318646 218898 318688 219134
rect 318368 218866 318688 218898
rect 349088 219454 349408 219486
rect 349088 219218 349130 219454
rect 349366 219218 349408 219454
rect 349088 219134 349408 219218
rect 349088 218898 349130 219134
rect 349366 218898 349408 219134
rect 349088 218866 349408 218898
rect 379808 219454 380128 219486
rect 379808 219218 379850 219454
rect 380086 219218 380128 219454
rect 379808 219134 380128 219218
rect 379808 218898 379850 219134
rect 380086 218898 380128 219134
rect 379808 218866 380128 218898
rect 410528 219454 410848 219486
rect 410528 219218 410570 219454
rect 410806 219218 410848 219454
rect 410528 219134 410848 219218
rect 410528 218898 410570 219134
rect 410806 218898 410848 219134
rect 410528 218866 410848 218898
rect 441248 219454 441568 219486
rect 441248 219218 441290 219454
rect 441526 219218 441568 219454
rect 441248 219134 441568 219218
rect 441248 218898 441290 219134
rect 441526 218898 441568 219134
rect 441248 218866 441568 218898
rect 471968 219454 472288 219486
rect 471968 219218 472010 219454
rect 472246 219218 472288 219454
rect 471968 219134 472288 219218
rect 471968 218898 472010 219134
rect 472246 218898 472288 219134
rect 471968 218866 472288 218898
rect 118688 201454 119008 201486
rect 118688 201218 118730 201454
rect 118966 201218 119008 201454
rect 118688 201134 119008 201218
rect 118688 200898 118730 201134
rect 118966 200898 119008 201134
rect 118688 200866 119008 200898
rect 149408 201454 149728 201486
rect 149408 201218 149450 201454
rect 149686 201218 149728 201454
rect 149408 201134 149728 201218
rect 149408 200898 149450 201134
rect 149686 200898 149728 201134
rect 149408 200866 149728 200898
rect 180128 201454 180448 201486
rect 180128 201218 180170 201454
rect 180406 201218 180448 201454
rect 180128 201134 180448 201218
rect 180128 200898 180170 201134
rect 180406 200898 180448 201134
rect 180128 200866 180448 200898
rect 210848 201454 211168 201486
rect 210848 201218 210890 201454
rect 211126 201218 211168 201454
rect 210848 201134 211168 201218
rect 210848 200898 210890 201134
rect 211126 200898 211168 201134
rect 210848 200866 211168 200898
rect 241568 201454 241888 201486
rect 241568 201218 241610 201454
rect 241846 201218 241888 201454
rect 241568 201134 241888 201218
rect 241568 200898 241610 201134
rect 241846 200898 241888 201134
rect 241568 200866 241888 200898
rect 272288 201454 272608 201486
rect 272288 201218 272330 201454
rect 272566 201218 272608 201454
rect 272288 201134 272608 201218
rect 272288 200898 272330 201134
rect 272566 200898 272608 201134
rect 272288 200866 272608 200898
rect 303008 201454 303328 201486
rect 303008 201218 303050 201454
rect 303286 201218 303328 201454
rect 303008 201134 303328 201218
rect 303008 200898 303050 201134
rect 303286 200898 303328 201134
rect 303008 200866 303328 200898
rect 333728 201454 334048 201486
rect 333728 201218 333770 201454
rect 334006 201218 334048 201454
rect 333728 201134 334048 201218
rect 333728 200898 333770 201134
rect 334006 200898 334048 201134
rect 333728 200866 334048 200898
rect 364448 201454 364768 201486
rect 364448 201218 364490 201454
rect 364726 201218 364768 201454
rect 364448 201134 364768 201218
rect 364448 200898 364490 201134
rect 364726 200898 364768 201134
rect 364448 200866 364768 200898
rect 395168 201454 395488 201486
rect 395168 201218 395210 201454
rect 395446 201218 395488 201454
rect 395168 201134 395488 201218
rect 395168 200898 395210 201134
rect 395446 200898 395488 201134
rect 395168 200866 395488 200898
rect 425888 201454 426208 201486
rect 425888 201218 425930 201454
rect 426166 201218 426208 201454
rect 425888 201134 426208 201218
rect 425888 200898 425930 201134
rect 426166 200898 426208 201134
rect 425888 200866 426208 200898
rect 456608 201454 456928 201486
rect 456608 201218 456650 201454
rect 456886 201218 456928 201454
rect 456608 201134 456928 201218
rect 456608 200898 456650 201134
rect 456886 200898 456928 201134
rect 456608 200866 456928 200898
rect 134048 183454 134368 183486
rect 134048 183218 134090 183454
rect 134326 183218 134368 183454
rect 134048 183134 134368 183218
rect 134048 182898 134090 183134
rect 134326 182898 134368 183134
rect 134048 182866 134368 182898
rect 164768 183454 165088 183486
rect 164768 183218 164810 183454
rect 165046 183218 165088 183454
rect 164768 183134 165088 183218
rect 164768 182898 164810 183134
rect 165046 182898 165088 183134
rect 164768 182866 165088 182898
rect 195488 183454 195808 183486
rect 195488 183218 195530 183454
rect 195766 183218 195808 183454
rect 195488 183134 195808 183218
rect 195488 182898 195530 183134
rect 195766 182898 195808 183134
rect 195488 182866 195808 182898
rect 226208 183454 226528 183486
rect 226208 183218 226250 183454
rect 226486 183218 226528 183454
rect 226208 183134 226528 183218
rect 226208 182898 226250 183134
rect 226486 182898 226528 183134
rect 226208 182866 226528 182898
rect 256928 183454 257248 183486
rect 256928 183218 256970 183454
rect 257206 183218 257248 183454
rect 256928 183134 257248 183218
rect 256928 182898 256970 183134
rect 257206 182898 257248 183134
rect 256928 182866 257248 182898
rect 287648 183454 287968 183486
rect 287648 183218 287690 183454
rect 287926 183218 287968 183454
rect 287648 183134 287968 183218
rect 287648 182898 287690 183134
rect 287926 182898 287968 183134
rect 287648 182866 287968 182898
rect 318368 183454 318688 183486
rect 318368 183218 318410 183454
rect 318646 183218 318688 183454
rect 318368 183134 318688 183218
rect 318368 182898 318410 183134
rect 318646 182898 318688 183134
rect 318368 182866 318688 182898
rect 349088 183454 349408 183486
rect 349088 183218 349130 183454
rect 349366 183218 349408 183454
rect 349088 183134 349408 183218
rect 349088 182898 349130 183134
rect 349366 182898 349408 183134
rect 349088 182866 349408 182898
rect 379808 183454 380128 183486
rect 379808 183218 379850 183454
rect 380086 183218 380128 183454
rect 379808 183134 380128 183218
rect 379808 182898 379850 183134
rect 380086 182898 380128 183134
rect 379808 182866 380128 182898
rect 410528 183454 410848 183486
rect 410528 183218 410570 183454
rect 410806 183218 410848 183454
rect 410528 183134 410848 183218
rect 410528 182898 410570 183134
rect 410806 182898 410848 183134
rect 410528 182866 410848 182898
rect 441248 183454 441568 183486
rect 441248 183218 441290 183454
rect 441526 183218 441568 183454
rect 441248 183134 441568 183218
rect 441248 182898 441290 183134
rect 441526 182898 441568 183134
rect 441248 182866 441568 182898
rect 471968 183454 472288 183486
rect 471968 183218 472010 183454
rect 472246 183218 472288 183454
rect 471968 183134 472288 183218
rect 471968 182898 472010 183134
rect 472246 182898 472288 183134
rect 471968 182866 472288 182898
rect 118688 165454 119008 165486
rect 118688 165218 118730 165454
rect 118966 165218 119008 165454
rect 118688 165134 119008 165218
rect 118688 164898 118730 165134
rect 118966 164898 119008 165134
rect 118688 164866 119008 164898
rect 149408 165454 149728 165486
rect 149408 165218 149450 165454
rect 149686 165218 149728 165454
rect 149408 165134 149728 165218
rect 149408 164898 149450 165134
rect 149686 164898 149728 165134
rect 149408 164866 149728 164898
rect 180128 165454 180448 165486
rect 180128 165218 180170 165454
rect 180406 165218 180448 165454
rect 180128 165134 180448 165218
rect 180128 164898 180170 165134
rect 180406 164898 180448 165134
rect 180128 164866 180448 164898
rect 210848 165454 211168 165486
rect 210848 165218 210890 165454
rect 211126 165218 211168 165454
rect 210848 165134 211168 165218
rect 210848 164898 210890 165134
rect 211126 164898 211168 165134
rect 210848 164866 211168 164898
rect 241568 165454 241888 165486
rect 241568 165218 241610 165454
rect 241846 165218 241888 165454
rect 241568 165134 241888 165218
rect 241568 164898 241610 165134
rect 241846 164898 241888 165134
rect 241568 164866 241888 164898
rect 272288 165454 272608 165486
rect 272288 165218 272330 165454
rect 272566 165218 272608 165454
rect 272288 165134 272608 165218
rect 272288 164898 272330 165134
rect 272566 164898 272608 165134
rect 272288 164866 272608 164898
rect 303008 165454 303328 165486
rect 303008 165218 303050 165454
rect 303286 165218 303328 165454
rect 303008 165134 303328 165218
rect 303008 164898 303050 165134
rect 303286 164898 303328 165134
rect 303008 164866 303328 164898
rect 333728 165454 334048 165486
rect 333728 165218 333770 165454
rect 334006 165218 334048 165454
rect 333728 165134 334048 165218
rect 333728 164898 333770 165134
rect 334006 164898 334048 165134
rect 333728 164866 334048 164898
rect 364448 165454 364768 165486
rect 364448 165218 364490 165454
rect 364726 165218 364768 165454
rect 364448 165134 364768 165218
rect 364448 164898 364490 165134
rect 364726 164898 364768 165134
rect 364448 164866 364768 164898
rect 395168 165454 395488 165486
rect 395168 165218 395210 165454
rect 395446 165218 395488 165454
rect 395168 165134 395488 165218
rect 395168 164898 395210 165134
rect 395446 164898 395488 165134
rect 395168 164866 395488 164898
rect 425888 165454 426208 165486
rect 425888 165218 425930 165454
rect 426166 165218 426208 165454
rect 425888 165134 426208 165218
rect 425888 164898 425930 165134
rect 426166 164898 426208 165134
rect 425888 164866 426208 164898
rect 456608 165454 456928 165486
rect 456608 165218 456650 165454
rect 456886 165218 456928 165454
rect 456608 165134 456928 165218
rect 456608 164898 456650 165134
rect 456886 164898 456928 165134
rect 456608 164866 456928 164898
rect 134048 147454 134368 147486
rect 134048 147218 134090 147454
rect 134326 147218 134368 147454
rect 134048 147134 134368 147218
rect 134048 146898 134090 147134
rect 134326 146898 134368 147134
rect 134048 146866 134368 146898
rect 164768 147454 165088 147486
rect 164768 147218 164810 147454
rect 165046 147218 165088 147454
rect 164768 147134 165088 147218
rect 164768 146898 164810 147134
rect 165046 146898 165088 147134
rect 164768 146866 165088 146898
rect 195488 147454 195808 147486
rect 195488 147218 195530 147454
rect 195766 147218 195808 147454
rect 195488 147134 195808 147218
rect 195488 146898 195530 147134
rect 195766 146898 195808 147134
rect 195488 146866 195808 146898
rect 226208 147454 226528 147486
rect 226208 147218 226250 147454
rect 226486 147218 226528 147454
rect 226208 147134 226528 147218
rect 226208 146898 226250 147134
rect 226486 146898 226528 147134
rect 226208 146866 226528 146898
rect 256928 147454 257248 147486
rect 256928 147218 256970 147454
rect 257206 147218 257248 147454
rect 256928 147134 257248 147218
rect 256928 146898 256970 147134
rect 257206 146898 257248 147134
rect 256928 146866 257248 146898
rect 287648 147454 287968 147486
rect 287648 147218 287690 147454
rect 287926 147218 287968 147454
rect 287648 147134 287968 147218
rect 287648 146898 287690 147134
rect 287926 146898 287968 147134
rect 287648 146866 287968 146898
rect 318368 147454 318688 147486
rect 318368 147218 318410 147454
rect 318646 147218 318688 147454
rect 318368 147134 318688 147218
rect 318368 146898 318410 147134
rect 318646 146898 318688 147134
rect 318368 146866 318688 146898
rect 349088 147454 349408 147486
rect 349088 147218 349130 147454
rect 349366 147218 349408 147454
rect 349088 147134 349408 147218
rect 349088 146898 349130 147134
rect 349366 146898 349408 147134
rect 349088 146866 349408 146898
rect 379808 147454 380128 147486
rect 379808 147218 379850 147454
rect 380086 147218 380128 147454
rect 379808 147134 380128 147218
rect 379808 146898 379850 147134
rect 380086 146898 380128 147134
rect 379808 146866 380128 146898
rect 410528 147454 410848 147486
rect 410528 147218 410570 147454
rect 410806 147218 410848 147454
rect 410528 147134 410848 147218
rect 410528 146898 410570 147134
rect 410806 146898 410848 147134
rect 410528 146866 410848 146898
rect 441248 147454 441568 147486
rect 441248 147218 441290 147454
rect 441526 147218 441568 147454
rect 441248 147134 441568 147218
rect 441248 146898 441290 147134
rect 441526 146898 441568 147134
rect 441248 146866 441568 146898
rect 471968 147454 472288 147486
rect 471968 147218 472010 147454
rect 472246 147218 472288 147454
rect 471968 147134 472288 147218
rect 471968 146898 472010 147134
rect 472246 146898 472288 147134
rect 471968 146866 472288 146898
rect 106043 125628 106109 125629
rect 106043 125564 106044 125628
rect 106108 125564 106109 125628
rect 106043 125563 106109 125564
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 101995 99516 102061 99517
rect 101995 99452 101996 99516
rect 102060 99452 102061 99516
rect 101995 99451 102061 99452
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 111454 110414 126400
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 115174 114134 126400
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 118894 117854 126400
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 122614 121574 126400
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 93454 128414 126400
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 97174 132134 126400
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 100894 135854 126400
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 104614 139574 126400
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 111454 146414 126400
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 115174 150134 126400
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 118894 153854 126400
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 122614 157574 126400
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 93454 164414 126400
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 97174 168134 126400
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 100894 171854 126400
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 104614 175574 126400
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 111454 182414 126400
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 115174 186134 126400
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 118894 189854 126400
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 122614 193574 126400
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 126400
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 97174 204134 126400
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 100894 207854 126400
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 104614 211574 126400
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 111454 218414 126400
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 115174 222134 126400
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 118894 225854 126400
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 122614 229574 126400
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 126400
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 126400
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 100894 243854 126400
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 104614 247574 126400
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 111454 254414 126400
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 115174 258134 126400
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 118894 261854 126400
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 122614 265574 126400
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 93454 272414 126400
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 97174 276134 126400
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 100894 279854 126400
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 104614 283574 126400
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 111454 290414 126400
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 115174 294134 126400
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 118894 297854 126400
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 122614 301574 126400
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 93454 308414 126400
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 97174 312134 126400
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 100894 315854 126400
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 104614 319574 126400
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 111454 326414 126400
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 115174 330134 126400
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 118894 333854 126400
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 122614 337574 126400
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 93454 344414 126400
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 97174 348134 126400
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 100894 351854 126400
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 104614 355574 126400
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 111454 362414 126400
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 115174 366134 126400
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 118894 369854 126400
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 122614 373574 126400
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 93454 380414 126400
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 97174 384134 126400
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 100894 387854 126400
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 104614 391574 126400
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 111454 398414 126400
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 115174 402134 126400
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 118894 405854 126400
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 122614 409574 126400
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 93454 416414 126400
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 97174 420134 126400
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 100894 423854 126400
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 104614 427574 126400
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 111454 434414 126400
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 115174 438134 126400
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 118894 441854 126400
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 122614 445574 126400
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 93454 452414 126400
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 97174 456134 126400
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 100894 459854 126400
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 104614 463574 126400
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 111454 470414 126400
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 115174 474134 126400
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 118894 477854 126400
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 122614 481574 126400
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 481774 111757 481834 574907
rect 481771 111756 481837 111757
rect 481771 111692 481772 111756
rect 481836 111692 481837 111756
rect 481771 111691 481837 111692
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 485822 85509 485882 574907
rect 487328 561454 487648 561486
rect 487328 561218 487370 561454
rect 487606 561218 487648 561454
rect 487328 561134 487648 561218
rect 487328 560898 487370 561134
rect 487606 560898 487648 561134
rect 487328 560866 487648 560898
rect 487328 525454 487648 525486
rect 487328 525218 487370 525454
rect 487606 525218 487648 525454
rect 487328 525134 487648 525218
rect 487328 524898 487370 525134
rect 487606 524898 487648 525134
rect 487328 524866 487648 524898
rect 487328 489454 487648 489486
rect 487328 489218 487370 489454
rect 487606 489218 487648 489454
rect 487328 489134 487648 489218
rect 487328 488898 487370 489134
rect 487606 488898 487648 489134
rect 487328 488866 487648 488898
rect 487328 453454 487648 453486
rect 487328 453218 487370 453454
rect 487606 453218 487648 453454
rect 487328 453134 487648 453218
rect 487328 452898 487370 453134
rect 487606 452898 487648 453134
rect 487328 452866 487648 452898
rect 487328 417454 487648 417486
rect 487328 417218 487370 417454
rect 487606 417218 487648 417454
rect 487328 417134 487648 417218
rect 487328 416898 487370 417134
rect 487606 416898 487648 417134
rect 487328 416866 487648 416898
rect 487328 381454 487648 381486
rect 487328 381218 487370 381454
rect 487606 381218 487648 381454
rect 487328 381134 487648 381218
rect 487328 380898 487370 381134
rect 487606 380898 487648 381134
rect 487328 380866 487648 380898
rect 487328 345454 487648 345486
rect 487328 345218 487370 345454
rect 487606 345218 487648 345454
rect 487328 345134 487648 345218
rect 487328 344898 487370 345134
rect 487606 344898 487648 345134
rect 487328 344866 487648 344898
rect 487328 309454 487648 309486
rect 487328 309218 487370 309454
rect 487606 309218 487648 309454
rect 487328 309134 487648 309218
rect 487328 308898 487370 309134
rect 487606 308898 487648 309134
rect 487328 308866 487648 308898
rect 487328 273454 487648 273486
rect 487328 273218 487370 273454
rect 487606 273218 487648 273454
rect 487328 273134 487648 273218
rect 487328 272898 487370 273134
rect 487606 272898 487648 273134
rect 487328 272866 487648 272898
rect 487328 237454 487648 237486
rect 487328 237218 487370 237454
rect 487606 237218 487648 237454
rect 487328 237134 487648 237218
rect 487328 236898 487370 237134
rect 487606 236898 487648 237134
rect 487328 236866 487648 236898
rect 487328 201454 487648 201486
rect 487328 201218 487370 201454
rect 487606 201218 487648 201454
rect 487328 201134 487648 201218
rect 487328 200898 487370 201134
rect 487606 200898 487648 201134
rect 487328 200866 487648 200898
rect 487328 165454 487648 165486
rect 487328 165218 487370 165454
rect 487606 165218 487648 165454
rect 487328 165134 487648 165218
rect 487328 164898 487370 165134
rect 487606 164898 487648 165134
rect 487328 164866 487648 164898
rect 487794 93454 488414 126400
rect 489686 97885 489746 574910
rect 489867 574908 489868 574910
rect 489932 574908 489933 574972
rect 489867 574907 489933 574908
rect 492811 574972 492877 574973
rect 492811 574908 492812 574972
rect 492876 574908 492877 574972
rect 492811 574907 492877 574908
rect 496859 574972 496925 574973
rect 496859 574908 496860 574972
rect 496924 574908 496925 574972
rect 496859 574907 496925 574908
rect 500907 574972 500973 574973
rect 500907 574908 500908 574972
rect 500972 574908 500973 574972
rect 500907 574907 500973 574908
rect 505139 574972 505205 574973
rect 505139 574908 505140 574972
rect 505204 574908 505205 574972
rect 509187 574972 509253 574973
rect 509187 574970 509188 574972
rect 505139 574907 505205 574908
rect 509006 574910 509188 574970
rect 489683 97884 489749 97885
rect 489683 97820 489684 97884
rect 489748 97820 489749 97884
rect 489683 97819 489749 97820
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 485819 85508 485885 85509
rect 485819 85444 485820 85508
rect 485884 85444 485885 85508
rect 485819 85443 485885 85444
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 97174 492134 126400
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 492814 71773 492874 574907
rect 495234 100894 495854 126400
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 492811 71772 492877 71773
rect 492811 71708 492812 71772
rect 492876 71708 492877 71772
rect 492811 71707 492877 71708
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 496862 45525 496922 574907
rect 498954 104614 499574 126400
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 496859 45524 496925 45525
rect 496859 45460 496860 45524
rect 496924 45460 496925 45524
rect 496859 45459 496925 45460
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 68058
rect 500910 59261 500970 574907
rect 502688 543454 503008 543486
rect 502688 543218 502730 543454
rect 502966 543218 503008 543454
rect 502688 543134 503008 543218
rect 502688 542898 502730 543134
rect 502966 542898 503008 543134
rect 502688 542866 503008 542898
rect 502688 507454 503008 507486
rect 502688 507218 502730 507454
rect 502966 507218 503008 507454
rect 502688 507134 503008 507218
rect 502688 506898 502730 507134
rect 502966 506898 503008 507134
rect 502688 506866 503008 506898
rect 502688 471454 503008 471486
rect 502688 471218 502730 471454
rect 502966 471218 503008 471454
rect 502688 471134 503008 471218
rect 502688 470898 502730 471134
rect 502966 470898 503008 471134
rect 502688 470866 503008 470898
rect 502688 435454 503008 435486
rect 502688 435218 502730 435454
rect 502966 435218 503008 435454
rect 502688 435134 503008 435218
rect 502688 434898 502730 435134
rect 502966 434898 503008 435134
rect 502688 434866 503008 434898
rect 502688 399454 503008 399486
rect 502688 399218 502730 399454
rect 502966 399218 503008 399454
rect 502688 399134 503008 399218
rect 502688 398898 502730 399134
rect 502966 398898 503008 399134
rect 502688 398866 503008 398898
rect 502688 363454 503008 363486
rect 502688 363218 502730 363454
rect 502966 363218 503008 363454
rect 502688 363134 503008 363218
rect 502688 362898 502730 363134
rect 502966 362898 503008 363134
rect 502688 362866 503008 362898
rect 502688 327454 503008 327486
rect 502688 327218 502730 327454
rect 502966 327218 503008 327454
rect 502688 327134 503008 327218
rect 502688 326898 502730 327134
rect 502966 326898 503008 327134
rect 502688 326866 503008 326898
rect 502688 291454 503008 291486
rect 502688 291218 502730 291454
rect 502966 291218 503008 291454
rect 502688 291134 503008 291218
rect 502688 290898 502730 291134
rect 502966 290898 503008 291134
rect 502688 290866 503008 290898
rect 502688 255454 503008 255486
rect 502688 255218 502730 255454
rect 502966 255218 503008 255454
rect 502688 255134 503008 255218
rect 502688 254898 502730 255134
rect 502966 254898 503008 255134
rect 502688 254866 503008 254898
rect 502688 219454 503008 219486
rect 502688 219218 502730 219454
rect 502966 219218 503008 219454
rect 502688 219134 503008 219218
rect 502688 218898 502730 219134
rect 502966 218898 503008 219134
rect 502688 218866 503008 218898
rect 502688 183454 503008 183486
rect 502688 183218 502730 183454
rect 502966 183218 503008 183454
rect 502688 183134 503008 183218
rect 502688 182898 502730 183134
rect 502966 182898 503008 183134
rect 502688 182866 503008 182898
rect 502688 147454 503008 147486
rect 502688 147218 502730 147454
rect 502966 147218 503008 147454
rect 502688 147134 503008 147218
rect 502688 146898 502730 147134
rect 502966 146898 503008 147134
rect 502688 146866 503008 146898
rect 500907 59260 500973 59261
rect 500907 59196 500908 59260
rect 500972 59196 500973 59260
rect 500907 59195 500973 59196
rect 505142 33149 505202 574907
rect 505794 111454 506414 126400
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505139 33148 505205 33149
rect 505139 33084 505140 33148
rect 505204 33084 505205 33148
rect 505139 33083 505205 33084
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 3454 506414 38898
rect 509006 6930 509066 574910
rect 509187 574908 509188 574910
rect 509252 574908 509253 574972
rect 509187 574907 509253 574908
rect 513971 574972 514037 574973
rect 513971 574908 513972 574972
rect 514036 574908 514037 574972
rect 513971 574907 514037 574908
rect 509514 115174 510134 126400
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509006 6901 509250 6930
rect 509006 6900 509253 6901
rect 509006 6870 509188 6900
rect 509187 6836 509188 6870
rect 509252 6836 509253 6900
rect 509187 6835 509253 6836
rect 509514 6854 510134 6938
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 118894 513854 126400
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513974 20637 514034 574907
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 516954 122614 517574 126400
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 513971 20636 514037 20637
rect 513971 20572 513972 20636
rect 514036 20572 514037 20636
rect 513971 20571 514037 20572
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 72650 543218 72886 543454
rect 72650 542898 72886 543134
rect 72650 507218 72886 507454
rect 72650 506898 72886 507134
rect 72650 471218 72886 471454
rect 72650 470898 72886 471134
rect 72650 435218 72886 435454
rect 72650 434898 72886 435134
rect 72650 399218 72886 399454
rect 72650 398898 72886 399134
rect 72650 363218 72886 363454
rect 72650 362898 72886 363134
rect 72650 327218 72886 327454
rect 72650 326898 72886 327134
rect 72650 291218 72886 291454
rect 72650 290898 72886 291134
rect 72650 255218 72886 255454
rect 72650 254898 72886 255134
rect 72650 219218 72886 219454
rect 72650 218898 72886 219134
rect 72650 183218 72886 183454
rect 72650 182898 72886 183134
rect 72650 147218 72886 147454
rect 72650 146898 72886 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 88010 561218 88246 561454
rect 88010 560898 88246 561134
rect 88010 525218 88246 525454
rect 88010 524898 88246 525134
rect 88010 489218 88246 489454
rect 88010 488898 88246 489134
rect 88010 453218 88246 453454
rect 88010 452898 88246 453134
rect 88010 417218 88246 417454
rect 88010 416898 88246 417134
rect 88010 381218 88246 381454
rect 88010 380898 88246 381134
rect 88010 345218 88246 345454
rect 88010 344898 88246 345134
rect 88010 309218 88246 309454
rect 88010 308898 88246 309134
rect 88010 273218 88246 273454
rect 88010 272898 88246 273134
rect 88010 237218 88246 237454
rect 88010 236898 88246 237134
rect 88010 201218 88246 201454
rect 88010 200898 88246 201134
rect 88010 165218 88246 165454
rect 88010 164898 88246 165134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 103370 543218 103606 543454
rect 103370 542898 103606 543134
rect 103370 507218 103606 507454
rect 103370 506898 103606 507134
rect 103370 471218 103606 471454
rect 103370 470898 103606 471134
rect 103370 435218 103606 435454
rect 103370 434898 103606 435134
rect 103370 399218 103606 399454
rect 103370 398898 103606 399134
rect 103370 363218 103606 363454
rect 103370 362898 103606 363134
rect 103370 327218 103606 327454
rect 103370 326898 103606 327134
rect 103370 291218 103606 291454
rect 103370 290898 103606 291134
rect 103370 255218 103606 255454
rect 103370 254898 103606 255134
rect 103370 219218 103606 219454
rect 103370 218898 103606 219134
rect 103370 183218 103606 183454
rect 103370 182898 103606 183134
rect 103370 147218 103606 147454
rect 103370 146898 103606 147134
rect 118730 561218 118966 561454
rect 118730 560898 118966 561134
rect 149450 561218 149686 561454
rect 149450 560898 149686 561134
rect 180170 561218 180406 561454
rect 180170 560898 180406 561134
rect 210890 561218 211126 561454
rect 210890 560898 211126 561134
rect 241610 561218 241846 561454
rect 241610 560898 241846 561134
rect 272330 561218 272566 561454
rect 272330 560898 272566 561134
rect 303050 561218 303286 561454
rect 303050 560898 303286 561134
rect 333770 561218 334006 561454
rect 333770 560898 334006 561134
rect 364490 561218 364726 561454
rect 364490 560898 364726 561134
rect 395210 561218 395446 561454
rect 395210 560898 395446 561134
rect 425930 561218 426166 561454
rect 425930 560898 426166 561134
rect 456650 561218 456886 561454
rect 456650 560898 456886 561134
rect 134090 543218 134326 543454
rect 134090 542898 134326 543134
rect 164810 543218 165046 543454
rect 164810 542898 165046 543134
rect 195530 543218 195766 543454
rect 195530 542898 195766 543134
rect 226250 543218 226486 543454
rect 226250 542898 226486 543134
rect 256970 543218 257206 543454
rect 256970 542898 257206 543134
rect 287690 543218 287926 543454
rect 287690 542898 287926 543134
rect 318410 543218 318646 543454
rect 318410 542898 318646 543134
rect 349130 543218 349366 543454
rect 349130 542898 349366 543134
rect 379850 543218 380086 543454
rect 379850 542898 380086 543134
rect 410570 543218 410806 543454
rect 410570 542898 410806 543134
rect 441290 543218 441526 543454
rect 441290 542898 441526 543134
rect 472010 543218 472246 543454
rect 472010 542898 472246 543134
rect 118730 525218 118966 525454
rect 118730 524898 118966 525134
rect 149450 525218 149686 525454
rect 149450 524898 149686 525134
rect 180170 525218 180406 525454
rect 180170 524898 180406 525134
rect 210890 525218 211126 525454
rect 210890 524898 211126 525134
rect 241610 525218 241846 525454
rect 241610 524898 241846 525134
rect 272330 525218 272566 525454
rect 272330 524898 272566 525134
rect 303050 525218 303286 525454
rect 303050 524898 303286 525134
rect 333770 525218 334006 525454
rect 333770 524898 334006 525134
rect 364490 525218 364726 525454
rect 364490 524898 364726 525134
rect 395210 525218 395446 525454
rect 395210 524898 395446 525134
rect 425930 525218 426166 525454
rect 425930 524898 426166 525134
rect 456650 525218 456886 525454
rect 456650 524898 456886 525134
rect 134090 507218 134326 507454
rect 134090 506898 134326 507134
rect 164810 507218 165046 507454
rect 164810 506898 165046 507134
rect 195530 507218 195766 507454
rect 195530 506898 195766 507134
rect 226250 507218 226486 507454
rect 226250 506898 226486 507134
rect 256970 507218 257206 507454
rect 256970 506898 257206 507134
rect 287690 507218 287926 507454
rect 287690 506898 287926 507134
rect 318410 507218 318646 507454
rect 318410 506898 318646 507134
rect 349130 507218 349366 507454
rect 349130 506898 349366 507134
rect 379850 507218 380086 507454
rect 379850 506898 380086 507134
rect 410570 507218 410806 507454
rect 410570 506898 410806 507134
rect 441290 507218 441526 507454
rect 441290 506898 441526 507134
rect 472010 507218 472246 507454
rect 472010 506898 472246 507134
rect 118730 489218 118966 489454
rect 118730 488898 118966 489134
rect 149450 489218 149686 489454
rect 149450 488898 149686 489134
rect 180170 489218 180406 489454
rect 180170 488898 180406 489134
rect 210890 489218 211126 489454
rect 210890 488898 211126 489134
rect 241610 489218 241846 489454
rect 241610 488898 241846 489134
rect 272330 489218 272566 489454
rect 272330 488898 272566 489134
rect 303050 489218 303286 489454
rect 303050 488898 303286 489134
rect 333770 489218 334006 489454
rect 333770 488898 334006 489134
rect 364490 489218 364726 489454
rect 364490 488898 364726 489134
rect 395210 489218 395446 489454
rect 395210 488898 395446 489134
rect 425930 489218 426166 489454
rect 425930 488898 426166 489134
rect 456650 489218 456886 489454
rect 456650 488898 456886 489134
rect 134090 471218 134326 471454
rect 134090 470898 134326 471134
rect 164810 471218 165046 471454
rect 164810 470898 165046 471134
rect 195530 471218 195766 471454
rect 195530 470898 195766 471134
rect 226250 471218 226486 471454
rect 226250 470898 226486 471134
rect 256970 471218 257206 471454
rect 256970 470898 257206 471134
rect 287690 471218 287926 471454
rect 287690 470898 287926 471134
rect 318410 471218 318646 471454
rect 318410 470898 318646 471134
rect 349130 471218 349366 471454
rect 349130 470898 349366 471134
rect 379850 471218 380086 471454
rect 379850 470898 380086 471134
rect 410570 471218 410806 471454
rect 410570 470898 410806 471134
rect 441290 471218 441526 471454
rect 441290 470898 441526 471134
rect 472010 471218 472246 471454
rect 472010 470898 472246 471134
rect 118730 453218 118966 453454
rect 118730 452898 118966 453134
rect 149450 453218 149686 453454
rect 149450 452898 149686 453134
rect 180170 453218 180406 453454
rect 180170 452898 180406 453134
rect 210890 453218 211126 453454
rect 210890 452898 211126 453134
rect 241610 453218 241846 453454
rect 241610 452898 241846 453134
rect 272330 453218 272566 453454
rect 272330 452898 272566 453134
rect 303050 453218 303286 453454
rect 303050 452898 303286 453134
rect 333770 453218 334006 453454
rect 333770 452898 334006 453134
rect 364490 453218 364726 453454
rect 364490 452898 364726 453134
rect 395210 453218 395446 453454
rect 395210 452898 395446 453134
rect 425930 453218 426166 453454
rect 425930 452898 426166 453134
rect 456650 453218 456886 453454
rect 456650 452898 456886 453134
rect 134090 435218 134326 435454
rect 134090 434898 134326 435134
rect 164810 435218 165046 435454
rect 164810 434898 165046 435134
rect 195530 435218 195766 435454
rect 195530 434898 195766 435134
rect 226250 435218 226486 435454
rect 226250 434898 226486 435134
rect 256970 435218 257206 435454
rect 256970 434898 257206 435134
rect 287690 435218 287926 435454
rect 287690 434898 287926 435134
rect 318410 435218 318646 435454
rect 318410 434898 318646 435134
rect 349130 435218 349366 435454
rect 349130 434898 349366 435134
rect 379850 435218 380086 435454
rect 379850 434898 380086 435134
rect 410570 435218 410806 435454
rect 410570 434898 410806 435134
rect 441290 435218 441526 435454
rect 441290 434898 441526 435134
rect 472010 435218 472246 435454
rect 472010 434898 472246 435134
rect 118730 417218 118966 417454
rect 118730 416898 118966 417134
rect 149450 417218 149686 417454
rect 149450 416898 149686 417134
rect 180170 417218 180406 417454
rect 180170 416898 180406 417134
rect 210890 417218 211126 417454
rect 210890 416898 211126 417134
rect 241610 417218 241846 417454
rect 241610 416898 241846 417134
rect 272330 417218 272566 417454
rect 272330 416898 272566 417134
rect 303050 417218 303286 417454
rect 303050 416898 303286 417134
rect 333770 417218 334006 417454
rect 333770 416898 334006 417134
rect 364490 417218 364726 417454
rect 364490 416898 364726 417134
rect 395210 417218 395446 417454
rect 395210 416898 395446 417134
rect 425930 417218 426166 417454
rect 425930 416898 426166 417134
rect 456650 417218 456886 417454
rect 456650 416898 456886 417134
rect 134090 399218 134326 399454
rect 134090 398898 134326 399134
rect 164810 399218 165046 399454
rect 164810 398898 165046 399134
rect 195530 399218 195766 399454
rect 195530 398898 195766 399134
rect 226250 399218 226486 399454
rect 226250 398898 226486 399134
rect 256970 399218 257206 399454
rect 256970 398898 257206 399134
rect 287690 399218 287926 399454
rect 287690 398898 287926 399134
rect 318410 399218 318646 399454
rect 318410 398898 318646 399134
rect 349130 399218 349366 399454
rect 349130 398898 349366 399134
rect 379850 399218 380086 399454
rect 379850 398898 380086 399134
rect 410570 399218 410806 399454
rect 410570 398898 410806 399134
rect 441290 399218 441526 399454
rect 441290 398898 441526 399134
rect 472010 399218 472246 399454
rect 472010 398898 472246 399134
rect 118730 381218 118966 381454
rect 118730 380898 118966 381134
rect 149450 381218 149686 381454
rect 149450 380898 149686 381134
rect 180170 381218 180406 381454
rect 180170 380898 180406 381134
rect 210890 381218 211126 381454
rect 210890 380898 211126 381134
rect 241610 381218 241846 381454
rect 241610 380898 241846 381134
rect 272330 381218 272566 381454
rect 272330 380898 272566 381134
rect 303050 381218 303286 381454
rect 303050 380898 303286 381134
rect 333770 381218 334006 381454
rect 333770 380898 334006 381134
rect 364490 381218 364726 381454
rect 364490 380898 364726 381134
rect 395210 381218 395446 381454
rect 395210 380898 395446 381134
rect 425930 381218 426166 381454
rect 425930 380898 426166 381134
rect 456650 381218 456886 381454
rect 456650 380898 456886 381134
rect 134090 363218 134326 363454
rect 134090 362898 134326 363134
rect 164810 363218 165046 363454
rect 164810 362898 165046 363134
rect 195530 363218 195766 363454
rect 195530 362898 195766 363134
rect 226250 363218 226486 363454
rect 226250 362898 226486 363134
rect 256970 363218 257206 363454
rect 256970 362898 257206 363134
rect 287690 363218 287926 363454
rect 287690 362898 287926 363134
rect 318410 363218 318646 363454
rect 318410 362898 318646 363134
rect 349130 363218 349366 363454
rect 349130 362898 349366 363134
rect 379850 363218 380086 363454
rect 379850 362898 380086 363134
rect 410570 363218 410806 363454
rect 410570 362898 410806 363134
rect 441290 363218 441526 363454
rect 441290 362898 441526 363134
rect 472010 363218 472246 363454
rect 472010 362898 472246 363134
rect 118730 345218 118966 345454
rect 118730 344898 118966 345134
rect 149450 345218 149686 345454
rect 149450 344898 149686 345134
rect 180170 345218 180406 345454
rect 180170 344898 180406 345134
rect 210890 345218 211126 345454
rect 210890 344898 211126 345134
rect 241610 345218 241846 345454
rect 241610 344898 241846 345134
rect 272330 345218 272566 345454
rect 272330 344898 272566 345134
rect 303050 345218 303286 345454
rect 303050 344898 303286 345134
rect 333770 345218 334006 345454
rect 333770 344898 334006 345134
rect 364490 345218 364726 345454
rect 364490 344898 364726 345134
rect 395210 345218 395446 345454
rect 395210 344898 395446 345134
rect 425930 345218 426166 345454
rect 425930 344898 426166 345134
rect 456650 345218 456886 345454
rect 456650 344898 456886 345134
rect 134090 327218 134326 327454
rect 134090 326898 134326 327134
rect 164810 327218 165046 327454
rect 164810 326898 165046 327134
rect 195530 327218 195766 327454
rect 195530 326898 195766 327134
rect 226250 327218 226486 327454
rect 226250 326898 226486 327134
rect 256970 327218 257206 327454
rect 256970 326898 257206 327134
rect 287690 327218 287926 327454
rect 287690 326898 287926 327134
rect 318410 327218 318646 327454
rect 318410 326898 318646 327134
rect 349130 327218 349366 327454
rect 349130 326898 349366 327134
rect 379850 327218 380086 327454
rect 379850 326898 380086 327134
rect 410570 327218 410806 327454
rect 410570 326898 410806 327134
rect 441290 327218 441526 327454
rect 441290 326898 441526 327134
rect 472010 327218 472246 327454
rect 472010 326898 472246 327134
rect 118730 309218 118966 309454
rect 118730 308898 118966 309134
rect 149450 309218 149686 309454
rect 149450 308898 149686 309134
rect 180170 309218 180406 309454
rect 180170 308898 180406 309134
rect 210890 309218 211126 309454
rect 210890 308898 211126 309134
rect 241610 309218 241846 309454
rect 241610 308898 241846 309134
rect 272330 309218 272566 309454
rect 272330 308898 272566 309134
rect 303050 309218 303286 309454
rect 303050 308898 303286 309134
rect 333770 309218 334006 309454
rect 333770 308898 334006 309134
rect 364490 309218 364726 309454
rect 364490 308898 364726 309134
rect 395210 309218 395446 309454
rect 395210 308898 395446 309134
rect 425930 309218 426166 309454
rect 425930 308898 426166 309134
rect 456650 309218 456886 309454
rect 456650 308898 456886 309134
rect 134090 291218 134326 291454
rect 134090 290898 134326 291134
rect 164810 291218 165046 291454
rect 164810 290898 165046 291134
rect 195530 291218 195766 291454
rect 195530 290898 195766 291134
rect 226250 291218 226486 291454
rect 226250 290898 226486 291134
rect 256970 291218 257206 291454
rect 256970 290898 257206 291134
rect 287690 291218 287926 291454
rect 287690 290898 287926 291134
rect 318410 291218 318646 291454
rect 318410 290898 318646 291134
rect 349130 291218 349366 291454
rect 349130 290898 349366 291134
rect 379850 291218 380086 291454
rect 379850 290898 380086 291134
rect 410570 291218 410806 291454
rect 410570 290898 410806 291134
rect 441290 291218 441526 291454
rect 441290 290898 441526 291134
rect 472010 291218 472246 291454
rect 472010 290898 472246 291134
rect 118730 273218 118966 273454
rect 118730 272898 118966 273134
rect 149450 273218 149686 273454
rect 149450 272898 149686 273134
rect 180170 273218 180406 273454
rect 180170 272898 180406 273134
rect 210890 273218 211126 273454
rect 210890 272898 211126 273134
rect 241610 273218 241846 273454
rect 241610 272898 241846 273134
rect 272330 273218 272566 273454
rect 272330 272898 272566 273134
rect 303050 273218 303286 273454
rect 303050 272898 303286 273134
rect 333770 273218 334006 273454
rect 333770 272898 334006 273134
rect 364490 273218 364726 273454
rect 364490 272898 364726 273134
rect 395210 273218 395446 273454
rect 395210 272898 395446 273134
rect 425930 273218 426166 273454
rect 425930 272898 426166 273134
rect 456650 273218 456886 273454
rect 456650 272898 456886 273134
rect 134090 255218 134326 255454
rect 134090 254898 134326 255134
rect 164810 255218 165046 255454
rect 164810 254898 165046 255134
rect 195530 255218 195766 255454
rect 195530 254898 195766 255134
rect 226250 255218 226486 255454
rect 226250 254898 226486 255134
rect 256970 255218 257206 255454
rect 256970 254898 257206 255134
rect 287690 255218 287926 255454
rect 287690 254898 287926 255134
rect 318410 255218 318646 255454
rect 318410 254898 318646 255134
rect 349130 255218 349366 255454
rect 349130 254898 349366 255134
rect 379850 255218 380086 255454
rect 379850 254898 380086 255134
rect 410570 255218 410806 255454
rect 410570 254898 410806 255134
rect 441290 255218 441526 255454
rect 441290 254898 441526 255134
rect 472010 255218 472246 255454
rect 472010 254898 472246 255134
rect 118730 237218 118966 237454
rect 118730 236898 118966 237134
rect 149450 237218 149686 237454
rect 149450 236898 149686 237134
rect 180170 237218 180406 237454
rect 180170 236898 180406 237134
rect 210890 237218 211126 237454
rect 210890 236898 211126 237134
rect 241610 237218 241846 237454
rect 241610 236898 241846 237134
rect 272330 237218 272566 237454
rect 272330 236898 272566 237134
rect 303050 237218 303286 237454
rect 303050 236898 303286 237134
rect 333770 237218 334006 237454
rect 333770 236898 334006 237134
rect 364490 237218 364726 237454
rect 364490 236898 364726 237134
rect 395210 237218 395446 237454
rect 395210 236898 395446 237134
rect 425930 237218 426166 237454
rect 425930 236898 426166 237134
rect 456650 237218 456886 237454
rect 456650 236898 456886 237134
rect 134090 219218 134326 219454
rect 134090 218898 134326 219134
rect 164810 219218 165046 219454
rect 164810 218898 165046 219134
rect 195530 219218 195766 219454
rect 195530 218898 195766 219134
rect 226250 219218 226486 219454
rect 226250 218898 226486 219134
rect 256970 219218 257206 219454
rect 256970 218898 257206 219134
rect 287690 219218 287926 219454
rect 287690 218898 287926 219134
rect 318410 219218 318646 219454
rect 318410 218898 318646 219134
rect 349130 219218 349366 219454
rect 349130 218898 349366 219134
rect 379850 219218 380086 219454
rect 379850 218898 380086 219134
rect 410570 219218 410806 219454
rect 410570 218898 410806 219134
rect 441290 219218 441526 219454
rect 441290 218898 441526 219134
rect 472010 219218 472246 219454
rect 472010 218898 472246 219134
rect 118730 201218 118966 201454
rect 118730 200898 118966 201134
rect 149450 201218 149686 201454
rect 149450 200898 149686 201134
rect 180170 201218 180406 201454
rect 180170 200898 180406 201134
rect 210890 201218 211126 201454
rect 210890 200898 211126 201134
rect 241610 201218 241846 201454
rect 241610 200898 241846 201134
rect 272330 201218 272566 201454
rect 272330 200898 272566 201134
rect 303050 201218 303286 201454
rect 303050 200898 303286 201134
rect 333770 201218 334006 201454
rect 333770 200898 334006 201134
rect 364490 201218 364726 201454
rect 364490 200898 364726 201134
rect 395210 201218 395446 201454
rect 395210 200898 395446 201134
rect 425930 201218 426166 201454
rect 425930 200898 426166 201134
rect 456650 201218 456886 201454
rect 456650 200898 456886 201134
rect 134090 183218 134326 183454
rect 134090 182898 134326 183134
rect 164810 183218 165046 183454
rect 164810 182898 165046 183134
rect 195530 183218 195766 183454
rect 195530 182898 195766 183134
rect 226250 183218 226486 183454
rect 226250 182898 226486 183134
rect 256970 183218 257206 183454
rect 256970 182898 257206 183134
rect 287690 183218 287926 183454
rect 287690 182898 287926 183134
rect 318410 183218 318646 183454
rect 318410 182898 318646 183134
rect 349130 183218 349366 183454
rect 349130 182898 349366 183134
rect 379850 183218 380086 183454
rect 379850 182898 380086 183134
rect 410570 183218 410806 183454
rect 410570 182898 410806 183134
rect 441290 183218 441526 183454
rect 441290 182898 441526 183134
rect 472010 183218 472246 183454
rect 472010 182898 472246 183134
rect 118730 165218 118966 165454
rect 118730 164898 118966 165134
rect 149450 165218 149686 165454
rect 149450 164898 149686 165134
rect 180170 165218 180406 165454
rect 180170 164898 180406 165134
rect 210890 165218 211126 165454
rect 210890 164898 211126 165134
rect 241610 165218 241846 165454
rect 241610 164898 241846 165134
rect 272330 165218 272566 165454
rect 272330 164898 272566 165134
rect 303050 165218 303286 165454
rect 303050 164898 303286 165134
rect 333770 165218 334006 165454
rect 333770 164898 334006 165134
rect 364490 165218 364726 165454
rect 364490 164898 364726 165134
rect 395210 165218 395446 165454
rect 395210 164898 395446 165134
rect 425930 165218 426166 165454
rect 425930 164898 426166 165134
rect 456650 165218 456886 165454
rect 456650 164898 456886 165134
rect 134090 147218 134326 147454
rect 134090 146898 134326 147134
rect 164810 147218 165046 147454
rect 164810 146898 165046 147134
rect 195530 147218 195766 147454
rect 195530 146898 195766 147134
rect 226250 147218 226486 147454
rect 226250 146898 226486 147134
rect 256970 147218 257206 147454
rect 256970 146898 257206 147134
rect 287690 147218 287926 147454
rect 287690 146898 287926 147134
rect 318410 147218 318646 147454
rect 318410 146898 318646 147134
rect 349130 147218 349366 147454
rect 349130 146898 349366 147134
rect 379850 147218 380086 147454
rect 379850 146898 380086 147134
rect 410570 147218 410806 147454
rect 410570 146898 410806 147134
rect 441290 147218 441526 147454
rect 441290 146898 441526 147134
rect 472010 147218 472246 147454
rect 472010 146898 472246 147134
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 487370 561218 487606 561454
rect 487370 560898 487606 561134
rect 487370 525218 487606 525454
rect 487370 524898 487606 525134
rect 487370 489218 487606 489454
rect 487370 488898 487606 489134
rect 487370 453218 487606 453454
rect 487370 452898 487606 453134
rect 487370 417218 487606 417454
rect 487370 416898 487606 417134
rect 487370 381218 487606 381454
rect 487370 380898 487606 381134
rect 487370 345218 487606 345454
rect 487370 344898 487606 345134
rect 487370 309218 487606 309454
rect 487370 308898 487606 309134
rect 487370 273218 487606 273454
rect 487370 272898 487606 273134
rect 487370 237218 487606 237454
rect 487370 236898 487606 237134
rect 487370 201218 487606 201454
rect 487370 200898 487606 201134
rect 487370 165218 487606 165454
rect 487370 164898 487606 165134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 502730 543218 502966 543454
rect 502730 542898 502966 543134
rect 502730 507218 502966 507454
rect 502730 506898 502966 507134
rect 502730 471218 502966 471454
rect 502730 470898 502966 471134
rect 502730 435218 502966 435454
rect 502730 434898 502966 435134
rect 502730 399218 502966 399454
rect 502730 398898 502966 399134
rect 502730 363218 502966 363454
rect 502730 362898 502966 363134
rect 502730 327218 502966 327454
rect 502730 326898 502966 327134
rect 502730 291218 502966 291454
rect 502730 290898 502966 291134
rect 502730 255218 502966 255454
rect 502730 254898 502966 255134
rect 502730 219218 502966 219454
rect 502730 218898 502966 219134
rect 502730 183218 502966 183454
rect 502730 182898 502966 183134
rect 502730 147218 502966 147454
rect 502730 146898 502966 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 88010 561454
rect 88246 561218 118730 561454
rect 118966 561218 149450 561454
rect 149686 561218 180170 561454
rect 180406 561218 210890 561454
rect 211126 561218 241610 561454
rect 241846 561218 272330 561454
rect 272566 561218 303050 561454
rect 303286 561218 333770 561454
rect 334006 561218 364490 561454
rect 364726 561218 395210 561454
rect 395446 561218 425930 561454
rect 426166 561218 456650 561454
rect 456886 561218 487370 561454
rect 487606 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 88010 561134
rect 88246 560898 118730 561134
rect 118966 560898 149450 561134
rect 149686 560898 180170 561134
rect 180406 560898 210890 561134
rect 211126 560898 241610 561134
rect 241846 560898 272330 561134
rect 272566 560898 303050 561134
rect 303286 560898 333770 561134
rect 334006 560898 364490 561134
rect 364726 560898 395210 561134
rect 395446 560898 425930 561134
rect 426166 560898 456650 561134
rect 456886 560898 487370 561134
rect 487606 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 72650 543454
rect 72886 543218 103370 543454
rect 103606 543218 134090 543454
rect 134326 543218 164810 543454
rect 165046 543218 195530 543454
rect 195766 543218 226250 543454
rect 226486 543218 256970 543454
rect 257206 543218 287690 543454
rect 287926 543218 318410 543454
rect 318646 543218 349130 543454
rect 349366 543218 379850 543454
rect 380086 543218 410570 543454
rect 410806 543218 441290 543454
rect 441526 543218 472010 543454
rect 472246 543218 502730 543454
rect 502966 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 72650 543134
rect 72886 542898 103370 543134
rect 103606 542898 134090 543134
rect 134326 542898 164810 543134
rect 165046 542898 195530 543134
rect 195766 542898 226250 543134
rect 226486 542898 256970 543134
rect 257206 542898 287690 543134
rect 287926 542898 318410 543134
rect 318646 542898 349130 543134
rect 349366 542898 379850 543134
rect 380086 542898 410570 543134
rect 410806 542898 441290 543134
rect 441526 542898 472010 543134
rect 472246 542898 502730 543134
rect 502966 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 88010 525454
rect 88246 525218 118730 525454
rect 118966 525218 149450 525454
rect 149686 525218 180170 525454
rect 180406 525218 210890 525454
rect 211126 525218 241610 525454
rect 241846 525218 272330 525454
rect 272566 525218 303050 525454
rect 303286 525218 333770 525454
rect 334006 525218 364490 525454
rect 364726 525218 395210 525454
rect 395446 525218 425930 525454
rect 426166 525218 456650 525454
rect 456886 525218 487370 525454
rect 487606 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 88010 525134
rect 88246 524898 118730 525134
rect 118966 524898 149450 525134
rect 149686 524898 180170 525134
rect 180406 524898 210890 525134
rect 211126 524898 241610 525134
rect 241846 524898 272330 525134
rect 272566 524898 303050 525134
rect 303286 524898 333770 525134
rect 334006 524898 364490 525134
rect 364726 524898 395210 525134
rect 395446 524898 425930 525134
rect 426166 524898 456650 525134
rect 456886 524898 487370 525134
rect 487606 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 72650 507454
rect 72886 507218 103370 507454
rect 103606 507218 134090 507454
rect 134326 507218 164810 507454
rect 165046 507218 195530 507454
rect 195766 507218 226250 507454
rect 226486 507218 256970 507454
rect 257206 507218 287690 507454
rect 287926 507218 318410 507454
rect 318646 507218 349130 507454
rect 349366 507218 379850 507454
rect 380086 507218 410570 507454
rect 410806 507218 441290 507454
rect 441526 507218 472010 507454
rect 472246 507218 502730 507454
rect 502966 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 72650 507134
rect 72886 506898 103370 507134
rect 103606 506898 134090 507134
rect 134326 506898 164810 507134
rect 165046 506898 195530 507134
rect 195766 506898 226250 507134
rect 226486 506898 256970 507134
rect 257206 506898 287690 507134
rect 287926 506898 318410 507134
rect 318646 506898 349130 507134
rect 349366 506898 379850 507134
rect 380086 506898 410570 507134
rect 410806 506898 441290 507134
rect 441526 506898 472010 507134
rect 472246 506898 502730 507134
rect 502966 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 88010 489454
rect 88246 489218 118730 489454
rect 118966 489218 149450 489454
rect 149686 489218 180170 489454
rect 180406 489218 210890 489454
rect 211126 489218 241610 489454
rect 241846 489218 272330 489454
rect 272566 489218 303050 489454
rect 303286 489218 333770 489454
rect 334006 489218 364490 489454
rect 364726 489218 395210 489454
rect 395446 489218 425930 489454
rect 426166 489218 456650 489454
rect 456886 489218 487370 489454
rect 487606 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 88010 489134
rect 88246 488898 118730 489134
rect 118966 488898 149450 489134
rect 149686 488898 180170 489134
rect 180406 488898 210890 489134
rect 211126 488898 241610 489134
rect 241846 488898 272330 489134
rect 272566 488898 303050 489134
rect 303286 488898 333770 489134
rect 334006 488898 364490 489134
rect 364726 488898 395210 489134
rect 395446 488898 425930 489134
rect 426166 488898 456650 489134
rect 456886 488898 487370 489134
rect 487606 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 72650 471454
rect 72886 471218 103370 471454
rect 103606 471218 134090 471454
rect 134326 471218 164810 471454
rect 165046 471218 195530 471454
rect 195766 471218 226250 471454
rect 226486 471218 256970 471454
rect 257206 471218 287690 471454
rect 287926 471218 318410 471454
rect 318646 471218 349130 471454
rect 349366 471218 379850 471454
rect 380086 471218 410570 471454
rect 410806 471218 441290 471454
rect 441526 471218 472010 471454
rect 472246 471218 502730 471454
rect 502966 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 72650 471134
rect 72886 470898 103370 471134
rect 103606 470898 134090 471134
rect 134326 470898 164810 471134
rect 165046 470898 195530 471134
rect 195766 470898 226250 471134
rect 226486 470898 256970 471134
rect 257206 470898 287690 471134
rect 287926 470898 318410 471134
rect 318646 470898 349130 471134
rect 349366 470898 379850 471134
rect 380086 470898 410570 471134
rect 410806 470898 441290 471134
rect 441526 470898 472010 471134
rect 472246 470898 502730 471134
rect 502966 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 88010 453454
rect 88246 453218 118730 453454
rect 118966 453218 149450 453454
rect 149686 453218 180170 453454
rect 180406 453218 210890 453454
rect 211126 453218 241610 453454
rect 241846 453218 272330 453454
rect 272566 453218 303050 453454
rect 303286 453218 333770 453454
rect 334006 453218 364490 453454
rect 364726 453218 395210 453454
rect 395446 453218 425930 453454
rect 426166 453218 456650 453454
rect 456886 453218 487370 453454
rect 487606 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 88010 453134
rect 88246 452898 118730 453134
rect 118966 452898 149450 453134
rect 149686 452898 180170 453134
rect 180406 452898 210890 453134
rect 211126 452898 241610 453134
rect 241846 452898 272330 453134
rect 272566 452898 303050 453134
rect 303286 452898 333770 453134
rect 334006 452898 364490 453134
rect 364726 452898 395210 453134
rect 395446 452898 425930 453134
rect 426166 452898 456650 453134
rect 456886 452898 487370 453134
rect 487606 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 72650 435454
rect 72886 435218 103370 435454
rect 103606 435218 134090 435454
rect 134326 435218 164810 435454
rect 165046 435218 195530 435454
rect 195766 435218 226250 435454
rect 226486 435218 256970 435454
rect 257206 435218 287690 435454
rect 287926 435218 318410 435454
rect 318646 435218 349130 435454
rect 349366 435218 379850 435454
rect 380086 435218 410570 435454
rect 410806 435218 441290 435454
rect 441526 435218 472010 435454
rect 472246 435218 502730 435454
rect 502966 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 72650 435134
rect 72886 434898 103370 435134
rect 103606 434898 134090 435134
rect 134326 434898 164810 435134
rect 165046 434898 195530 435134
rect 195766 434898 226250 435134
rect 226486 434898 256970 435134
rect 257206 434898 287690 435134
rect 287926 434898 318410 435134
rect 318646 434898 349130 435134
rect 349366 434898 379850 435134
rect 380086 434898 410570 435134
rect 410806 434898 441290 435134
rect 441526 434898 472010 435134
rect 472246 434898 502730 435134
rect 502966 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88010 417454
rect 88246 417218 118730 417454
rect 118966 417218 149450 417454
rect 149686 417218 180170 417454
rect 180406 417218 210890 417454
rect 211126 417218 241610 417454
rect 241846 417218 272330 417454
rect 272566 417218 303050 417454
rect 303286 417218 333770 417454
rect 334006 417218 364490 417454
rect 364726 417218 395210 417454
rect 395446 417218 425930 417454
rect 426166 417218 456650 417454
rect 456886 417218 487370 417454
rect 487606 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88010 417134
rect 88246 416898 118730 417134
rect 118966 416898 149450 417134
rect 149686 416898 180170 417134
rect 180406 416898 210890 417134
rect 211126 416898 241610 417134
rect 241846 416898 272330 417134
rect 272566 416898 303050 417134
rect 303286 416898 333770 417134
rect 334006 416898 364490 417134
rect 364726 416898 395210 417134
rect 395446 416898 425930 417134
rect 426166 416898 456650 417134
rect 456886 416898 487370 417134
rect 487606 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 72650 399454
rect 72886 399218 103370 399454
rect 103606 399218 134090 399454
rect 134326 399218 164810 399454
rect 165046 399218 195530 399454
rect 195766 399218 226250 399454
rect 226486 399218 256970 399454
rect 257206 399218 287690 399454
rect 287926 399218 318410 399454
rect 318646 399218 349130 399454
rect 349366 399218 379850 399454
rect 380086 399218 410570 399454
rect 410806 399218 441290 399454
rect 441526 399218 472010 399454
rect 472246 399218 502730 399454
rect 502966 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 72650 399134
rect 72886 398898 103370 399134
rect 103606 398898 134090 399134
rect 134326 398898 164810 399134
rect 165046 398898 195530 399134
rect 195766 398898 226250 399134
rect 226486 398898 256970 399134
rect 257206 398898 287690 399134
rect 287926 398898 318410 399134
rect 318646 398898 349130 399134
rect 349366 398898 379850 399134
rect 380086 398898 410570 399134
rect 410806 398898 441290 399134
rect 441526 398898 472010 399134
rect 472246 398898 502730 399134
rect 502966 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 88010 381454
rect 88246 381218 118730 381454
rect 118966 381218 149450 381454
rect 149686 381218 180170 381454
rect 180406 381218 210890 381454
rect 211126 381218 241610 381454
rect 241846 381218 272330 381454
rect 272566 381218 303050 381454
rect 303286 381218 333770 381454
rect 334006 381218 364490 381454
rect 364726 381218 395210 381454
rect 395446 381218 425930 381454
rect 426166 381218 456650 381454
rect 456886 381218 487370 381454
rect 487606 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 88010 381134
rect 88246 380898 118730 381134
rect 118966 380898 149450 381134
rect 149686 380898 180170 381134
rect 180406 380898 210890 381134
rect 211126 380898 241610 381134
rect 241846 380898 272330 381134
rect 272566 380898 303050 381134
rect 303286 380898 333770 381134
rect 334006 380898 364490 381134
rect 364726 380898 395210 381134
rect 395446 380898 425930 381134
rect 426166 380898 456650 381134
rect 456886 380898 487370 381134
rect 487606 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 72650 363454
rect 72886 363218 103370 363454
rect 103606 363218 134090 363454
rect 134326 363218 164810 363454
rect 165046 363218 195530 363454
rect 195766 363218 226250 363454
rect 226486 363218 256970 363454
rect 257206 363218 287690 363454
rect 287926 363218 318410 363454
rect 318646 363218 349130 363454
rect 349366 363218 379850 363454
rect 380086 363218 410570 363454
rect 410806 363218 441290 363454
rect 441526 363218 472010 363454
rect 472246 363218 502730 363454
rect 502966 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 72650 363134
rect 72886 362898 103370 363134
rect 103606 362898 134090 363134
rect 134326 362898 164810 363134
rect 165046 362898 195530 363134
rect 195766 362898 226250 363134
rect 226486 362898 256970 363134
rect 257206 362898 287690 363134
rect 287926 362898 318410 363134
rect 318646 362898 349130 363134
rect 349366 362898 379850 363134
rect 380086 362898 410570 363134
rect 410806 362898 441290 363134
rect 441526 362898 472010 363134
rect 472246 362898 502730 363134
rect 502966 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 88010 345454
rect 88246 345218 118730 345454
rect 118966 345218 149450 345454
rect 149686 345218 180170 345454
rect 180406 345218 210890 345454
rect 211126 345218 241610 345454
rect 241846 345218 272330 345454
rect 272566 345218 303050 345454
rect 303286 345218 333770 345454
rect 334006 345218 364490 345454
rect 364726 345218 395210 345454
rect 395446 345218 425930 345454
rect 426166 345218 456650 345454
rect 456886 345218 487370 345454
rect 487606 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 88010 345134
rect 88246 344898 118730 345134
rect 118966 344898 149450 345134
rect 149686 344898 180170 345134
rect 180406 344898 210890 345134
rect 211126 344898 241610 345134
rect 241846 344898 272330 345134
rect 272566 344898 303050 345134
rect 303286 344898 333770 345134
rect 334006 344898 364490 345134
rect 364726 344898 395210 345134
rect 395446 344898 425930 345134
rect 426166 344898 456650 345134
rect 456886 344898 487370 345134
rect 487606 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 72650 327454
rect 72886 327218 103370 327454
rect 103606 327218 134090 327454
rect 134326 327218 164810 327454
rect 165046 327218 195530 327454
rect 195766 327218 226250 327454
rect 226486 327218 256970 327454
rect 257206 327218 287690 327454
rect 287926 327218 318410 327454
rect 318646 327218 349130 327454
rect 349366 327218 379850 327454
rect 380086 327218 410570 327454
rect 410806 327218 441290 327454
rect 441526 327218 472010 327454
rect 472246 327218 502730 327454
rect 502966 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 72650 327134
rect 72886 326898 103370 327134
rect 103606 326898 134090 327134
rect 134326 326898 164810 327134
rect 165046 326898 195530 327134
rect 195766 326898 226250 327134
rect 226486 326898 256970 327134
rect 257206 326898 287690 327134
rect 287926 326898 318410 327134
rect 318646 326898 349130 327134
rect 349366 326898 379850 327134
rect 380086 326898 410570 327134
rect 410806 326898 441290 327134
rect 441526 326898 472010 327134
rect 472246 326898 502730 327134
rect 502966 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 88010 309454
rect 88246 309218 118730 309454
rect 118966 309218 149450 309454
rect 149686 309218 180170 309454
rect 180406 309218 210890 309454
rect 211126 309218 241610 309454
rect 241846 309218 272330 309454
rect 272566 309218 303050 309454
rect 303286 309218 333770 309454
rect 334006 309218 364490 309454
rect 364726 309218 395210 309454
rect 395446 309218 425930 309454
rect 426166 309218 456650 309454
rect 456886 309218 487370 309454
rect 487606 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 88010 309134
rect 88246 308898 118730 309134
rect 118966 308898 149450 309134
rect 149686 308898 180170 309134
rect 180406 308898 210890 309134
rect 211126 308898 241610 309134
rect 241846 308898 272330 309134
rect 272566 308898 303050 309134
rect 303286 308898 333770 309134
rect 334006 308898 364490 309134
rect 364726 308898 395210 309134
rect 395446 308898 425930 309134
rect 426166 308898 456650 309134
rect 456886 308898 487370 309134
rect 487606 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 72650 291454
rect 72886 291218 103370 291454
rect 103606 291218 134090 291454
rect 134326 291218 164810 291454
rect 165046 291218 195530 291454
rect 195766 291218 226250 291454
rect 226486 291218 256970 291454
rect 257206 291218 287690 291454
rect 287926 291218 318410 291454
rect 318646 291218 349130 291454
rect 349366 291218 379850 291454
rect 380086 291218 410570 291454
rect 410806 291218 441290 291454
rect 441526 291218 472010 291454
rect 472246 291218 502730 291454
rect 502966 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 72650 291134
rect 72886 290898 103370 291134
rect 103606 290898 134090 291134
rect 134326 290898 164810 291134
rect 165046 290898 195530 291134
rect 195766 290898 226250 291134
rect 226486 290898 256970 291134
rect 257206 290898 287690 291134
rect 287926 290898 318410 291134
rect 318646 290898 349130 291134
rect 349366 290898 379850 291134
rect 380086 290898 410570 291134
rect 410806 290898 441290 291134
rect 441526 290898 472010 291134
rect 472246 290898 502730 291134
rect 502966 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 88010 273454
rect 88246 273218 118730 273454
rect 118966 273218 149450 273454
rect 149686 273218 180170 273454
rect 180406 273218 210890 273454
rect 211126 273218 241610 273454
rect 241846 273218 272330 273454
rect 272566 273218 303050 273454
rect 303286 273218 333770 273454
rect 334006 273218 364490 273454
rect 364726 273218 395210 273454
rect 395446 273218 425930 273454
rect 426166 273218 456650 273454
rect 456886 273218 487370 273454
rect 487606 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 88010 273134
rect 88246 272898 118730 273134
rect 118966 272898 149450 273134
rect 149686 272898 180170 273134
rect 180406 272898 210890 273134
rect 211126 272898 241610 273134
rect 241846 272898 272330 273134
rect 272566 272898 303050 273134
rect 303286 272898 333770 273134
rect 334006 272898 364490 273134
rect 364726 272898 395210 273134
rect 395446 272898 425930 273134
rect 426166 272898 456650 273134
rect 456886 272898 487370 273134
rect 487606 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 72650 255454
rect 72886 255218 103370 255454
rect 103606 255218 134090 255454
rect 134326 255218 164810 255454
rect 165046 255218 195530 255454
rect 195766 255218 226250 255454
rect 226486 255218 256970 255454
rect 257206 255218 287690 255454
rect 287926 255218 318410 255454
rect 318646 255218 349130 255454
rect 349366 255218 379850 255454
rect 380086 255218 410570 255454
rect 410806 255218 441290 255454
rect 441526 255218 472010 255454
rect 472246 255218 502730 255454
rect 502966 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 72650 255134
rect 72886 254898 103370 255134
rect 103606 254898 134090 255134
rect 134326 254898 164810 255134
rect 165046 254898 195530 255134
rect 195766 254898 226250 255134
rect 226486 254898 256970 255134
rect 257206 254898 287690 255134
rect 287926 254898 318410 255134
rect 318646 254898 349130 255134
rect 349366 254898 379850 255134
rect 380086 254898 410570 255134
rect 410806 254898 441290 255134
rect 441526 254898 472010 255134
rect 472246 254898 502730 255134
rect 502966 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 88010 237454
rect 88246 237218 118730 237454
rect 118966 237218 149450 237454
rect 149686 237218 180170 237454
rect 180406 237218 210890 237454
rect 211126 237218 241610 237454
rect 241846 237218 272330 237454
rect 272566 237218 303050 237454
rect 303286 237218 333770 237454
rect 334006 237218 364490 237454
rect 364726 237218 395210 237454
rect 395446 237218 425930 237454
rect 426166 237218 456650 237454
rect 456886 237218 487370 237454
rect 487606 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 88010 237134
rect 88246 236898 118730 237134
rect 118966 236898 149450 237134
rect 149686 236898 180170 237134
rect 180406 236898 210890 237134
rect 211126 236898 241610 237134
rect 241846 236898 272330 237134
rect 272566 236898 303050 237134
rect 303286 236898 333770 237134
rect 334006 236898 364490 237134
rect 364726 236898 395210 237134
rect 395446 236898 425930 237134
rect 426166 236898 456650 237134
rect 456886 236898 487370 237134
rect 487606 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 72650 219454
rect 72886 219218 103370 219454
rect 103606 219218 134090 219454
rect 134326 219218 164810 219454
rect 165046 219218 195530 219454
rect 195766 219218 226250 219454
rect 226486 219218 256970 219454
rect 257206 219218 287690 219454
rect 287926 219218 318410 219454
rect 318646 219218 349130 219454
rect 349366 219218 379850 219454
rect 380086 219218 410570 219454
rect 410806 219218 441290 219454
rect 441526 219218 472010 219454
rect 472246 219218 502730 219454
rect 502966 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 72650 219134
rect 72886 218898 103370 219134
rect 103606 218898 134090 219134
rect 134326 218898 164810 219134
rect 165046 218898 195530 219134
rect 195766 218898 226250 219134
rect 226486 218898 256970 219134
rect 257206 218898 287690 219134
rect 287926 218898 318410 219134
rect 318646 218898 349130 219134
rect 349366 218898 379850 219134
rect 380086 218898 410570 219134
rect 410806 218898 441290 219134
rect 441526 218898 472010 219134
rect 472246 218898 502730 219134
rect 502966 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 88010 201454
rect 88246 201218 118730 201454
rect 118966 201218 149450 201454
rect 149686 201218 180170 201454
rect 180406 201218 210890 201454
rect 211126 201218 241610 201454
rect 241846 201218 272330 201454
rect 272566 201218 303050 201454
rect 303286 201218 333770 201454
rect 334006 201218 364490 201454
rect 364726 201218 395210 201454
rect 395446 201218 425930 201454
rect 426166 201218 456650 201454
rect 456886 201218 487370 201454
rect 487606 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 88010 201134
rect 88246 200898 118730 201134
rect 118966 200898 149450 201134
rect 149686 200898 180170 201134
rect 180406 200898 210890 201134
rect 211126 200898 241610 201134
rect 241846 200898 272330 201134
rect 272566 200898 303050 201134
rect 303286 200898 333770 201134
rect 334006 200898 364490 201134
rect 364726 200898 395210 201134
rect 395446 200898 425930 201134
rect 426166 200898 456650 201134
rect 456886 200898 487370 201134
rect 487606 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 72650 183454
rect 72886 183218 103370 183454
rect 103606 183218 134090 183454
rect 134326 183218 164810 183454
rect 165046 183218 195530 183454
rect 195766 183218 226250 183454
rect 226486 183218 256970 183454
rect 257206 183218 287690 183454
rect 287926 183218 318410 183454
rect 318646 183218 349130 183454
rect 349366 183218 379850 183454
rect 380086 183218 410570 183454
rect 410806 183218 441290 183454
rect 441526 183218 472010 183454
rect 472246 183218 502730 183454
rect 502966 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 72650 183134
rect 72886 182898 103370 183134
rect 103606 182898 134090 183134
rect 134326 182898 164810 183134
rect 165046 182898 195530 183134
rect 195766 182898 226250 183134
rect 226486 182898 256970 183134
rect 257206 182898 287690 183134
rect 287926 182898 318410 183134
rect 318646 182898 349130 183134
rect 349366 182898 379850 183134
rect 380086 182898 410570 183134
rect 410806 182898 441290 183134
rect 441526 182898 472010 183134
rect 472246 182898 502730 183134
rect 502966 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 88010 165454
rect 88246 165218 118730 165454
rect 118966 165218 149450 165454
rect 149686 165218 180170 165454
rect 180406 165218 210890 165454
rect 211126 165218 241610 165454
rect 241846 165218 272330 165454
rect 272566 165218 303050 165454
rect 303286 165218 333770 165454
rect 334006 165218 364490 165454
rect 364726 165218 395210 165454
rect 395446 165218 425930 165454
rect 426166 165218 456650 165454
rect 456886 165218 487370 165454
rect 487606 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 88010 165134
rect 88246 164898 118730 165134
rect 118966 164898 149450 165134
rect 149686 164898 180170 165134
rect 180406 164898 210890 165134
rect 211126 164898 241610 165134
rect 241846 164898 272330 165134
rect 272566 164898 303050 165134
rect 303286 164898 333770 165134
rect 334006 164898 364490 165134
rect 364726 164898 395210 165134
rect 395446 164898 425930 165134
rect 426166 164898 456650 165134
rect 456886 164898 487370 165134
rect 487606 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 72650 147454
rect 72886 147218 103370 147454
rect 103606 147218 134090 147454
rect 134326 147218 164810 147454
rect 165046 147218 195530 147454
rect 195766 147218 226250 147454
rect 226486 147218 256970 147454
rect 257206 147218 287690 147454
rect 287926 147218 318410 147454
rect 318646 147218 349130 147454
rect 349366 147218 379850 147454
rect 380086 147218 410570 147454
rect 410806 147218 441290 147454
rect 441526 147218 472010 147454
rect 472246 147218 502730 147454
rect 502966 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 72650 147134
rect 72886 146898 103370 147134
rect 103606 146898 134090 147134
rect 134326 146898 164810 147134
rect 165046 146898 195530 147134
rect 195766 146898 226250 147134
rect 226486 146898 256970 147134
rect 257206 146898 287690 147134
rect 287926 146898 318410 147134
rect 318646 146898 349130 147134
rect 349366 146898 379850 147134
rect 380086 146898 410570 147134
rect 410806 146898 441290 147134
rect 441526 146898 472010 147134
rect 472246 146898 502730 147134
rect 502966 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1635447575
transform 1 0 68400 0 1 128400
box 382 0 446738 447200
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 126400 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 577600 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 577600 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 577600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 577600 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 577600 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 577600 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 577600 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 577600 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 577600 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 577600 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 577600 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 577600 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 577600 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 126400 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 577600 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 577600 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 577600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 577600 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 577600 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 577600 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 577600 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 577600 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 577600 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 577600 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 577600 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 577600 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 577600 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 126400 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 577600 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 577600 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 577600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 577600 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 577600 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 577600 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 577600 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 577600 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 577600 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 577600 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 577600 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 577600 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 577600 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 126400 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 577600 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 577600 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 577600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 577600 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 577600 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 577600 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 577600 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 577600 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 577600 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 577600 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 577600 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 577600 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 577600 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 126400 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 577600 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 577600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 577600 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 577600 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 577600 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 577600 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 577600 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 577600 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 577600 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 577600 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 577600 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 577600 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 126400 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 577600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 577600 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 577600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 577600 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 577600 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 577600 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 577600 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 577600 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 577600 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 577600 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 577600 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 577600 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 577600 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 126400 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 577600 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 577600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 577600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 577600 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 577600 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 577600 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 577600 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 577600 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 577600 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 577600 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 577600 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 577600 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 126400 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 577600 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 577600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 577600 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 577600 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 577600 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 577600 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 577600 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 577600 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 577600 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 577600 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 577600 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 577600 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
