magic
tech sky130A
magscale 1 2
timestamp 1636060364
<< locali >>
rect 84301 545207 84335 545377
rect 515505 39899 515539 40001
rect 155141 38743 155175 39525
rect 541173 39287 541207 39593
rect 53849 3383 53883 3893
rect 546785 3043 546819 3417
rect 552673 2975 552707 3349
rect 582389 3043 582423 39321
rect 552765 2839 552799 2941
rect 552615 2805 552799 2839
<< viali >>
rect 84301 545377 84335 545411
rect 84301 545173 84335 545207
rect 515505 40001 515539 40035
rect 515505 39865 515539 39899
rect 541173 39593 541207 39627
rect 155141 39525 155175 39559
rect 541173 39253 541207 39287
rect 582389 39321 582423 39355
rect 155141 38709 155175 38743
rect 53849 3893 53883 3927
rect 53849 3349 53883 3383
rect 546785 3417 546819 3451
rect 546785 3009 546819 3043
rect 552673 3349 552707 3383
rect 582389 3009 582423 3043
rect 552673 2941 552707 2975
rect 552765 2941 552799 2975
rect 552581 2805 552615 2839
<< metal1 >>
rect 273162 700952 273168 701004
rect 273220 700992 273226 701004
rect 397454 700992 397460 701004
rect 273220 700964 397460 700992
rect 273220 700952 273226 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 154114 700884 154120 700936
rect 154172 700924 154178 700936
rect 268378 700924 268384 700936
rect 154172 700896 268384 700924
rect 154172 700884 154178 700896
rect 268378 700884 268384 700896
rect 268436 700884 268442 700936
rect 278682 700884 278688 700936
rect 278740 700924 278746 700936
rect 413646 700924 413652 700936
rect 278740 700896 413652 700924
rect 278740 700884 278746 700896
rect 413646 700884 413652 700896
rect 413704 700884 413710 700936
rect 137830 700816 137836 700868
rect 137888 700856 137894 700868
rect 325694 700856 325700 700868
rect 137888 700828 325700 700856
rect 137888 700816 137894 700828
rect 325694 700816 325700 700828
rect 325752 700816 325758 700868
rect 331858 700816 331864 700868
rect 331916 700856 331922 700868
rect 494790 700856 494796 700868
rect 331916 700828 494796 700856
rect 331916 700816 331922 700828
rect 494790 700816 494796 700828
rect 494848 700816 494854 700868
rect 89162 700748 89168 700800
rect 89220 700788 89226 700800
rect 93118 700788 93124 700800
rect 89220 700760 93124 700788
rect 89220 700748 89226 700760
rect 93118 700748 93124 700760
rect 93176 700748 93182 700800
rect 260742 700748 260748 700800
rect 260800 700788 260806 700800
rect 462314 700788 462320 700800
rect 260800 700760 462320 700788
rect 260800 700748 260806 700760
rect 462314 700748 462320 700760
rect 462372 700748 462378 700800
rect 218974 700680 218980 700732
rect 219032 700720 219038 700732
rect 255958 700720 255964 700732
rect 219032 700692 255964 700720
rect 219032 700680 219038 700692
rect 255958 700680 255964 700692
rect 256016 700680 256022 700732
rect 264882 700680 264888 700732
rect 264940 700720 264946 700732
rect 478506 700720 478512 700732
rect 264940 700692 478512 700720
rect 264940 700680 264946 700692
rect 478506 700680 478512 700692
rect 478564 700680 478570 700732
rect 105446 700612 105452 700664
rect 105504 700652 105510 700664
rect 333974 700652 333980 700664
rect 105504 700624 333980 700652
rect 105504 700612 105510 700624
rect 333974 700612 333980 700624
rect 334032 700612 334038 700664
rect 72970 700544 72976 700596
rect 73028 700584 73034 700596
rect 338114 700584 338120 700596
rect 73028 700556 338120 700584
rect 73028 700544 73034 700556
rect 338114 700544 338120 700556
rect 338172 700544 338178 700596
rect 246942 700476 246948 700528
rect 247000 700516 247006 700528
rect 527174 700516 527180 700528
rect 247000 700488 527180 700516
rect 247000 700476 247006 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 24302 700408 24308 700460
rect 24360 700448 24366 700460
rect 65518 700448 65524 700460
rect 24360 700420 65524 700448
rect 24360 700408 24366 700420
rect 65518 700408 65524 700420
rect 65576 700408 65582 700460
rect 170306 700408 170312 700460
rect 170364 700448 170370 700460
rect 180058 700448 180064 700460
rect 170364 700420 180064 700448
rect 170364 700408 170370 700420
rect 180058 700408 180064 700420
rect 180116 700408 180122 700460
rect 235166 700408 235172 700460
rect 235224 700448 235230 700460
rect 242158 700448 242164 700460
rect 235224 700420 242164 700448
rect 235224 700408 235230 700420
rect 242158 700408 242164 700420
rect 242216 700408 242222 700460
rect 251082 700408 251088 700460
rect 251140 700448 251146 700460
rect 543458 700448 543464 700460
rect 251140 700420 543464 700448
rect 251140 700408 251146 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 347774 700380 347780 700392
rect 40552 700352 347780 700380
rect 40552 700340 40558 700352
rect 347774 700340 347780 700352
rect 347832 700340 347838 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 351914 700312 351920 700324
rect 8168 700284 351920 700312
rect 8168 700272 8174 700284
rect 351914 700272 351920 700284
rect 351972 700272 351978 700324
rect 400858 700272 400864 700324
rect 400916 700312 400922 700324
rect 429838 700312 429844 700324
rect 400916 700284 429844 700312
rect 400916 700272 400922 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 538858 700272 538864 700324
rect 538916 700312 538922 700324
rect 559650 700312 559656 700324
rect 538916 700284 559656 700312
rect 538916 700272 538922 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 202782 700204 202788 700256
rect 202840 700244 202846 700256
rect 311894 700244 311900 700256
rect 202840 700216 311900 700244
rect 202840 700204 202846 700216
rect 311894 700204 311900 700216
rect 311952 700204 311958 700256
rect 324958 700204 324964 700256
rect 325016 700244 325022 700256
rect 364978 700244 364984 700256
rect 325016 700216 364984 700244
rect 325016 700204 325022 700216
rect 364978 700204 364984 700216
rect 365036 700204 365042 700256
rect 291102 700136 291108 700188
rect 291160 700176 291166 700188
rect 348786 700176 348792 700188
rect 291160 700148 348792 700176
rect 291160 700136 291166 700148
rect 348786 700136 348792 700148
rect 348844 700136 348850 700188
rect 286962 700068 286968 700120
rect 287020 700108 287026 700120
rect 332502 700108 332508 700120
rect 287020 700080 332508 700108
rect 287020 700068 287026 700080
rect 332502 700068 332508 700080
rect 332560 700068 332566 700120
rect 267642 700000 267648 700052
rect 267700 700040 267706 700052
rect 299474 700040 299480 700052
rect 267700 700012 299480 700040
rect 267700 700000 267706 700012
rect 299474 700000 299480 700012
rect 299532 700000 299538 700052
rect 283834 699932 283840 699984
rect 283892 699972 283898 699984
rect 303614 699972 303620 699984
rect 283892 699944 303620 699972
rect 283892 699932 283898 699944
rect 303614 699932 303620 699944
rect 303672 699932 303678 699984
rect 234522 696940 234528 696992
rect 234580 696980 234586 696992
rect 580166 696980 580172 696992
rect 234580 696952 580172 696980
rect 234580 696940 234586 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 238662 683204 238668 683256
rect 238720 683244 238726 683256
rect 580166 683244 580172 683256
rect 238720 683216 580172 683244
rect 238720 683204 238726 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 360194 683176 360200 683188
rect 3476 683148 360200 683176
rect 3476 683136 3482 683148
rect 360194 683136 360200 683148
rect 360252 683136 360258 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 61378 670732 61384 670744
rect 3568 670704 61384 670732
rect 3568 670692 3574 670704
rect 61378 670692 61384 670704
rect 61436 670692 61442 670744
rect 230382 670692 230388 670744
rect 230440 670732 230446 670744
rect 580166 670732 580172 670744
rect 230440 670704 580172 670732
rect 230440 670692 230446 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 364334 656928 364340 656940
rect 3476 656900 364340 656928
rect 3476 656888 3482 656900
rect 364334 656888 364340 656900
rect 364392 656888 364398 656940
rect 220722 643084 220728 643136
rect 220780 643124 220786 643136
rect 580166 643124 580172 643136
rect 220780 643096 580172 643124
rect 220780 643084 220786 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 373994 632108 374000 632120
rect 3476 632080 374000 632108
rect 3476 632068 3482 632080
rect 373994 632068 374000 632080
rect 374052 632068 374058 632120
rect 224862 630640 224868 630692
rect 224920 630680 224926 630692
rect 580166 630680 580172 630692
rect 224920 630652 580172 630680
rect 224920 630640 224926 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 68278 618304 68284 618316
rect 3200 618276 68284 618304
rect 3200 618264 3206 618276
rect 68278 618264 68284 618276
rect 68336 618264 68342 618316
rect 216582 616836 216588 616888
rect 216640 616876 216646 616888
rect 580166 616876 580172 616888
rect 216640 616848 580172 616876
rect 216640 616836 216646 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 378134 605860 378140 605872
rect 3292 605832 378140 605860
rect 3292 605820 3298 605832
rect 378134 605820 378140 605832
rect 378192 605820 378198 605872
rect 208302 590656 208308 590708
rect 208360 590696 208366 590708
rect 579798 590696 579804 590708
rect 208360 590668 579804 590696
rect 208360 590656 208366 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 386414 579680 386420 579692
rect 3384 579652 386420 579680
rect 3384 579640 3390 579652
rect 386414 579640 386420 579652
rect 386472 579640 386478 579692
rect 212442 576852 212448 576904
rect 212500 576892 212506 576904
rect 580166 576892 580172 576904
rect 212500 576864 580172 576892
rect 212500 576852 212506 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 202782 563048 202788 563100
rect 202840 563088 202846 563100
rect 579798 563088 579804 563100
rect 202840 563060 579804 563088
rect 202840 563048 202846 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 391934 553432 391940 553444
rect 3476 553404 391940 553432
rect 3476 553392 3482 553404
rect 391934 553392 391940 553404
rect 391992 553392 391998 553444
rect 282270 551284 282276 551336
rect 282328 551324 282334 551336
rect 324958 551324 324964 551336
rect 282328 551296 324964 551324
rect 282328 551284 282334 551296
rect 324958 551284 324964 551296
rect 325016 551284 325022 551336
rect 268378 550536 268384 550588
rect 268436 550576 268442 550588
rect 329926 550576 329932 550588
rect 268436 550548 329932 550576
rect 268436 550536 268442 550548
rect 329926 550536 329932 550548
rect 329984 550536 329990 550588
rect 242158 550468 242164 550520
rect 242216 550508 242222 550520
rect 307938 550508 307944 550520
rect 242216 550480 307944 550508
rect 242216 550468 242222 550480
rect 307938 550468 307944 550480
rect 307996 550468 308002 550520
rect 255774 550400 255780 550452
rect 255832 550440 255838 550452
rect 331858 550440 331864 550452
rect 255832 550412 331864 550440
rect 255832 550400 255838 550412
rect 331858 550400 331864 550412
rect 331916 550400 331922 550452
rect 268930 550332 268936 550384
rect 268988 550372 268994 550384
rect 400858 550372 400864 550384
rect 268988 550344 400864 550372
rect 268988 550332 268994 550344
rect 400858 550332 400864 550344
rect 400916 550332 400922 550384
rect 180058 550264 180064 550316
rect 180116 550304 180122 550316
rect 321554 550304 321560 550316
rect 180116 550276 321560 550304
rect 180116 550264 180122 550276
rect 321554 550264 321560 550276
rect 321612 550264 321618 550316
rect 93118 550196 93124 550248
rect 93176 550236 93182 550248
rect 343174 550236 343180 550248
rect 93176 550208 343180 550236
rect 93176 550196 93182 550208
rect 343174 550196 343180 550208
rect 343232 550196 343238 550248
rect 65518 550128 65524 550180
rect 65576 550168 65582 550180
rect 356422 550168 356428 550180
rect 65576 550140 356428 550168
rect 65576 550128 65582 550140
rect 356422 550128 356428 550140
rect 356480 550128 356486 550180
rect 242526 550060 242532 550112
rect 242584 550100 242590 550112
rect 538858 550100 538864 550112
rect 242584 550072 538864 550100
rect 242584 550060 242590 550072
rect 538858 550060 538864 550072
rect 538916 550060 538922 550112
rect 61378 549992 61384 550044
rect 61436 550032 61442 550044
rect 370038 550032 370044 550044
rect 61436 550004 370044 550032
rect 61436 549992 61442 550004
rect 370038 549992 370044 550004
rect 370096 549992 370102 550044
rect 68278 549924 68284 549976
rect 68336 549964 68342 549976
rect 382826 549964 382832 549976
rect 68336 549936 382832 549964
rect 68336 549924 68342 549936
rect 382826 549924 382832 549936
rect 382884 549924 382890 549976
rect 3510 549856 3516 549908
rect 3568 549896 3574 549908
rect 396166 549896 396172 549908
rect 3568 549868 396172 549896
rect 3568 549856 3574 549868
rect 396166 549856 396172 549868
rect 396224 549856 396230 549908
rect 255958 549788 255964 549840
rect 256016 549828 256022 549840
rect 316770 549828 316776 549840
rect 256016 549800 316776 549828
rect 256016 549788 256022 549800
rect 316770 549788 316776 549800
rect 316828 549788 316834 549840
rect 295242 549720 295248 549772
rect 295300 549760 295306 549772
rect 299566 549760 299572 549772
rect 295300 549732 299572 549760
rect 295300 549720 295306 549732
rect 299566 549720 299572 549732
rect 299624 549720 299630 549772
rect 172054 549176 172060 549228
rect 172112 549216 172118 549228
rect 431310 549216 431316 549228
rect 172112 549188 431316 549216
rect 172112 549176 172118 549188
rect 431310 549176 431316 549188
rect 431368 549176 431374 549228
rect 198550 549108 198556 549160
rect 198608 549148 198614 549160
rect 554038 549148 554044 549160
rect 198608 549120 554044 549148
rect 198608 549108 198614 549120
rect 554038 549108 554044 549120
rect 554096 549108 554102 549160
rect 40862 549040 40868 549092
rect 40920 549080 40926 549092
rect 404814 549080 404820 549092
rect 40920 549052 404820 549080
rect 40920 549040 40926 549052
rect 404814 549040 404820 549052
rect 404872 549040 404878 549092
rect 180702 548972 180708 549024
rect 180760 549012 180766 549024
rect 565170 549012 565176 549024
rect 180760 548984 565176 549012
rect 180760 548972 180766 548984
rect 565170 548972 565176 548984
rect 565228 548972 565234 549024
rect 132402 548904 132408 548956
rect 132460 548944 132466 548956
rect 180794 548944 180800 548956
rect 132460 548916 180800 548944
rect 132460 548904 132466 548916
rect 180794 548904 180800 548916
rect 180852 548904 180858 548956
rect 185302 548904 185308 548956
rect 185360 548944 185366 548956
rect 576210 548944 576216 548956
rect 185360 548916 576216 548944
rect 185360 548904 185366 548916
rect 576210 548904 576216 548916
rect 576268 548904 576274 548956
rect 11790 548836 11796 548888
rect 11848 548876 11854 548888
rect 409230 548876 409236 548888
rect 11848 548848 409236 548876
rect 11848 548836 11854 548848
rect 409230 548836 409236 548848
rect 409288 548836 409294 548888
rect 167730 548768 167736 548820
rect 167788 548808 167794 548820
rect 574830 548808 574836 548820
rect 167788 548780 574836 548808
rect 167788 548768 167794 548780
rect 574830 548768 574836 548780
rect 574888 548768 574894 548820
rect 150066 548700 150072 548752
rect 150124 548740 150130 548752
rect 561030 548740 561036 548752
rect 150124 548712 561036 548740
rect 150124 548700 150130 548712
rect 561030 548700 561036 548712
rect 561088 548700 561094 548752
rect 154298 548632 154304 548684
rect 154356 548672 154362 548684
rect 573450 548672 573456 548684
rect 154356 548644 573456 548672
rect 154356 548632 154362 548644
rect 573450 548632 573456 548644
rect 573508 548632 573514 548684
rect 40678 548564 40684 548616
rect 40736 548604 40742 548616
rect 462498 548604 462504 548616
rect 40736 548576 462504 548604
rect 40736 548564 40742 548576
rect 462498 548564 462504 548576
rect 462556 548564 462562 548616
rect 17310 548496 17316 548548
rect 17368 548536 17374 548548
rect 448882 548536 448888 548548
rect 17368 548508 448888 548536
rect 17368 548496 17374 548508
rect 448882 548496 448888 548508
rect 448940 548496 448946 548548
rect 22738 548428 22744 548480
rect 22796 548468 22802 548480
rect 470870 548468 470876 548480
rect 22796 548440 470876 548468
rect 22796 548428 22802 548440
rect 470870 548428 470876 548440
rect 470928 548428 470934 548480
rect 471514 548428 471520 548480
rect 471572 548468 471578 548480
rect 541342 548468 541348 548480
rect 471572 548440 541348 548468
rect 471572 548428 471578 548440
rect 541342 548428 541348 548440
rect 541400 548428 541406 548480
rect 25590 548360 25596 548412
rect 25648 548400 25654 548412
rect 475286 548400 475292 548412
rect 25648 548372 475292 548400
rect 25648 548360 25654 548372
rect 475286 548360 475292 548372
rect 475344 548360 475350 548412
rect 29638 548292 29644 548344
rect 29696 548332 29702 548344
rect 488534 548332 488540 548344
rect 29696 548304 488540 548332
rect 29696 548292 29702 548304
rect 488534 548292 488540 548304
rect 488592 548292 488598 548344
rect 101674 548224 101680 548276
rect 101732 548264 101738 548276
rect 562318 548264 562324 548276
rect 101732 548236 562324 548264
rect 101732 548224 101738 548236
rect 562318 548224 562324 548236
rect 562376 548224 562382 548276
rect 15930 548156 15936 548208
rect 15988 548196 15994 548208
rect 484394 548196 484400 548208
rect 15988 548168 484400 548196
rect 15988 548156 15994 548168
rect 484394 548156 484400 548168
rect 484452 548156 484458 548208
rect 32398 548088 32404 548140
rect 32456 548128 32462 548140
rect 501690 548128 501696 548140
rect 32456 548100 501696 548128
rect 32456 548088 32462 548100
rect 501690 548088 501696 548100
rect 501748 548088 501754 548140
rect 17218 548020 17224 548072
rect 17276 548060 17282 548072
rect 497274 548060 497280 548072
rect 17276 548032 497280 548060
rect 17276 548020 17282 548032
rect 497274 548020 497280 548032
rect 497332 548020 497338 548072
rect 75270 547952 75276 548004
rect 75328 547992 75334 548004
rect 558178 547992 558184 548004
rect 75328 547964 558184 547992
rect 75328 547952 75334 547964
rect 558178 547952 558184 547964
rect 558236 547952 558242 548004
rect 25498 547884 25504 547936
rect 25556 547924 25562 547936
rect 514846 547924 514852 547936
rect 25556 547896 514852 547924
rect 25556 547884 25562 547896
rect 514846 547884 514852 547896
rect 514904 547884 514910 547936
rect 189718 547748 189724 547800
rect 189776 547788 189782 547800
rect 548610 547788 548616 547800
rect 189776 547760 548616 547788
rect 189776 547748 189782 547760
rect 548610 547748 548616 547760
rect 548668 547748 548674 547800
rect 35250 547680 35256 547732
rect 35308 547720 35314 547732
rect 414106 547720 414112 547732
rect 35308 547692 414112 547720
rect 35308 547680 35314 547692
rect 414106 547680 414112 547692
rect 414164 547680 414170 547732
rect 36630 547612 36636 547664
rect 36688 547652 36694 547664
rect 426802 547652 426808 547664
rect 36688 547624 426808 547652
rect 36688 547612 36694 547624
rect 426802 547612 426808 547624
rect 426860 547612 426866 547664
rect 35158 547544 35164 547596
rect 35216 547584 35222 547596
rect 431218 547584 431224 547596
rect 35216 547556 431224 547584
rect 35216 547544 35222 547556
rect 431218 547544 431224 547556
rect 431276 547544 431282 547596
rect 431310 547544 431316 547596
rect 431368 547584 431374 547596
rect 580442 547584 580448 547596
rect 431368 547556 580448 547584
rect 431368 547544 431374 547556
rect 580442 547544 580448 547556
rect 580500 547544 580506 547596
rect 39390 547476 39396 547528
rect 39448 547516 39454 547528
rect 440234 547516 440240 547528
rect 39448 547488 440240 547516
rect 39448 547476 39454 547488
rect 440234 547476 440240 547488
rect 440292 547476 440298 547528
rect 39298 547408 39304 547460
rect 39356 547448 39362 547460
rect 457622 547448 457628 547460
rect 39356 547420 457628 547448
rect 39356 547408 39362 547420
rect 457622 547408 457628 547420
rect 457680 547408 457686 547460
rect 33778 547340 33784 547392
rect 33836 547380 33842 547392
rect 453206 547380 453212 547392
rect 33836 547352 453212 547380
rect 33836 547340 33842 547352
rect 453206 547340 453212 547352
rect 453264 547340 453270 547392
rect 136910 547272 136916 547324
rect 136968 547312 136974 547324
rect 558270 547312 558276 547324
rect 136968 547284 558276 547312
rect 136968 547272 136974 547284
rect 558270 547272 558276 547284
rect 558328 547272 558334 547324
rect 123662 547204 123668 547256
rect 123720 547244 123726 547256
rect 556890 547244 556896 547256
rect 123720 547216 556896 547244
rect 123720 547204 123726 547216
rect 556890 547204 556896 547216
rect 556948 547204 556954 547256
rect 110322 547136 110328 547188
rect 110380 547176 110386 547188
rect 555510 547176 555516 547188
rect 110380 547148 555516 547176
rect 110380 547136 110386 547148
rect 555510 547136 555516 547148
rect 555568 547136 555574 547188
rect 97258 547068 97264 547120
rect 97316 547108 97322 547120
rect 551370 547108 551376 547120
rect 97316 547080 551376 547108
rect 97316 547068 97322 547080
rect 551370 547068 551376 547080
rect 551428 547068 551434 547120
rect 83918 547000 83924 547052
rect 83976 547040 83982 547052
rect 544378 547040 544384 547052
rect 83976 547012 544384 547040
rect 83976 547000 83982 547012
rect 544378 547000 544384 547012
rect 544436 547000 544442 547052
rect 4890 546932 4896 546984
rect 4948 546972 4954 546984
rect 466454 546972 466460 546984
rect 4948 546944 466460 546972
rect 4948 546932 4954 546944
rect 466454 546932 466460 546944
rect 466512 546932 466518 546984
rect 7650 546864 7656 546916
rect 7708 546904 7714 546916
rect 479702 546904 479708 546916
rect 7708 546876 479708 546904
rect 7708 546864 7714 546876
rect 479702 546864 479708 546876
rect 479760 546864 479766 546916
rect 88242 546796 88248 546848
rect 88300 546836 88306 546848
rect 560938 546836 560944 546848
rect 88300 546808 560944 546836
rect 88300 546796 88306 546808
rect 560938 546796 560944 546808
rect 560996 546796 561002 546848
rect 70854 546728 70860 546780
rect 70912 546768 70918 546780
rect 548518 546768 548524 546780
rect 70912 546740 548524 546768
rect 70912 546728 70918 546740
rect 548518 546728 548524 546740
rect 548576 546728 548582 546780
rect 11698 546660 11704 546712
rect 11756 546700 11762 546712
rect 492858 546700 492864 546712
rect 11756 546672 492864 546700
rect 11756 546660 11762 546672
rect 492858 546660 492864 546672
rect 492916 546660 492922 546712
rect 21358 546592 21364 546644
rect 21416 546632 21422 546644
rect 506566 546632 506572 546644
rect 21416 546604 506572 546632
rect 21416 546592 21422 546604
rect 506566 546592 506572 546604
rect 506624 546592 506630 546644
rect 62022 546524 62028 546576
rect 62080 546564 62086 546576
rect 556798 546564 556804 546576
rect 62080 546536 556804 546564
rect 62080 546524 62086 546536
rect 556798 546524 556804 546536
rect 556856 546524 556862 546576
rect 4798 546456 4804 546508
rect 4856 546496 4862 546508
rect 519262 546496 519268 546508
rect 4856 546468 519268 546496
rect 4856 546456 4862 546468
rect 519262 546456 519268 546468
rect 519320 546456 519326 546508
rect 180794 546388 180800 546440
rect 180852 546428 180858 546440
rect 580258 546428 580264 546440
rect 180852 546400 580264 546428
rect 180852 546388 180858 546400
rect 580258 546388 580264 546400
rect 580316 546388 580322 546440
rect 194134 546320 194140 546372
rect 194192 546360 194198 546372
rect 544470 546360 544476 546372
rect 194192 546332 544476 546360
rect 194192 546320 194198 546332
rect 544470 546320 544476 546332
rect 544528 546320 544534 546372
rect 33870 546252 33876 546304
rect 33928 546292 33934 546304
rect 400398 546292 400404 546304
rect 33928 546264 400404 546292
rect 33928 546252 33934 546264
rect 400398 546252 400404 546264
rect 400456 546252 400462 546304
rect 176148 546184 176154 546236
rect 176206 546224 176212 546236
rect 545850 546224 545856 546236
rect 176206 546196 545856 546224
rect 176206 546184 176212 546196
rect 545850 546184 545856 546196
rect 545908 546184 545914 546236
rect 40770 546116 40776 546168
rect 40828 546156 40834 546168
rect 418154 546156 418160 546168
rect 40828 546128 418160 546156
rect 40828 546116 40834 546128
rect 418154 546116 418160 546128
rect 418212 546116 418218 546168
rect 163314 546048 163320 546100
rect 163372 546088 163378 546100
rect 562410 546088 562416 546100
rect 163372 546060 562416 546088
rect 163372 546048 163378 546060
rect 562410 546048 562416 546060
rect 562468 546048 562474 546100
rect 145650 545980 145656 546032
rect 145708 546020 145714 546032
rect 547230 546020 547236 546032
rect 145708 545992 547236 546020
rect 145708 545980 145714 545992
rect 547230 545980 547236 545992
rect 547288 545980 547294 546032
rect 36538 545912 36544 545964
rect 36596 545952 36602 545964
rect 444466 545952 444472 545964
rect 36596 545924 444472 545952
rect 36596 545912 36602 545924
rect 444466 545912 444472 545924
rect 444524 545912 444530 545964
rect 10318 545844 10324 545896
rect 10376 545884 10382 545896
rect 422478 545884 422484 545896
rect 10376 545856 422484 545884
rect 10376 545844 10382 545856
rect 422478 545844 422484 545856
rect 422536 545844 422542 545896
rect 14550 545776 14556 545828
rect 14608 545816 14614 545828
rect 435634 545816 435640 545828
rect 14608 545788 435640 545816
rect 14608 545776 14614 545788
rect 435634 545776 435640 545788
rect 435692 545776 435698 545828
rect 158714 545708 158720 545760
rect 158772 545748 158778 545760
rect 580350 545748 580356 545760
rect 158772 545720 580356 545748
rect 158772 545708 158778 545720
rect 580350 545708 580356 545720
rect 580408 545708 580414 545760
rect 141234 545640 141240 545692
rect 141292 545680 141298 545692
rect 569310 545680 569316 545692
rect 141292 545652 569316 545680
rect 141292 545640 141298 545652
rect 569310 545640 569316 545652
rect 569368 545640 569374 545692
rect 128078 545572 128084 545624
rect 128136 545612 128142 545624
rect 566550 545612 566556 545624
rect 128136 545584 566556 545612
rect 128136 545572 128142 545584
rect 566550 545572 566556 545584
rect 566608 545572 566614 545624
rect 114830 545504 114836 545556
rect 114888 545544 114894 545556
rect 565078 545544 565084 545556
rect 114888 545516 565084 545544
rect 114888 545504 114894 545516
rect 565078 545504 565084 545516
rect 565136 545504 565142 545556
rect 64846 545448 74534 545476
rect 57606 545368 57612 545420
rect 57664 545408 57670 545420
rect 64846 545408 64874 545448
rect 57664 545380 64874 545408
rect 57664 545368 57670 545380
rect 66254 545368 66260 545420
rect 66312 545368 66318 545420
rect 66272 545340 66300 545368
rect 66272 545312 70348 545340
rect 70320 545136 70348 545312
rect 74506 545272 74534 545448
rect 119246 545436 119252 545488
rect 119304 545476 119310 545488
rect 576118 545476 576124 545488
rect 119304 545448 576124 545476
rect 119304 545436 119310 545448
rect 576118 545436 576124 545448
rect 576176 545436 576182 545488
rect 79594 545368 79600 545420
rect 79652 545408 79658 545420
rect 84289 545411 84347 545417
rect 84289 545408 84301 545411
rect 79652 545380 84301 545408
rect 79652 545368 79658 545380
rect 84289 545377 84301 545380
rect 84335 545377 84347 545411
rect 84289 545371 84347 545377
rect 92842 545368 92848 545420
rect 92900 545368 92906 545420
rect 106090 545368 106096 545420
rect 106148 545408 106154 545420
rect 574738 545408 574744 545420
rect 106148 545380 574744 545408
rect 106148 545368 106154 545380
rect 574738 545368 574744 545380
rect 574796 545368 574802 545420
rect 92860 545340 92888 545368
rect 573358 545340 573364 545352
rect 92860 545312 573364 545340
rect 573358 545300 573364 545312
rect 573416 545300 573422 545352
rect 545758 545272 545764 545284
rect 74506 545244 545764 545272
rect 545758 545232 545764 545244
rect 545816 545232 545822 545284
rect 84289 545207 84347 545213
rect 84289 545173 84301 545207
rect 84335 545204 84347 545207
rect 569218 545204 569224 545216
rect 84335 545176 569224 545204
rect 84335 545173 84347 545176
rect 84289 545167 84347 545173
rect 569218 545164 569224 545176
rect 569276 545164 569282 545216
rect 566458 545136 566464 545148
rect 70320 545108 566464 545136
rect 566458 545096 566464 545108
rect 566516 545096 566522 545148
rect 544470 538160 544476 538212
rect 544528 538200 544534 538212
rect 580166 538200 580172 538212
rect 544528 538172 580172 538200
rect 544528 538160 544534 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 3326 528504 3332 528556
rect 3384 528544 3390 528556
rect 33870 528544 33876 528556
rect 3384 528516 33876 528544
rect 3384 528504 3390 528516
rect 33870 528504 33876 528516
rect 33928 528504 33934 528556
rect 554038 525716 554044 525768
rect 554096 525756 554102 525768
rect 580166 525756 580172 525768
rect 554096 525728 580172 525756
rect 554096 525716 554102 525728
rect 580166 525716 580172 525728
rect 580224 525716 580230 525768
rect 3142 516060 3148 516112
rect 3200 516100 3206 516112
rect 11790 516100 11796 516112
rect 3200 516072 11796 516100
rect 3200 516060 3206 516072
rect 11790 516060 11796 516072
rect 11848 516060 11854 516112
rect 548610 511912 548616 511964
rect 548668 511952 548674 511964
rect 580166 511952 580172 511964
rect 548668 511924 580172 511952
rect 548668 511912 548674 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 2958 502256 2964 502308
rect 3016 502296 3022 502308
rect 40862 502296 40868 502308
rect 3016 502268 40868 502296
rect 3016 502256 3022 502268
rect 40862 502256 40868 502268
rect 40920 502256 40926 502308
rect 565170 485732 565176 485784
rect 565228 485772 565234 485784
rect 580166 485772 580172 485784
rect 565228 485744 580172 485772
rect 565228 485732 565234 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 3234 476008 3240 476060
rect 3292 476048 3298 476060
rect 35250 476048 35256 476060
rect 3292 476020 35256 476048
rect 3292 476008 3298 476020
rect 35250 476008 35256 476020
rect 35308 476008 35314 476060
rect 576210 471928 576216 471980
rect 576268 471968 576274 471980
rect 580166 471968 580172 471980
rect 576268 471940 580172 471968
rect 576268 471928 576274 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 3050 463632 3056 463684
rect 3108 463672 3114 463684
rect 10318 463672 10324 463684
rect 3108 463644 10324 463672
rect 3108 463632 3114 463644
rect 10318 463632 10324 463644
rect 10376 463632 10382 463684
rect 545850 458124 545856 458176
rect 545908 458164 545914 458176
rect 580166 458164 580172 458176
rect 545908 458136 580172 458164
rect 545908 458124 545914 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 40770 449868 40776 449880
rect 3384 449840 40776 449868
rect 3384 449828 3390 449840
rect 40770 449828 40776 449840
rect 40828 449828 40834 449880
rect 574830 431876 574836 431928
rect 574888 431916 574894 431928
rect 580166 431916 580172 431928
rect 574888 431888 580172 431916
rect 574888 431876 574894 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 36630 423620 36636 423632
rect 3384 423592 36636 423620
rect 3384 423580 3390 423592
rect 36630 423580 36636 423592
rect 36688 423580 36694 423632
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 14550 411244 14556 411256
rect 3016 411216 14556 411244
rect 3016 411204 3022 411216
rect 14550 411204 14556 411216
rect 14608 411204 14614 411256
rect 562410 405628 562416 405680
rect 562468 405668 562474 405680
rect 580166 405668 580172 405680
rect 562468 405640 580172 405668
rect 562468 405628 562474 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 35158 398800 35164 398812
rect 3384 398772 35164 398800
rect 3384 398760 3390 398772
rect 35158 398760 35164 398772
rect 35216 398760 35222 398812
rect 573450 379448 573456 379500
rect 573508 379488 573514 379500
rect 580166 379488 580172 379500
rect 573508 379460 580172 379488
rect 573508 379448 573514 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 39390 372552 39396 372564
rect 3384 372524 39396 372552
rect 3384 372512 3390 372524
rect 39390 372512 39396 372524
rect 39448 372512 39454 372564
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 17310 358748 17316 358760
rect 3384 358720 17316 358748
rect 3384 358708 3390 358720
rect 17310 358708 17316 358720
rect 17368 358708 17374 358760
rect 561030 353200 561036 353252
rect 561088 353240 561094 353252
rect 580166 353240 580172 353252
rect 561088 353212 580172 353240
rect 561088 353200 561094 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 36538 346372 36544 346384
rect 3384 346344 36544 346372
rect 3384 346332 3390 346344
rect 36538 346332 36544 346344
rect 36596 346332 36602 346384
rect 569310 325592 569316 325644
rect 569368 325632 569374 325644
rect 579890 325632 579896 325644
rect 569368 325604 579896 325632
rect 569368 325592 569374 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 33778 320124 33784 320136
rect 3384 320096 33784 320124
rect 3384 320084 3390 320096
rect 33778 320084 33784 320096
rect 33836 320084 33842 320136
rect 547230 313216 547236 313268
rect 547288 313256 547294 313268
rect 580166 313256 580172 313268
rect 547288 313228 580172 313256
rect 547288 313216 547294 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 40678 306320 40684 306332
rect 3384 306292 40684 306320
rect 3384 306280 3390 306292
rect 40678 306280 40684 306292
rect 40736 306280 40742 306332
rect 558270 299412 558276 299464
rect 558328 299452 558334 299464
rect 579614 299452 579620 299464
rect 558328 299424 579620 299452
rect 558328 299412 558334 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 3326 293904 3332 293956
rect 3384 293944 3390 293956
rect 39298 293944 39304 293956
rect 3384 293916 39304 293944
rect 3384 293904 3390 293916
rect 39298 293904 39304 293916
rect 39356 293904 39362 293956
rect 566550 273164 566556 273216
rect 566608 273204 566614 273216
rect 579890 273204 579896 273216
rect 566608 273176 579896 273204
rect 566608 273164 566614 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 2774 267248 2780 267300
rect 2832 267288 2838 267300
rect 4890 267288 4896 267300
rect 2832 267260 4896 267288
rect 2832 267248 2838 267260
rect 4890 267248 4896 267260
rect 4948 267248 4954 267300
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 25590 255252 25596 255264
rect 3200 255224 25596 255252
rect 3200 255212 3206 255224
rect 25590 255212 25596 255224
rect 25648 255212 25654 255264
rect 556890 245556 556896 245608
rect 556948 245596 556954 245608
rect 580166 245596 580172 245608
rect 556948 245568 580172 245596
rect 556948 245556 556954 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 22738 241448 22744 241460
rect 3292 241420 22744 241448
rect 3292 241408 3298 241420
rect 22738 241408 22744 241420
rect 22796 241408 22802 241460
rect 565078 233180 565084 233232
rect 565136 233220 565142 233232
rect 579982 233220 579988 233232
rect 565136 233192 579988 233220
rect 565136 233180 565142 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 576118 219376 576124 219428
rect 576176 219416 576182 219428
rect 580166 219416 580172 219428
rect 576176 219388 580172 219416
rect 576176 219376 576182 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3326 214956 3332 215008
rect 3384 214996 3390 215008
rect 7650 214996 7656 215008
rect 3384 214968 7656 214996
rect 3384 214956 3390 214968
rect 7650 214956 7656 214968
rect 7708 214956 7714 215008
rect 555510 206932 555516 206984
rect 555568 206972 555574 206984
rect 579798 206972 579804 206984
rect 555568 206944 579804 206972
rect 555568 206932 555574 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 29638 202824 29644 202836
rect 3108 202796 29644 202824
rect 3108 202784 3114 202796
rect 29638 202784 29644 202796
rect 29696 202784 29702 202836
rect 562318 193128 562324 193180
rect 562376 193168 562382 193180
rect 580166 193168 580172 193180
rect 562376 193140 580172 193168
rect 562376 193128 562382 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 15930 189020 15936 189032
rect 3200 188992 15936 189020
rect 3200 188980 3206 188992
rect 15930 188980 15936 188992
rect 15988 188980 15994 189032
rect 574738 179324 574744 179376
rect 574796 179364 574802 179376
rect 580166 179364 580172 179376
rect 574796 179336 580172 179364
rect 574796 179324 574802 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 551370 166948 551376 167000
rect 551428 166988 551434 167000
rect 580166 166988 580172 167000
rect 551428 166960 580172 166988
rect 551428 166948 551434 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 11698 164200 11704 164212
rect 3384 164172 11704 164200
rect 3384 164160 3390 164172
rect 11698 164160 11704 164172
rect 11756 164160 11762 164212
rect 560938 153144 560944 153196
rect 560996 153184 561002 153196
rect 580166 153184 580172 153196
rect 560996 153156 580172 153184
rect 560996 153144 561002 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3602 150356 3608 150408
rect 3660 150396 3666 150408
rect 32398 150396 32404 150408
rect 3660 150368 32404 150396
rect 3660 150356 3666 150368
rect 32398 150356 32404 150368
rect 32456 150356 32462 150408
rect 573358 139340 573364 139392
rect 573416 139380 573422 139392
rect 580166 139380 580172 139392
rect 573416 139352 580172 139380
rect 573416 139340 573422 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3326 137912 3332 137964
rect 3384 137952 3390 137964
rect 17218 137952 17224 137964
rect 3384 137924 17224 137952
rect 3384 137912 3390 137924
rect 17218 137912 17224 137924
rect 17276 137912 17282 137964
rect 544378 126896 544384 126948
rect 544436 126936 544442 126948
rect 580166 126936 580172 126948
rect 544436 126908 580172 126936
rect 544436 126896 544442 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 558178 113092 558184 113144
rect 558236 113132 558242 113144
rect 579798 113132 579804 113144
rect 558236 113104 579804 113132
rect 558236 113092 558242 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 21358 111772 21364 111784
rect 3200 111744 21364 111772
rect 3200 111732 3206 111744
rect 21358 111732 21364 111744
rect 21416 111732 21422 111784
rect 569218 100648 569224 100700
rect 569276 100688 569282 100700
rect 580166 100688 580172 100700
rect 569276 100660 580172 100688
rect 569276 100648 569282 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3234 97928 3240 97980
rect 3292 97968 3298 97980
rect 25498 97968 25504 97980
rect 3292 97940 25504 97968
rect 3292 97928 3298 97940
rect 25498 97928 25504 97940
rect 25556 97928 25562 97980
rect 548518 86912 548524 86964
rect 548576 86952 548582 86964
rect 580166 86952 580172 86964
rect 548576 86924 580172 86952
rect 548576 86912 548582 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3326 85484 3332 85536
rect 3384 85524 3390 85536
rect 18598 85524 18604 85536
rect 3384 85496 18604 85524
rect 3384 85484 3390 85496
rect 18598 85484 18604 85496
rect 18656 85484 18662 85536
rect 556798 73108 556804 73160
rect 556856 73148 556862 73160
rect 580166 73148 580172 73160
rect 556856 73120 580172 73148
rect 556856 73108 556862 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 2774 71612 2780 71664
rect 2832 71652 2838 71664
rect 4798 71652 4804 71664
rect 2832 71624 4804 71652
rect 2832 71612 2838 71624
rect 4798 71612 4804 71624
rect 4856 71612 4862 71664
rect 566458 60664 566464 60716
rect 566516 60704 566522 60716
rect 580166 60704 580172 60716
rect 566516 60676 580172 60704
rect 566516 60664 566522 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 545758 46860 545764 46912
rect 545816 46900 545822 46912
rect 580166 46900 580172 46912
rect 545816 46872 580172 46900
rect 545816 46860 545822 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 7558 45540 7564 45552
rect 3568 45512 7564 45540
rect 3568 45500 3574 45512
rect 7558 45500 7564 45512
rect 7616 45500 7622 45552
rect 133966 41828 133972 41880
rect 134024 41868 134030 41880
rect 135116 41868 135122 41880
rect 134024 41840 135122 41868
rect 134024 41828 134030 41840
rect 135116 41828 135122 41840
rect 135174 41828 135180 41880
rect 179984 40072 181024 40100
rect 20622 39992 20628 40044
rect 20680 40032 20686 40044
rect 58710 40032 58716 40044
rect 20680 40004 58716 40032
rect 20680 39992 20686 40004
rect 58710 39992 58716 40004
rect 58768 39992 58774 40044
rect 75822 39992 75828 40044
rect 75880 40032 75886 40044
rect 106550 40032 106556 40044
rect 75880 40004 106556 40032
rect 75880 39992 75886 40004
rect 106550 39992 106556 40004
rect 106608 39992 106614 40044
rect 110322 39992 110328 40044
rect 110380 40032 110386 40044
rect 136082 40032 136088 40044
rect 110380 40004 136088 40032
rect 110380 39992 110386 40004
rect 136082 39992 136088 40004
rect 136140 39992 136146 40044
rect 136542 39992 136548 40044
rect 136600 40032 136606 40044
rect 158438 40032 158444 40044
rect 136600 40004 158444 40032
rect 136600 39992 136606 40004
rect 158438 39992 158444 40004
rect 158496 39992 158502 40044
rect 158622 39992 158628 40044
rect 158680 40032 158686 40044
rect 177758 40032 177764 40044
rect 158680 40004 177764 40032
rect 158680 39992 158686 40004
rect 177758 39992 177764 40004
rect 177816 39992 177822 40044
rect 177942 39992 177948 40044
rect 178000 40032 178006 40044
rect 179984 40032 180012 40072
rect 178000 40004 180012 40032
rect 178000 39992 178006 40004
rect 180058 39992 180064 40044
rect 180116 40032 180122 40044
rect 180886 40032 180892 40044
rect 180116 40004 180892 40032
rect 180116 39992 180122 40004
rect 180886 39992 180892 40004
rect 180944 39992 180950 40044
rect 180996 40032 181024 40072
rect 195146 40032 195152 40044
rect 180996 40004 195152 40032
rect 195146 39992 195152 40004
rect 195204 39992 195210 40044
rect 200022 39992 200028 40044
rect 200080 40032 200086 40044
rect 213454 40032 213460 40044
rect 200080 40004 213460 40032
rect 200080 39992 200086 40004
rect 213454 39992 213460 40004
rect 213512 39992 213518 40044
rect 223482 39992 223488 40044
rect 223540 40032 223546 40044
rect 233786 40032 233792 40044
rect 223540 40004 233792 40032
rect 223540 39992 223546 40004
rect 233786 39992 233792 40004
rect 233844 39992 233850 40044
rect 242802 39992 242808 40044
rect 242860 40032 242866 40044
rect 250070 40032 250076 40044
rect 242860 40004 250076 40032
rect 242860 39992 242866 40004
rect 250070 39992 250076 40004
rect 250128 39992 250134 40044
rect 253842 39992 253848 40044
rect 253900 40032 253906 40044
rect 260282 40032 260288 40044
rect 253900 40004 260288 40032
rect 253900 39992 253906 40004
rect 260282 39992 260288 40004
rect 260340 39992 260346 40044
rect 277302 39992 277308 40044
rect 277360 40032 277366 40044
rect 279602 40032 279608 40044
rect 277360 40004 279608 40032
rect 277360 39992 277366 40004
rect 279602 39992 279608 40004
rect 279660 39992 279666 40044
rect 286962 39992 286968 40044
rect 287020 40032 287026 40044
rect 288802 40032 288808 40044
rect 287020 40004 288808 40032
rect 287020 39992 287026 40004
rect 288802 39992 288808 40004
rect 288860 39992 288866 40044
rect 315298 39992 315304 40044
rect 315356 40032 315362 40044
rect 316126 40032 316132 40044
rect 315356 40004 316132 40032
rect 315356 39992 315362 40004
rect 316126 39992 316132 40004
rect 316184 39992 316190 40044
rect 509786 39992 509792 40044
rect 509844 40032 509850 40044
rect 515493 40035 515551 40041
rect 515493 40032 515505 40035
rect 509844 40004 515505 40032
rect 509844 39992 509850 40004
rect 515493 40001 515505 40004
rect 515539 40001 515551 40035
rect 515493 39995 515551 40001
rect 538306 39992 538312 40044
rect 538364 40032 538370 40044
rect 565078 40032 565084 40044
rect 538364 40004 565084 40032
rect 538364 39992 538370 40004
rect 565078 39992 565084 40004
rect 565136 39992 565142 40044
rect 26142 39924 26148 39976
rect 26200 39964 26206 39976
rect 63770 39964 63776 39976
rect 26200 39936 63776 39964
rect 26200 39924 26206 39936
rect 63770 39924 63776 39936
rect 63828 39924 63834 39976
rect 74442 39924 74448 39976
rect 74500 39964 74506 39976
rect 105538 39964 105544 39976
rect 74500 39936 105544 39964
rect 74500 39924 74506 39936
rect 105538 39924 105544 39936
rect 105596 39924 105602 39976
rect 107562 39924 107568 39976
rect 107620 39964 107626 39976
rect 134058 39964 134064 39976
rect 107620 39936 134064 39964
rect 107620 39924 107626 39936
rect 134058 39924 134064 39936
rect 134116 39924 134122 39976
rect 144822 39924 144828 39976
rect 144880 39964 144886 39976
rect 166626 39964 166632 39976
rect 144880 39936 166632 39964
rect 144880 39924 144886 39936
rect 166626 39924 166632 39936
rect 166684 39924 166690 39976
rect 169570 39924 169576 39976
rect 169628 39964 169634 39976
rect 186958 39964 186964 39976
rect 169628 39936 186964 39964
rect 169628 39924 169634 39936
rect 186958 39924 186964 39936
rect 187016 39924 187022 39976
rect 190362 39924 190368 39976
rect 190420 39964 190426 39976
rect 205266 39964 205272 39976
rect 190420 39936 205272 39964
rect 190420 39924 190426 39936
rect 205266 39924 205272 39936
rect 205324 39924 205330 39976
rect 205542 39924 205548 39976
rect 205600 39964 205606 39976
rect 218514 39964 218520 39976
rect 205600 39936 218520 39964
rect 205600 39924 205606 39936
rect 218514 39924 218520 39936
rect 218572 39924 218578 39976
rect 222102 39924 222108 39976
rect 222160 39964 222166 39976
rect 232774 39964 232780 39976
rect 222160 39936 232780 39964
rect 222160 39924 222166 39936
rect 232774 39924 232780 39936
rect 232832 39924 232838 39976
rect 275922 39924 275928 39976
rect 275980 39964 275986 39976
rect 278590 39964 278596 39976
rect 275980 39936 278596 39964
rect 275980 39924 275986 39936
rect 278590 39924 278596 39936
rect 278648 39924 278654 39976
rect 285582 39924 285588 39976
rect 285640 39964 285646 39976
rect 287790 39964 287796 39976
rect 285640 39936 287796 39964
rect 285640 39924 285646 39936
rect 287790 39924 287796 39936
rect 287848 39924 287854 39976
rect 495526 39924 495532 39976
rect 495584 39964 495590 39976
rect 495584 39936 509234 39964
rect 495584 39924 495590 39936
rect 23382 39856 23388 39908
rect 23440 39896 23446 39908
rect 61746 39896 61752 39908
rect 23440 39868 61752 39896
rect 23440 39856 23446 39868
rect 61746 39856 61752 39868
rect 61804 39856 61810 39908
rect 68922 39856 68928 39908
rect 68980 39896 68986 39908
rect 100386 39896 100392 39908
rect 68980 39868 100392 39896
rect 68980 39856 68986 39868
rect 100386 39856 100392 39868
rect 100444 39856 100450 39908
rect 103422 39856 103428 39908
rect 103480 39896 103486 39908
rect 129918 39896 129924 39908
rect 103480 39868 129924 39896
rect 103480 39856 103486 39868
rect 129918 39856 129924 39868
rect 129976 39856 129982 39908
rect 142062 39856 142068 39908
rect 142120 39896 142126 39908
rect 163498 39896 163504 39908
rect 142120 39868 163504 39896
rect 142120 39856 142126 39868
rect 163498 39856 163504 39868
rect 163556 39856 163562 39908
rect 165522 39856 165528 39908
rect 165580 39896 165586 39908
rect 183922 39896 183928 39908
rect 165580 39868 183928 39896
rect 165580 39856 165586 39868
rect 183922 39856 183928 39868
rect 183980 39856 183986 39908
rect 187602 39856 187608 39908
rect 187660 39896 187666 39908
rect 203242 39896 203248 39908
rect 187660 39868 203248 39896
rect 187660 39856 187666 39868
rect 203242 39856 203248 39868
rect 203300 39856 203306 39908
rect 204162 39856 204168 39908
rect 204220 39896 204226 39908
rect 217502 39896 217508 39908
rect 204220 39868 217508 39896
rect 204220 39856 204226 39868
rect 217502 39856 217508 39868
rect 217560 39856 217566 39908
rect 217962 39856 217968 39908
rect 218020 39896 218026 39908
rect 228726 39896 228732 39908
rect 218020 39868 228732 39896
rect 218020 39856 218026 39868
rect 228726 39856 228732 39868
rect 228784 39856 228790 39908
rect 235902 39856 235908 39908
rect 235960 39896 235966 39908
rect 243998 39896 244004 39908
rect 235960 39868 244004 39896
rect 235960 39856 235966 39868
rect 243998 39856 244004 39868
rect 244056 39856 244062 39908
rect 509206 39896 509234 39936
rect 513834 39924 513840 39976
rect 513892 39964 513898 39976
rect 524966 39964 524972 39976
rect 513892 39936 524972 39964
rect 513892 39924 513898 39936
rect 524966 39924 524972 39936
rect 525024 39924 525030 39976
rect 532234 39924 532240 39976
rect 532292 39964 532298 39976
rect 560938 39964 560944 39976
rect 532292 39936 560944 39964
rect 532292 39924 532298 39936
rect 560938 39924 560944 39936
rect 560996 39924 561002 39976
rect 515398 39896 515404 39908
rect 509206 39868 515404 39896
rect 515398 39856 515404 39868
rect 515456 39856 515462 39908
rect 515493 39899 515551 39905
rect 515493 39865 515505 39899
rect 515539 39896 515551 39899
rect 540422 39896 540428 39908
rect 515539 39868 540428 39896
rect 515539 39865 515551 39868
rect 515493 39859 515551 39865
rect 540422 39856 540428 39868
rect 540480 39856 540486 39908
rect 542354 39856 542360 39908
rect 542412 39896 542418 39908
rect 548610 39896 548616 39908
rect 542412 39868 548616 39896
rect 542412 39856 542418 39868
rect 548610 39856 548616 39868
rect 548668 39856 548674 39908
rect 19242 39788 19248 39840
rect 19300 39828 19306 39840
rect 57698 39828 57704 39840
rect 19300 39800 57704 39828
rect 19300 39788 19306 39800
rect 57698 39788 57704 39800
rect 57756 39788 57762 39840
rect 60642 39788 60648 39840
rect 60700 39828 60706 39840
rect 93302 39828 93308 39840
rect 60700 39800 93308 39828
rect 60700 39788 60706 39800
rect 93302 39788 93308 39800
rect 93360 39788 93366 39840
rect 95142 39788 95148 39840
rect 95200 39828 95206 39840
rect 123846 39828 123852 39840
rect 95200 39800 123852 39828
rect 95200 39788 95206 39800
rect 123846 39788 123852 39800
rect 123904 39788 123910 39840
rect 124122 39788 124128 39840
rect 124180 39828 124186 39840
rect 148226 39828 148232 39840
rect 124180 39800 148232 39828
rect 124180 39788 124186 39800
rect 148226 39788 148232 39800
rect 148284 39788 148290 39840
rect 153010 39788 153016 39840
rect 153068 39828 153074 39840
rect 173710 39828 173716 39840
rect 153068 39800 173716 39828
rect 153068 39788 153074 39800
rect 173710 39788 173716 39800
rect 173768 39788 173774 39840
rect 173802 39788 173808 39840
rect 173860 39828 173866 39840
rect 191006 39828 191012 39840
rect 173860 39800 191012 39828
rect 173860 39788 173866 39800
rect 191006 39788 191012 39800
rect 191064 39788 191070 39840
rect 195882 39788 195888 39840
rect 195940 39828 195946 39840
rect 210418 39828 210424 39840
rect 195940 39800 210424 39828
rect 195940 39788 195946 39800
rect 210418 39788 210424 39800
rect 210476 39788 210482 39840
rect 211062 39788 211068 39840
rect 211120 39828 211126 39840
rect 222562 39828 222568 39840
rect 211120 39800 222568 39828
rect 211120 39788 211126 39800
rect 222562 39788 222568 39800
rect 222620 39788 222626 39840
rect 224862 39788 224868 39840
rect 224920 39828 224926 39840
rect 234798 39828 234804 39840
rect 224920 39800 234804 39828
rect 224920 39788 224926 39800
rect 234798 39788 234804 39800
rect 234856 39788 234862 39840
rect 237282 39788 237288 39840
rect 237340 39828 237346 39840
rect 246022 39828 246028 39840
rect 237340 39800 246028 39828
rect 237340 39788 237346 39800
rect 246022 39788 246028 39800
rect 246080 39788 246086 39840
rect 248322 39788 248328 39840
rect 248380 39828 248386 39840
rect 255130 39828 255136 39840
rect 248380 39800 255136 39828
rect 248380 39788 248386 39800
rect 255130 39788 255136 39800
rect 255188 39788 255194 39840
rect 501690 39788 501696 39840
rect 501748 39828 501754 39840
rect 532694 39828 532700 39840
rect 501748 39800 532700 39828
rect 501748 39788 501754 39800
rect 532694 39788 532700 39800
rect 532752 39788 532758 39840
rect 535270 39788 535276 39840
rect 535328 39828 535334 39840
rect 562318 39828 562324 39840
rect 535328 39800 562324 39828
rect 535328 39788 535334 39800
rect 562318 39788 562324 39800
rect 562376 39788 562382 39840
rect 9582 39720 9588 39772
rect 9640 39760 9646 39772
rect 49510 39760 49516 39772
rect 9640 39732 49516 39760
rect 9640 39720 9646 39732
rect 49510 39720 49516 39732
rect 49568 39720 49574 39772
rect 63402 39720 63408 39772
rect 63460 39760 63466 39772
rect 96338 39760 96344 39772
rect 63460 39732 96344 39760
rect 63460 39720 63466 39732
rect 96338 39720 96344 39732
rect 96396 39720 96402 39772
rect 106182 39720 106188 39772
rect 106240 39760 106246 39772
rect 132954 39760 132960 39772
rect 106240 39732 132960 39760
rect 106240 39720 106246 39732
rect 132954 39720 132960 39732
rect 133012 39720 133018 39772
rect 139302 39720 139308 39772
rect 139360 39760 139366 39772
rect 161474 39760 161480 39772
rect 139360 39732 161480 39760
rect 139360 39720 139366 39732
rect 161474 39720 161480 39732
rect 161532 39720 161538 39772
rect 162762 39720 162768 39772
rect 162820 39760 162826 39772
rect 181898 39760 181904 39772
rect 162820 39732 181904 39760
rect 162820 39720 162826 39732
rect 181898 39720 181904 39732
rect 181956 39720 181962 39772
rect 184842 39720 184848 39772
rect 184900 39760 184906 39772
rect 200206 39760 200212 39772
rect 184900 39732 200212 39760
rect 184900 39720 184906 39732
rect 200206 39720 200212 39732
rect 200264 39720 200270 39772
rect 201402 39720 201408 39772
rect 201460 39760 201466 39772
rect 214466 39760 214472 39772
rect 201460 39732 214472 39760
rect 201460 39720 201466 39732
rect 214466 39720 214472 39732
rect 214524 39720 214530 39772
rect 219250 39720 219256 39772
rect 219308 39760 219314 39772
rect 229738 39760 229744 39772
rect 219308 39732 229744 39760
rect 219308 39720 219314 39732
rect 229738 39720 229744 39732
rect 229796 39720 229802 39772
rect 230382 39720 230388 39772
rect 230440 39760 230446 39772
rect 239858 39760 239864 39772
rect 230440 39732 239864 39760
rect 230440 39720 230446 39732
rect 239858 39720 239864 39732
rect 239916 39720 239922 39772
rect 241422 39720 241428 39772
rect 241480 39760 241486 39772
rect 249058 39760 249064 39772
rect 241480 39732 249064 39760
rect 241480 39720 241486 39732
rect 249058 39720 249064 39732
rect 249116 39720 249122 39772
rect 257982 39720 257988 39772
rect 258040 39760 258046 39772
rect 263318 39760 263324 39772
rect 258040 39732 263324 39760
rect 258040 39720 258046 39732
rect 263318 39720 263324 39732
rect 263376 39720 263382 39772
rect 498562 39720 498568 39772
rect 498620 39760 498626 39772
rect 518158 39760 518164 39772
rect 498620 39732 518164 39760
rect 498620 39720 498626 39732
rect 518158 39720 518164 39732
rect 518216 39720 518222 39772
rect 526070 39720 526076 39772
rect 526128 39760 526134 39772
rect 558178 39760 558184 39772
rect 526128 39732 558184 39760
rect 526128 39720 526134 39732
rect 558178 39720 558184 39732
rect 558236 39720 558242 39772
rect 10962 39652 10968 39704
rect 11020 39692 11026 39704
rect 50522 39692 50528 39704
rect 11020 39664 50528 39692
rect 11020 39652 11026 39664
rect 50522 39652 50528 39664
rect 50580 39652 50586 39704
rect 67542 39652 67548 39704
rect 67600 39692 67606 39704
rect 99374 39692 99380 39704
rect 67600 39664 99380 39692
rect 67600 39652 67606 39664
rect 99374 39652 99380 39664
rect 99432 39652 99438 39704
rect 100662 39652 100668 39704
rect 100720 39692 100726 39704
rect 127894 39692 127900 39704
rect 100720 39664 127900 39692
rect 100720 39652 100726 39664
rect 127894 39652 127900 39664
rect 127952 39652 127958 39704
rect 135162 39652 135168 39704
rect 135220 39692 135226 39704
rect 157426 39692 157432 39704
rect 135220 39664 157432 39692
rect 135220 39652 135226 39664
rect 157426 39652 157432 39664
rect 157484 39652 157490 39704
rect 160002 39652 160008 39704
rect 160060 39692 160066 39704
rect 178770 39692 178776 39704
rect 160060 39664 178776 39692
rect 160060 39652 160066 39664
rect 178770 39652 178776 39664
rect 178828 39652 178834 39704
rect 180702 39652 180708 39704
rect 180760 39692 180766 39704
rect 197170 39692 197176 39704
rect 180760 39664 197176 39692
rect 180760 39652 180766 39664
rect 197170 39652 197176 39664
rect 197228 39652 197234 39704
rect 198642 39652 198648 39704
rect 198700 39692 198706 39704
rect 212534 39692 212540 39704
rect 198700 39664 212540 39692
rect 198700 39652 198706 39664
rect 212534 39652 212540 39664
rect 212592 39652 212598 39704
rect 219342 39652 219348 39704
rect 219400 39692 219406 39704
rect 230750 39692 230756 39704
rect 219400 39664 230756 39692
rect 219400 39652 219406 39664
rect 230750 39652 230756 39664
rect 230808 39652 230814 39704
rect 233142 39652 233148 39704
rect 233200 39692 233206 39704
rect 241974 39692 241980 39704
rect 233200 39664 241980 39692
rect 233200 39652 233206 39664
rect 241974 39652 241980 39664
rect 242032 39652 242038 39704
rect 244182 39652 244188 39704
rect 244240 39692 244246 39704
rect 252094 39692 252100 39704
rect 244240 39664 252100 39692
rect 244240 39652 244246 39664
rect 252094 39652 252100 39664
rect 252152 39652 252158 39704
rect 267642 39652 267648 39704
rect 267700 39692 267706 39704
rect 271506 39692 271512 39704
rect 267700 39664 271512 39692
rect 267700 39652 267706 39664
rect 271506 39652 271512 39664
rect 271564 39652 271570 39704
rect 488442 39652 488448 39704
rect 488500 39692 488506 39704
rect 497458 39692 497464 39704
rect 488500 39664 497464 39692
rect 488500 39652 488506 39664
rect 497458 39652 497464 39664
rect 497516 39652 497522 39704
rect 512822 39652 512828 39704
rect 512880 39692 512886 39704
rect 512880 39664 541296 39692
rect 512880 39652 512886 39664
rect 16482 39584 16488 39636
rect 16540 39624 16546 39636
rect 55582 39624 55588 39636
rect 16540 39596 55588 39624
rect 16540 39584 16546 39596
rect 55582 39584 55588 39596
rect 55640 39584 55646 39636
rect 64138 39584 64144 39636
rect 64196 39624 64202 39636
rect 69842 39624 69848 39636
rect 64196 39596 69848 39624
rect 64196 39584 64202 39596
rect 69842 39584 69848 39596
rect 69900 39584 69906 39636
rect 70302 39584 70308 39636
rect 70360 39624 70366 39636
rect 102410 39624 102416 39636
rect 70360 39596 102416 39624
rect 70360 39584 70366 39596
rect 102410 39584 102416 39596
rect 102468 39584 102474 39636
rect 103330 39584 103336 39636
rect 103388 39624 103394 39636
rect 130930 39624 130936 39636
rect 103388 39596 130936 39624
rect 103388 39584 103394 39596
rect 130930 39584 130936 39596
rect 130988 39584 130994 39636
rect 137922 39584 137928 39636
rect 137980 39624 137986 39636
rect 160462 39624 160468 39636
rect 137980 39596 160468 39624
rect 137980 39584 137986 39596
rect 160462 39584 160468 39596
rect 160520 39584 160526 39636
rect 164142 39584 164148 39636
rect 164200 39624 164206 39636
rect 182910 39624 182916 39636
rect 164200 39596 182916 39624
rect 164200 39584 164206 39596
rect 182910 39584 182916 39596
rect 182968 39584 182974 39636
rect 183462 39584 183468 39636
rect 183520 39624 183526 39636
rect 199194 39624 199200 39636
rect 183520 39596 199200 39624
rect 183520 39584 183526 39596
rect 199194 39584 199200 39596
rect 199252 39584 199258 39636
rect 202690 39584 202696 39636
rect 202748 39624 202754 39636
rect 216490 39624 216496 39636
rect 202748 39596 216496 39624
rect 202748 39584 202754 39596
rect 216490 39584 216496 39596
rect 216548 39584 216554 39636
rect 216582 39584 216588 39636
rect 216640 39624 216646 39636
rect 227714 39624 227720 39636
rect 216640 39596 227720 39624
rect 216640 39584 216646 39596
rect 227714 39584 227720 39596
rect 227772 39584 227778 39636
rect 231762 39584 231768 39636
rect 231820 39624 231826 39636
rect 240962 39624 240968 39636
rect 231820 39596 240968 39624
rect 231820 39584 231826 39596
rect 240962 39584 240968 39596
rect 241020 39584 241026 39636
rect 264882 39584 264888 39636
rect 264940 39624 264946 39636
rect 269390 39624 269396 39636
rect 264940 39596 269396 39624
rect 264940 39584 264946 39596
rect 269390 39584 269396 39596
rect 269448 39584 269454 39636
rect 464982 39584 464988 39636
rect 465040 39624 465046 39636
rect 490006 39624 490012 39636
rect 465040 39596 490012 39624
rect 465040 39584 465046 39596
rect 490006 39584 490012 39596
rect 490064 39584 490070 39636
rect 491478 39584 491484 39636
rect 491536 39624 491542 39636
rect 512638 39624 512644 39636
rect 491536 39596 512644 39624
rect 491536 39584 491542 39596
rect 512638 39584 512644 39596
rect 512696 39584 512702 39636
rect 515950 39584 515956 39636
rect 516008 39624 516014 39636
rect 541161 39627 541219 39633
rect 541161 39624 541173 39627
rect 516008 39596 541173 39624
rect 516008 39584 516014 39596
rect 541161 39593 541173 39596
rect 541207 39593 541219 39627
rect 541268 39624 541296 39664
rect 541342 39652 541348 39704
rect 541400 39692 541406 39704
rect 548518 39692 548524 39704
rect 541400 39664 548524 39692
rect 541400 39652 541406 39664
rect 548518 39652 548524 39664
rect 548576 39652 548582 39704
rect 544378 39624 544384 39636
rect 541268 39596 544384 39624
rect 541161 39587 541219 39593
rect 544378 39584 544384 39596
rect 544436 39584 544442 39636
rect 13722 39516 13728 39568
rect 13780 39556 13786 39568
rect 53558 39556 53564 39568
rect 13780 39528 53564 39556
rect 13780 39516 13786 39528
rect 53558 39516 53564 39528
rect 53616 39516 53622 39568
rect 53742 39516 53748 39568
rect 53800 39556 53806 39568
rect 87138 39556 87144 39568
rect 53800 39528 87144 39556
rect 53800 39516 53806 39528
rect 87138 39516 87144 39528
rect 87196 39516 87202 39568
rect 88242 39516 88248 39568
rect 88300 39556 88306 39568
rect 117682 39556 117688 39568
rect 88300 39528 117688 39556
rect 88300 39516 88306 39528
rect 117682 39516 117688 39528
rect 117740 39516 117746 39568
rect 119982 39516 119988 39568
rect 120040 39556 120046 39568
rect 145190 39556 145196 39568
rect 120040 39528 145196 39556
rect 120040 39516 120046 39528
rect 145190 39516 145196 39528
rect 145248 39516 145254 39568
rect 146938 39516 146944 39568
rect 146996 39556 147002 39568
rect 154390 39556 154396 39568
rect 146996 39528 154396 39556
rect 146996 39516 147002 39528
rect 154390 39516 154396 39528
rect 154448 39516 154454 39568
rect 155129 39559 155187 39565
rect 155129 39525 155141 39559
rect 155175 39556 155187 39559
rect 167638 39556 167644 39568
rect 155175 39528 167644 39556
rect 155175 39525 155187 39528
rect 155129 39519 155187 39525
rect 167638 39516 167644 39528
rect 167696 39516 167702 39568
rect 169662 39516 169668 39568
rect 169720 39556 169726 39568
rect 187970 39556 187976 39568
rect 169720 39528 187976 39556
rect 169720 39516 169726 39528
rect 187970 39516 187976 39528
rect 188028 39516 188034 39568
rect 188982 39516 188988 39568
rect 189040 39556 189046 39568
rect 204254 39556 204260 39568
rect 189040 39528 204260 39556
rect 189040 39516 189046 39528
rect 204254 39516 204260 39528
rect 204312 39516 204318 39568
rect 206922 39516 206928 39568
rect 206980 39556 206986 39568
rect 219526 39556 219532 39568
rect 206980 39528 219532 39556
rect 206980 39516 206986 39528
rect 219526 39516 219532 39528
rect 219584 39516 219590 39568
rect 220722 39516 220728 39568
rect 220780 39556 220786 39568
rect 231854 39556 231860 39568
rect 220780 39528 231860 39556
rect 220780 39516 220786 39528
rect 231854 39516 231860 39528
rect 231912 39516 231918 39568
rect 234522 39516 234528 39568
rect 234580 39556 234586 39568
rect 242986 39556 242992 39568
rect 234580 39528 242992 39556
rect 234580 39516 234586 39528
rect 242986 39516 242992 39528
rect 243044 39516 243050 39568
rect 245562 39516 245568 39568
rect 245620 39556 245626 39568
rect 253106 39556 253112 39568
rect 245620 39528 253112 39556
rect 245620 39516 245626 39528
rect 253106 39516 253112 39528
rect 253164 39516 253170 39568
rect 256602 39516 256608 39568
rect 256660 39556 256666 39568
rect 262306 39556 262312 39568
rect 256660 39528 262312 39556
rect 256660 39516 256666 39528
rect 262306 39516 262312 39528
rect 262364 39516 262370 39568
rect 477218 39516 477224 39568
rect 477276 39556 477282 39568
rect 502978 39556 502984 39568
rect 477276 39528 502984 39556
rect 477276 39516 477282 39528
rect 502978 39516 502984 39528
rect 503036 39516 503042 39568
rect 503714 39516 503720 39568
rect 503772 39556 503778 39568
rect 522298 39556 522304 39568
rect 503772 39528 522304 39556
rect 503772 39516 503778 39528
rect 522298 39516 522304 39528
rect 522356 39516 522362 39568
rect 523034 39516 523040 39568
rect 523092 39556 523098 39568
rect 556798 39556 556804 39568
rect 523092 39528 556804 39556
rect 523092 39516 523098 39528
rect 556798 39516 556804 39528
rect 556856 39516 556862 39568
rect 12342 39448 12348 39500
rect 12400 39488 12406 39500
rect 51534 39488 51540 39500
rect 12400 39460 51540 39488
rect 12400 39448 12406 39460
rect 51534 39448 51540 39460
rect 51592 39448 51598 39500
rect 56502 39448 56508 39500
rect 56560 39488 56566 39500
rect 90266 39488 90272 39500
rect 56560 39460 90272 39488
rect 56560 39448 56566 39460
rect 90266 39448 90272 39460
rect 90324 39448 90330 39500
rect 92382 39448 92388 39500
rect 92440 39488 92446 39500
rect 120810 39488 120816 39500
rect 92440 39460 120816 39488
rect 92440 39448 92446 39460
rect 120810 39448 120816 39460
rect 120868 39448 120874 39500
rect 121362 39448 121368 39500
rect 121420 39488 121426 39500
rect 146294 39488 146300 39500
rect 121420 39460 146300 39488
rect 121420 39448 121426 39460
rect 146294 39448 146300 39460
rect 146352 39448 146358 39500
rect 148962 39448 148968 39500
rect 149020 39488 149026 39500
rect 169754 39488 169760 39500
rect 149020 39460 169760 39488
rect 149020 39448 149026 39460
rect 169754 39448 169760 39460
rect 169812 39448 169818 39500
rect 171042 39448 171048 39500
rect 171100 39488 171106 39500
rect 189074 39488 189080 39500
rect 171100 39460 189080 39488
rect 171100 39448 171106 39460
rect 189074 39448 189080 39460
rect 189132 39448 189138 39500
rect 194410 39448 194416 39500
rect 194468 39488 194474 39500
rect 208394 39488 208400 39500
rect 194468 39460 208400 39488
rect 194468 39448 194474 39460
rect 208394 39448 208400 39460
rect 208452 39448 208458 39500
rect 215202 39448 215208 39500
rect 215260 39488 215266 39500
rect 226702 39488 226708 39500
rect 215260 39460 226708 39488
rect 215260 39448 215266 39460
rect 226702 39448 226708 39460
rect 226760 39448 226766 39500
rect 235810 39448 235816 39500
rect 235868 39488 235874 39500
rect 245010 39488 245016 39500
rect 235868 39460 245016 39488
rect 235868 39448 235874 39460
rect 245010 39448 245016 39460
rect 245068 39448 245074 39500
rect 246942 39448 246948 39500
rect 247000 39488 247006 39500
rect 254118 39488 254124 39500
rect 247000 39460 254124 39488
rect 247000 39448 247006 39460
rect 254118 39448 254124 39460
rect 254176 39448 254182 39500
rect 255222 39448 255228 39500
rect 255280 39488 255286 39500
rect 261294 39488 261300 39500
rect 255280 39460 261300 39488
rect 255280 39448 255286 39460
rect 261294 39448 261300 39460
rect 261352 39448 261358 39500
rect 266998 39448 267004 39500
rect 267056 39488 267062 39500
rect 270494 39488 270500 39500
rect 267056 39460 270500 39488
rect 267056 39448 267062 39460
rect 270494 39448 270500 39460
rect 270552 39448 270558 39500
rect 332686 39448 332692 39500
rect 332744 39488 332750 39500
rect 335998 39488 336004 39500
rect 332744 39460 336004 39488
rect 332744 39448 332750 39460
rect 335998 39448 336004 39460
rect 336056 39448 336062 39500
rect 480254 39448 480260 39500
rect 480312 39488 480318 39500
rect 507854 39488 507860 39500
rect 480312 39460 507860 39488
rect 480312 39448 480318 39460
rect 507854 39448 507860 39460
rect 507912 39448 507918 39500
rect 516962 39448 516968 39500
rect 517020 39488 517026 39500
rect 550634 39488 550640 39500
rect 517020 39460 550640 39488
rect 517020 39448 517026 39460
rect 550634 39448 550640 39460
rect 550692 39448 550698 39500
rect 6822 39380 6828 39432
rect 6880 39420 6886 39432
rect 47486 39420 47492 39432
rect 6880 39392 47492 39420
rect 6880 39380 6886 39392
rect 47486 39380 47492 39392
rect 47544 39380 47550 39432
rect 57882 39380 57888 39432
rect 57940 39420 57946 39432
rect 91278 39420 91284 39432
rect 57940 39392 91284 39420
rect 57940 39380 57946 39392
rect 91278 39380 91284 39392
rect 91336 39380 91342 39432
rect 99282 39380 99288 39432
rect 99340 39420 99346 39432
rect 126974 39420 126980 39432
rect 99340 39392 126980 39420
rect 99340 39380 99346 39392
rect 126974 39380 126980 39392
rect 127032 39380 127038 39432
rect 132402 39380 132408 39432
rect 132460 39420 132466 39432
rect 155402 39420 155408 39432
rect 132460 39392 155408 39420
rect 132460 39380 132466 39392
rect 155402 39380 155408 39392
rect 155460 39380 155466 39432
rect 155862 39380 155868 39432
rect 155920 39420 155926 39432
rect 175734 39420 175740 39432
rect 155920 39392 175740 39420
rect 155920 39380 155926 39392
rect 175734 39380 175740 39392
rect 175792 39380 175798 39432
rect 179322 39380 179328 39432
rect 179380 39420 179386 39432
rect 196158 39420 196164 39432
rect 179380 39392 196164 39420
rect 179380 39380 179386 39392
rect 196158 39380 196164 39392
rect 196216 39380 196222 39432
rect 197262 39380 197268 39432
rect 197320 39420 197326 39432
rect 211430 39420 211436 39432
rect 197320 39392 211436 39420
rect 197320 39380 197326 39392
rect 211430 39380 211436 39392
rect 211488 39380 211494 39432
rect 213822 39380 213828 39432
rect 213880 39420 213886 39432
rect 225690 39420 225696 39432
rect 213880 39392 225696 39420
rect 213880 39380 213886 39392
rect 225690 39380 225696 39392
rect 225748 39380 225754 39432
rect 229002 39380 229008 39432
rect 229060 39420 229066 39432
rect 238846 39420 238852 39432
rect 229060 39392 238852 39420
rect 229060 39380 229066 39392
rect 238846 39380 238852 39392
rect 238904 39380 238910 39432
rect 244090 39380 244096 39432
rect 244148 39420 244154 39432
rect 251174 39420 251180 39432
rect 244148 39392 251180 39420
rect 244148 39380 244154 39392
rect 251174 39380 251180 39392
rect 251232 39380 251238 39432
rect 434438 39380 434444 39432
rect 434496 39420 434502 39432
rect 443546 39420 443552 39432
rect 434496 39392 443552 39420
rect 434496 39380 434502 39392
rect 443546 39380 443552 39392
rect 443604 39380 443610 39432
rect 458910 39380 458916 39432
rect 458968 39420 458974 39432
rect 483014 39420 483020 39432
rect 458968 39392 483020 39420
rect 458968 39380 458974 39392
rect 483014 39380 483020 39392
rect 483072 39380 483078 39432
rect 483290 39380 483296 39432
rect 483348 39420 483354 39432
rect 511994 39420 512000 39432
rect 483348 39392 512000 39420
rect 483348 39380 483354 39392
rect 511994 39380 512000 39392
rect 512052 39380 512058 39432
rect 519998 39380 520004 39432
rect 520056 39420 520062 39432
rect 554774 39420 554780 39432
rect 520056 39392 554780 39420
rect 520056 39380 520062 39392
rect 554774 39380 554780 39392
rect 554832 39380 554838 39432
rect 4062 39312 4068 39364
rect 4120 39352 4126 39364
rect 45554 39352 45560 39364
rect 4120 39324 45560 39352
rect 4120 39312 4126 39324
rect 45554 39312 45560 39324
rect 45612 39312 45618 39364
rect 49602 39312 49608 39364
rect 49660 39352 49666 39364
rect 84194 39352 84200 39364
rect 49660 39324 84200 39352
rect 49660 39312 49666 39324
rect 84194 39312 84200 39324
rect 84252 39312 84258 39364
rect 85482 39312 85488 39364
rect 85540 39352 85546 39364
rect 114646 39352 114652 39364
rect 85540 39324 114652 39352
rect 85540 39312 85546 39324
rect 114646 39312 114652 39324
rect 114704 39312 114710 39364
rect 117222 39312 117228 39364
rect 117280 39352 117286 39364
rect 142154 39352 142160 39364
rect 117280 39324 142160 39352
rect 117280 39312 117286 39324
rect 142154 39312 142160 39324
rect 142212 39312 142218 39364
rect 144730 39312 144736 39364
rect 144788 39352 144794 39364
rect 165614 39352 165620 39364
rect 144788 39324 165620 39352
rect 144788 39312 144794 39324
rect 165614 39312 165620 39324
rect 165672 39312 165678 39364
rect 166902 39312 166908 39364
rect 166960 39352 166966 39364
rect 184934 39352 184940 39364
rect 166960 39324 184940 39352
rect 166960 39312 166966 39324
rect 184934 39312 184940 39324
rect 184992 39312 184998 39364
rect 186130 39312 186136 39364
rect 186188 39352 186194 39364
rect 202230 39352 202236 39364
rect 186188 39324 202236 39352
rect 186188 39312 186194 39324
rect 202230 39312 202236 39324
rect 202288 39312 202294 39364
rect 210970 39312 210976 39364
rect 211028 39352 211034 39364
rect 223574 39352 223580 39364
rect 211028 39324 223580 39352
rect 211028 39312 211034 39324
rect 223574 39312 223580 39324
rect 223632 39312 223638 39364
rect 227530 39312 227536 39364
rect 227588 39352 227594 39364
rect 237834 39352 237840 39364
rect 227588 39324 237840 39352
rect 227588 39312 227594 39324
rect 237834 39312 237840 39324
rect 237892 39312 237898 39364
rect 238662 39312 238668 39364
rect 238720 39352 238726 39364
rect 247034 39352 247040 39364
rect 238720 39324 247040 39352
rect 238720 39312 238726 39324
rect 247034 39312 247040 39324
rect 247092 39312 247098 39364
rect 277210 39312 277216 39364
rect 277268 39352 277274 39364
rect 280614 39352 280620 39364
rect 277268 39324 280620 39352
rect 277268 39312 277274 39324
rect 280614 39312 280620 39324
rect 280672 39312 280678 39364
rect 343818 39312 343824 39364
rect 343876 39352 343882 39364
rect 349246 39352 349252 39364
rect 343876 39324 349252 39352
rect 343876 39312 343882 39324
rect 349246 39312 349252 39324
rect 349304 39312 349310 39364
rect 437474 39312 437480 39364
rect 437532 39352 437538 39364
rect 454678 39352 454684 39364
rect 437532 39324 454684 39352
rect 437532 39312 437538 39324
rect 454678 39312 454684 39324
rect 454736 39312 454742 39364
rect 455874 39312 455880 39364
rect 455932 39352 455938 39364
rect 465718 39352 465724 39364
rect 455932 39324 465724 39352
rect 455932 39312 455938 39324
rect 465718 39312 465724 39324
rect 465776 39312 465782 39364
rect 474182 39312 474188 39364
rect 474240 39352 474246 39364
rect 474240 39324 489914 39352
rect 474240 39312 474246 39324
rect 31662 39244 31668 39296
rect 31720 39284 31726 39296
rect 68830 39284 68836 39296
rect 31720 39256 68836 39284
rect 31720 39244 31726 39256
rect 68830 39244 68836 39256
rect 68888 39244 68894 39296
rect 71774 39244 71780 39296
rect 71832 39284 71838 39296
rect 73982 39284 73988 39296
rect 71832 39256 73988 39284
rect 71832 39244 71838 39256
rect 73982 39244 73988 39256
rect 74040 39244 74046 39296
rect 75178 39244 75184 39296
rect 75236 39284 75242 39296
rect 82078 39284 82084 39296
rect 75236 39256 82084 39284
rect 75236 39244 75242 39256
rect 82078 39244 82084 39256
rect 82136 39244 82142 39296
rect 111610 39284 111616 39296
rect 82464 39256 111616 39284
rect 28902 39176 28908 39228
rect 28960 39216 28966 39228
rect 65794 39216 65800 39228
rect 28960 39188 65800 39216
rect 28960 39176 28966 39188
rect 65794 39176 65800 39188
rect 65852 39176 65858 39228
rect 68278 39176 68284 39228
rect 68336 39216 68342 39228
rect 68336 39188 78536 39216
rect 68336 39176 68342 39188
rect 35802 39108 35808 39160
rect 35860 39148 35866 39160
rect 71866 39148 71872 39160
rect 35860 39120 71872 39148
rect 35860 39108 35866 39120
rect 71866 39108 71872 39120
rect 71924 39108 71930 39160
rect 72418 39108 72424 39160
rect 72476 39148 72482 39160
rect 73062 39148 73068 39160
rect 72476 39120 73068 39148
rect 72476 39108 72482 39120
rect 73062 39108 73068 39120
rect 73120 39108 73126 39160
rect 39298 39040 39304 39092
rect 39356 39080 39362 39092
rect 74994 39080 75000 39092
rect 39356 39052 75000 39080
rect 39356 39040 39362 39052
rect 74994 39040 75000 39052
rect 75052 39040 75058 39092
rect 78508 39080 78536 39188
rect 81342 39176 81348 39228
rect 81400 39216 81406 39228
rect 82464 39216 82492 39256
rect 111610 39244 111616 39256
rect 111668 39244 111674 39296
rect 113082 39244 113088 39296
rect 113140 39284 113146 39296
rect 139118 39284 139124 39296
rect 113140 39256 139124 39284
rect 113140 39244 113146 39256
rect 139118 39244 139124 39256
rect 139176 39244 139182 39296
rect 143442 39244 143448 39296
rect 143500 39284 143506 39296
rect 164602 39284 164608 39296
rect 143500 39256 164608 39284
rect 143500 39244 143506 39256
rect 164602 39244 164608 39256
rect 164660 39244 164666 39296
rect 172422 39244 172428 39296
rect 172480 39284 172486 39296
rect 189994 39284 190000 39296
rect 172480 39256 190000 39284
rect 172480 39244 172486 39256
rect 189994 39244 190000 39256
rect 190052 39244 190058 39296
rect 193122 39244 193128 39296
rect 193180 39284 193186 39296
rect 207290 39284 207296 39296
rect 193180 39256 207296 39284
rect 193180 39244 193186 39256
rect 207290 39244 207296 39256
rect 207348 39244 207354 39296
rect 208302 39244 208308 39296
rect 208360 39284 208366 39296
rect 220538 39284 220544 39296
rect 208360 39256 220544 39284
rect 208360 39244 208366 39256
rect 220538 39244 220544 39256
rect 220596 39244 220602 39296
rect 227622 39244 227628 39296
rect 227680 39284 227686 39296
rect 236822 39284 236828 39296
rect 227680 39256 236828 39284
rect 227680 39244 227686 39256
rect 236822 39244 236828 39256
rect 236880 39244 236886 39296
rect 489886 39284 489914 39324
rect 510798 39312 510804 39364
rect 510856 39352 510862 39364
rect 542998 39352 543004 39364
rect 510856 39324 543004 39352
rect 510856 39312 510862 39324
rect 542998 39312 543004 39324
rect 543056 39312 543062 39364
rect 543642 39312 543648 39364
rect 543700 39352 543706 39364
rect 582377 39355 582435 39361
rect 582377 39352 582389 39355
rect 543700 39324 582389 39352
rect 543700 39312 543706 39324
rect 582377 39321 582389 39324
rect 582423 39321 582435 39355
rect 582377 39315 582435 39321
rect 500954 39284 500960 39296
rect 489886 39256 500960 39284
rect 500954 39244 500960 39256
rect 501012 39244 501018 39296
rect 528094 39244 528100 39296
rect 528152 39284 528158 39296
rect 540238 39284 540244 39296
rect 528152 39256 540244 39284
rect 528152 39244 528158 39256
rect 540238 39244 540244 39256
rect 540296 39244 540302 39296
rect 541161 39287 541219 39293
rect 541161 39253 541173 39287
rect 541207 39284 541219 39287
rect 547230 39284 547236 39296
rect 541207 39256 547236 39284
rect 541207 39253 541219 39256
rect 541161 39247 541219 39253
rect 547230 39244 547236 39256
rect 547288 39244 547294 39296
rect 108574 39216 108580 39228
rect 81400 39188 82492 39216
rect 84166 39188 108580 39216
rect 81400 39176 81406 39188
rect 78582 39108 78588 39160
rect 78640 39148 78646 39160
rect 84166 39148 84194 39188
rect 108574 39176 108580 39188
rect 108632 39176 108638 39228
rect 114462 39176 114468 39228
rect 114520 39216 114526 39228
rect 140130 39216 140136 39228
rect 114520 39188 140136 39216
rect 114520 39176 114526 39188
rect 140130 39176 140136 39188
rect 140188 39176 140194 39228
rect 140682 39176 140688 39228
rect 140740 39216 140746 39228
rect 162486 39216 162492 39228
rect 140740 39188 162492 39216
rect 140740 39176 140746 39188
rect 162486 39176 162492 39188
rect 162544 39176 162550 39228
rect 168282 39176 168288 39228
rect 168340 39216 168346 39228
rect 185946 39216 185952 39228
rect 168340 39188 185952 39216
rect 168340 39176 168346 39188
rect 185946 39176 185952 39188
rect 186004 39176 186010 39228
rect 191742 39176 191748 39228
rect 191800 39216 191806 39228
rect 206278 39216 206284 39228
rect 191800 39188 206284 39216
rect 191800 39176 191806 39188
rect 206278 39176 206284 39188
rect 206336 39176 206342 39228
rect 209682 39176 209688 39228
rect 209740 39216 209746 39228
rect 221550 39216 221556 39228
rect 209740 39188 221556 39216
rect 209740 39176 209746 39188
rect 221550 39176 221556 39188
rect 221608 39176 221614 39228
rect 226242 39176 226248 39228
rect 226300 39216 226306 39228
rect 235718 39216 235724 39228
rect 226300 39188 235724 39216
rect 226300 39176 226306 39188
rect 235718 39176 235724 39188
rect 235776 39176 235782 39228
rect 274542 39176 274548 39228
rect 274600 39216 274606 39228
rect 277578 39216 277584 39228
rect 274600 39188 277584 39216
rect 274600 39176 274606 39188
rect 277578 39176 277584 39188
rect 277636 39176 277642 39228
rect 534258 39176 534264 39228
rect 534316 39216 534322 39228
rect 541618 39216 541624 39228
rect 534316 39188 541624 39216
rect 534316 39176 534322 39188
rect 541618 39176 541624 39188
rect 541676 39176 541682 39228
rect 78640 39120 84194 39148
rect 78640 39108 78646 39120
rect 84838 39108 84844 39160
rect 84896 39148 84902 39160
rect 112622 39148 112628 39160
rect 84896 39120 112628 39148
rect 84896 39108 84902 39120
rect 112622 39108 112628 39120
rect 112680 39108 112686 39160
rect 115842 39108 115848 39160
rect 115900 39148 115906 39160
rect 141142 39148 141148 39160
rect 115900 39120 141148 39148
rect 115900 39108 115906 39120
rect 141142 39108 141148 39120
rect 141200 39108 141206 39160
rect 147582 39108 147588 39160
rect 147640 39148 147646 39160
rect 168650 39148 168656 39160
rect 147640 39120 168656 39148
rect 147640 39108 147646 39120
rect 168650 39108 168656 39120
rect 168708 39108 168714 39160
rect 175182 39108 175188 39160
rect 175240 39148 175246 39160
rect 192018 39148 192024 39160
rect 175240 39120 192024 39148
rect 175240 39108 175246 39120
rect 192018 39108 192024 39120
rect 192076 39108 192082 39160
rect 194502 39108 194508 39160
rect 194560 39148 194566 39160
rect 209314 39148 209320 39160
rect 194560 39120 209320 39148
rect 194560 39108 194566 39120
rect 209314 39108 209320 39120
rect 209372 39108 209378 39160
rect 212442 39108 212448 39160
rect 212500 39148 212506 39160
rect 224586 39148 224592 39160
rect 212500 39120 224592 39148
rect 212500 39108 212506 39120
rect 224586 39108 224592 39120
rect 224644 39108 224650 39160
rect 78508 39052 79180 39080
rect 44082 38972 44088 39024
rect 44140 39012 44146 39024
rect 79042 39012 79048 39024
rect 44140 38984 79048 39012
rect 44140 38972 44146 38984
rect 79042 38972 79048 38984
rect 79100 38972 79106 39024
rect 79152 39012 79180 39052
rect 82078 39040 82084 39092
rect 82136 39080 82142 39092
rect 109586 39080 109592 39092
rect 82136 39052 109592 39080
rect 82136 39040 82142 39052
rect 109586 39040 109592 39052
rect 109644 39040 109650 39092
rect 111702 39040 111708 39092
rect 111760 39080 111766 39092
rect 137094 39080 137100 39092
rect 111760 39052 137100 39080
rect 111760 39040 111766 39052
rect 137094 39040 137100 39052
rect 137152 39040 137158 39092
rect 137278 39040 137284 39092
rect 137336 39080 137342 39092
rect 138106 39080 138112 39092
rect 137336 39052 138112 39080
rect 137336 39040 137342 39052
rect 138106 39040 138112 39052
rect 138164 39040 138170 39092
rect 153102 39040 153108 39092
rect 153160 39080 153166 39092
rect 172698 39080 172704 39092
rect 153160 39052 172704 39080
rect 153160 39040 153166 39052
rect 172698 39040 172704 39052
rect 172756 39040 172762 39092
rect 177850 39040 177856 39092
rect 177908 39080 177914 39092
rect 194042 39080 194048 39092
rect 177908 39052 194048 39080
rect 177908 39040 177914 39052
rect 194042 39040 194048 39052
rect 194100 39040 194106 39092
rect 202782 39040 202788 39092
rect 202840 39080 202846 39092
rect 215478 39080 215484 39092
rect 202840 39052 215484 39080
rect 202840 39040 202846 39052
rect 215478 39040 215484 39052
rect 215536 39040 215542 39092
rect 252370 39040 252376 39092
rect 252428 39080 252434 39092
rect 259270 39080 259276 39092
rect 252428 39052 259276 39080
rect 252428 39040 252434 39052
rect 259270 39040 259276 39052
rect 259328 39040 259334 39092
rect 259362 39040 259368 39092
rect 259420 39080 259426 39092
rect 264330 39080 264336 39092
rect 259420 39052 264336 39080
rect 259420 39040 259426 39052
rect 264330 39040 264336 39052
rect 264388 39040 264394 39092
rect 269022 39040 269028 39092
rect 269080 39080 269086 39092
rect 273530 39080 273536 39092
rect 269080 39052 273536 39080
rect 269080 39040 269086 39052
rect 273530 39040 273536 39052
rect 273588 39040 273594 39092
rect 85114 39012 85120 39024
rect 79152 38984 85120 39012
rect 85114 38972 85120 38984
rect 85172 38972 85178 39024
rect 91738 38972 91744 39024
rect 91796 39012 91802 39024
rect 118786 39012 118792 39024
rect 91796 38984 118792 39012
rect 91796 38972 91802 38984
rect 118786 38972 118792 38984
rect 118844 38972 118850 39024
rect 119890 38972 119896 39024
rect 119948 39012 119954 39024
rect 144178 39012 144184 39024
rect 119948 38984 144184 39012
rect 119948 38972 119954 38984
rect 144178 38972 144184 38984
rect 144236 38972 144242 39024
rect 150342 38972 150348 39024
rect 150400 39012 150406 39024
rect 170674 39012 170680 39024
rect 150400 38984 170680 39012
rect 150400 38972 150406 38984
rect 170674 38972 170680 38984
rect 170732 38972 170738 39024
rect 176562 38972 176568 39024
rect 176620 39012 176626 39024
rect 193030 39012 193036 39024
rect 176620 38984 193036 39012
rect 176620 38972 176626 38984
rect 193030 38972 193036 38984
rect 193088 38972 193094 39024
rect 240042 38972 240048 39024
rect 240100 39012 240106 39024
rect 248046 39012 248052 39024
rect 240100 38984 248052 39012
rect 240100 38972 240106 38984
rect 248046 38972 248052 38984
rect 248104 38972 248110 39024
rect 251082 38972 251088 39024
rect 251140 39012 251146 39024
rect 257246 39012 257252 39024
rect 251140 38984 257252 39012
rect 251140 38972 251146 38984
rect 257246 38972 257252 38984
rect 257304 38972 257310 39024
rect 260742 38972 260748 39024
rect 260800 39012 260806 39024
rect 265342 39012 265348 39024
rect 260800 38984 265348 39012
rect 260800 38972 260806 38984
rect 265342 38972 265348 38984
rect 265400 38972 265406 39024
rect 271782 38972 271788 39024
rect 271840 39012 271846 39024
rect 275554 39012 275560 39024
rect 271840 38984 275560 39012
rect 271840 38972 271846 38984
rect 275554 38972 275560 38984
rect 275612 38972 275618 39024
rect 282822 38972 282828 39024
rect 282880 39012 282886 39024
rect 284662 39012 284668 39024
rect 282880 38984 284668 39012
rect 282880 38972 282886 38984
rect 284662 38972 284668 38984
rect 284720 38972 284726 39024
rect 284938 38972 284944 39024
rect 284996 39012 285002 39024
rect 285674 39012 285680 39024
rect 284996 38984 285680 39012
rect 284996 38972 285002 38984
rect 285674 38972 285680 38984
rect 285732 38972 285738 39024
rect 289722 38972 289728 39024
rect 289780 39012 289786 39024
rect 290826 39012 290832 39024
rect 289780 38984 290832 39012
rect 289780 38972 289786 38984
rect 290826 38972 290832 38984
rect 290884 38972 290890 39024
rect 296714 38972 296720 39024
rect 296772 39012 296778 39024
rect 297910 39012 297916 39024
rect 296772 38984 297916 39012
rect 296772 38972 296778 38984
rect 297910 38972 297916 38984
rect 297968 38972 297974 39024
rect 303614 38972 303620 39024
rect 303672 39012 303678 39024
rect 304074 39012 304080 39024
rect 303672 38984 304080 39012
rect 303672 38972 303678 38984
rect 304074 38972 304080 38984
rect 304132 38972 304138 39024
rect 307202 38972 307208 39024
rect 307260 39012 307266 39024
rect 307662 39012 307668 39024
rect 307260 38984 307668 39012
rect 307260 38972 307266 38984
rect 307662 38972 307668 38984
rect 307720 38972 307726 39024
rect 311250 38972 311256 39024
rect 311308 39012 311314 39024
rect 311802 39012 311808 39024
rect 311308 38984 311808 39012
rect 311308 38972 311314 38984
rect 311802 38972 311808 38984
rect 311860 38972 311866 39024
rect 313274 38972 313280 39024
rect 313332 39012 313338 39024
rect 314562 39012 314568 39024
rect 313332 38984 314568 39012
rect 313332 38972 313338 38984
rect 314562 38972 314568 38984
rect 314620 38972 314626 39024
rect 316402 38972 316408 39024
rect 316460 39012 316466 39024
rect 317322 39012 317328 39024
rect 316460 38984 317328 39012
rect 316460 38972 316466 38984
rect 317322 38972 317328 38984
rect 317380 38972 317386 39024
rect 317414 38972 317420 39024
rect 317472 39012 317478 39024
rect 318702 39012 318708 39024
rect 317472 38984 318708 39012
rect 317472 38972 317478 38984
rect 318702 38972 318708 38984
rect 318760 38972 318766 39024
rect 320450 38972 320456 39024
rect 320508 39012 320514 39024
rect 321462 39012 321468 39024
rect 320508 38984 321468 39012
rect 320508 38972 320514 38984
rect 321462 38972 321468 38984
rect 321520 38972 321526 39024
rect 323486 38972 323492 39024
rect 323544 39012 323550 39024
rect 324222 39012 324228 39024
rect 323544 38984 324228 39012
rect 323544 38972 323550 38984
rect 324222 38972 324228 38984
rect 324280 38972 324286 39024
rect 324498 38972 324504 39024
rect 324556 39012 324562 39024
rect 325510 39012 325516 39024
rect 324556 38984 325516 39012
rect 324556 38972 324562 38984
rect 325510 38972 325516 38984
rect 325568 38972 325574 39024
rect 326522 38972 326528 39024
rect 326580 39012 326586 39024
rect 326982 39012 326988 39024
rect 326580 38984 326988 39012
rect 326580 38972 326586 38984
rect 326982 38972 326988 38984
rect 327040 38972 327046 39024
rect 327534 38972 327540 39024
rect 327592 39012 327598 39024
rect 328362 39012 328368 39024
rect 327592 38984 328368 39012
rect 327592 38972 327598 38984
rect 328362 38972 328368 38984
rect 328420 38972 328426 39024
rect 328546 38972 328552 39024
rect 328604 39012 328610 39024
rect 329742 39012 329748 39024
rect 328604 38984 329748 39012
rect 328604 38972 328610 38984
rect 329742 38972 329748 38984
rect 329800 38972 329806 39024
rect 330570 38972 330576 39024
rect 330628 39012 330634 39024
rect 331122 39012 331128 39024
rect 330628 38984 331128 39012
rect 330628 38972 330634 38984
rect 331122 38972 331128 38984
rect 331180 38972 331186 39024
rect 331674 38972 331680 39024
rect 331732 39012 331738 39024
rect 332502 39012 332508 39024
rect 331732 38984 332508 39012
rect 331732 38972 331738 38984
rect 332502 38972 332508 38984
rect 332560 38972 332566 39024
rect 333698 38972 333704 39024
rect 333756 39012 333762 39024
rect 334618 39012 334624 39024
rect 333756 38984 334624 39012
rect 333756 38972 333762 38984
rect 334618 38972 334624 38984
rect 334676 38972 334682 39024
rect 334710 38972 334716 39024
rect 334768 39012 334774 39024
rect 335262 39012 335268 39024
rect 334768 38984 335268 39012
rect 334768 38972 334774 38984
rect 335262 38972 335268 38984
rect 335320 38972 335326 39024
rect 335722 38972 335728 39024
rect 335780 39012 335786 39024
rect 336642 39012 336648 39024
rect 335780 38984 336648 39012
rect 335780 38972 335786 38984
rect 336642 38972 336648 38984
rect 336700 38972 336706 39024
rect 338758 38972 338764 39024
rect 338816 39012 338822 39024
rect 339402 39012 339408 39024
rect 338816 38984 339408 39012
rect 338816 38972 338822 38984
rect 339402 38972 339408 38984
rect 339460 38972 339466 39024
rect 339770 38972 339776 39024
rect 339828 39012 339834 39024
rect 340782 39012 340788 39024
rect 339828 38984 340788 39012
rect 339828 38972 339834 38984
rect 340782 38972 340788 38984
rect 340840 38972 340846 39024
rect 342806 38972 342812 39024
rect 342864 39012 342870 39024
rect 343542 39012 343548 39024
rect 342864 38984 343548 39012
rect 342864 38972 342870 38984
rect 343542 38972 343548 38984
rect 343600 38972 343606 39024
rect 345842 38972 345848 39024
rect 345900 39012 345906 39024
rect 346302 39012 346308 39024
rect 345900 38984 346308 39012
rect 345900 38972 345906 38984
rect 346302 38972 346308 38984
rect 346360 38972 346366 39024
rect 346946 38972 346952 39024
rect 347004 39012 347010 39024
rect 347682 39012 347688 39024
rect 347004 38984 347688 39012
rect 347004 38972 347010 38984
rect 347682 38972 347688 38984
rect 347740 38972 347746 39024
rect 347958 38972 347964 39024
rect 348016 39012 348022 39024
rect 348970 39012 348976 39024
rect 348016 38984 348976 39012
rect 348016 38972 348022 38984
rect 348970 38972 348976 38984
rect 349028 38972 349034 39024
rect 349982 38972 349988 39024
rect 350040 39012 350046 39024
rect 350442 39012 350448 39024
rect 350040 38984 350448 39012
rect 350040 38972 350046 38984
rect 350442 38972 350448 38984
rect 350500 38972 350506 39024
rect 350994 38972 351000 39024
rect 351052 39012 351058 39024
rect 351822 39012 351828 39024
rect 351052 38984 351828 39012
rect 351052 38972 351058 38984
rect 351822 38972 351828 38984
rect 351880 38972 351886 39024
rect 352006 38972 352012 39024
rect 352064 39012 352070 39024
rect 353202 39012 353208 39024
rect 352064 38984 353208 39012
rect 352064 38972 352070 38984
rect 353202 38972 353208 38984
rect 353260 38972 353266 39024
rect 354030 38972 354036 39024
rect 354088 39012 354094 39024
rect 354582 39012 354588 39024
rect 354088 38984 354588 39012
rect 354088 38972 354094 38984
rect 354582 38972 354588 38984
rect 354640 38972 354646 39024
rect 355042 38972 355048 39024
rect 355100 39012 355106 39024
rect 355962 39012 355968 39024
rect 355100 38984 355968 39012
rect 355100 38972 355106 38984
rect 355962 38972 355968 38984
rect 356020 38972 356026 39024
rect 356054 38972 356060 39024
rect 356112 39012 356118 39024
rect 357342 39012 357348 39024
rect 356112 38984 357348 39012
rect 356112 38972 356118 38984
rect 357342 38972 357348 38984
rect 357400 38972 357406 39024
rect 358078 38972 358084 39024
rect 358136 39012 358142 39024
rect 358722 39012 358728 39024
rect 358136 38984 358728 39012
rect 358136 38972 358142 38984
rect 358722 38972 358728 38984
rect 358780 38972 358786 39024
rect 359090 38972 359096 39024
rect 359148 39012 359154 39024
rect 360102 39012 360108 39024
rect 359148 38984 360108 39012
rect 359148 38972 359154 38984
rect 360102 38972 360108 38984
rect 360160 38972 360166 39024
rect 363230 38972 363236 39024
rect 363288 39012 363294 39024
rect 364242 39012 364248 39024
rect 363288 38984 364248 39012
rect 363288 38972 363294 38984
rect 364242 38972 364248 38984
rect 364300 38972 364306 39024
rect 366266 38972 366272 39024
rect 366324 39012 366330 39024
rect 367002 39012 367008 39024
rect 366324 38984 367008 39012
rect 366324 38972 366330 38984
rect 367002 38972 367008 38984
rect 367060 38972 367066 39024
rect 367278 38972 367284 39024
rect 367336 39012 367342 39024
rect 368290 39012 368296 39024
rect 367336 38984 368296 39012
rect 367336 38972 367342 38984
rect 368290 38972 368296 38984
rect 368348 38972 368354 39024
rect 369302 38972 369308 39024
rect 369360 39012 369366 39024
rect 369762 39012 369768 39024
rect 369360 38984 369768 39012
rect 369360 38972 369366 38984
rect 369762 38972 369768 38984
rect 369820 38972 369826 39024
rect 370314 38972 370320 39024
rect 370372 39012 370378 39024
rect 371142 39012 371148 39024
rect 370372 38984 371148 39012
rect 370372 38972 370378 38984
rect 371142 38972 371148 38984
rect 371200 38972 371206 39024
rect 371326 38972 371332 39024
rect 371384 39012 371390 39024
rect 372522 39012 372528 39024
rect 371384 38984 372528 39012
rect 371384 38972 371390 38984
rect 372522 38972 372528 38984
rect 372580 38972 372586 39024
rect 373350 38972 373356 39024
rect 373408 39012 373414 39024
rect 373902 39012 373908 39024
rect 373408 38984 373908 39012
rect 373408 38972 373414 38984
rect 373902 38972 373908 38984
rect 373960 38972 373966 39024
rect 374362 38972 374368 39024
rect 374420 39012 374426 39024
rect 375282 39012 375288 39024
rect 374420 38984 375288 39012
rect 374420 38972 374426 38984
rect 375282 38972 375288 38984
rect 375340 38972 375346 39024
rect 377490 38972 377496 39024
rect 377548 39012 377554 39024
rect 378042 39012 378048 39024
rect 377548 38984 378048 39012
rect 377548 38972 377554 38984
rect 378042 38972 378048 38984
rect 378100 38972 378106 39024
rect 378502 38972 378508 39024
rect 378560 39012 378566 39024
rect 379422 39012 379428 39024
rect 378560 38984 379428 39012
rect 378560 38972 378566 38984
rect 379422 38972 379428 38984
rect 379480 38972 379486 39024
rect 379514 38972 379520 39024
rect 379572 39012 379578 39024
rect 380710 39012 380716 39024
rect 379572 38984 380716 39012
rect 379572 38972 379578 38984
rect 380710 38972 380716 38984
rect 380768 38972 380774 39024
rect 382550 38972 382556 39024
rect 382608 39012 382614 39024
rect 383470 39012 383476 39024
rect 382608 38984 383476 39012
rect 382608 38972 382614 38984
rect 383470 38972 383476 38984
rect 383528 38972 383534 39024
rect 385586 38972 385592 39024
rect 385644 39012 385650 39024
rect 386322 39012 386328 39024
rect 385644 38984 386328 39012
rect 385644 38972 385650 38984
rect 386322 38972 386328 38984
rect 386380 38972 386386 39024
rect 386598 38972 386604 39024
rect 386656 39012 386662 39024
rect 387702 39012 387708 39024
rect 386656 38984 387708 39012
rect 386656 38972 386662 38984
rect 387702 38972 387708 38984
rect 387760 38972 387766 39024
rect 388622 38972 388628 39024
rect 388680 39012 388686 39024
rect 389082 39012 389088 39024
rect 388680 38984 389088 39012
rect 388680 38972 388686 38984
rect 389082 38972 389088 38984
rect 389140 38972 389146 39024
rect 389634 38972 389640 39024
rect 389692 39012 389698 39024
rect 390462 39012 390468 39024
rect 389692 38984 390468 39012
rect 389692 38972 389698 38984
rect 390462 38972 390468 38984
rect 390520 38972 390526 39024
rect 390646 38972 390652 39024
rect 390704 39012 390710 39024
rect 391750 39012 391756 39024
rect 390704 38984 391756 39012
rect 390704 38972 390710 38984
rect 391750 38972 391756 38984
rect 391808 38972 391814 39024
rect 392762 38972 392768 39024
rect 392820 39012 392826 39024
rect 393222 39012 393228 39024
rect 392820 38984 393228 39012
rect 392820 38972 392826 38984
rect 393222 38972 393228 38984
rect 393280 38972 393286 39024
rect 393774 38972 393780 39024
rect 393832 39012 393838 39024
rect 394602 39012 394608 39024
rect 393832 38984 394608 39012
rect 393832 38972 393838 38984
rect 394602 38972 394608 38984
rect 394660 38972 394666 39024
rect 396810 38972 396816 39024
rect 396868 39012 396874 39024
rect 397362 39012 397368 39024
rect 396868 38984 397368 39012
rect 396868 38972 396874 38984
rect 397362 38972 397368 38984
rect 397420 38972 397426 39024
rect 397822 38972 397828 39024
rect 397880 39012 397886 39024
rect 398742 39012 398748 39024
rect 397880 38984 398748 39012
rect 397880 38972 397886 38984
rect 398742 38972 398748 38984
rect 398800 38972 398806 39024
rect 398834 38972 398840 39024
rect 398892 39012 398898 39024
rect 400122 39012 400128 39024
rect 398892 38984 400128 39012
rect 398892 38972 398898 38984
rect 400122 38972 400128 38984
rect 400180 38972 400186 39024
rect 401870 38972 401876 39024
rect 401928 39012 401934 39024
rect 402882 39012 402888 39024
rect 401928 38984 402888 39012
rect 401928 38972 401934 38984
rect 402882 38972 402888 38984
rect 402940 38972 402946 39024
rect 404906 38972 404912 39024
rect 404964 39012 404970 39024
rect 405642 39012 405648 39024
rect 404964 38984 405648 39012
rect 404964 38972 404970 38984
rect 405642 38972 405648 38984
rect 405700 38972 405706 39024
rect 405918 38972 405924 39024
rect 405976 39012 405982 39024
rect 407022 39012 407028 39024
rect 405976 38984 407028 39012
rect 405976 38972 405982 38984
rect 407022 38972 407028 38984
rect 407080 38972 407086 39024
rect 409046 38972 409052 39024
rect 409104 39012 409110 39024
rect 409782 39012 409788 39024
rect 409104 38984 409788 39012
rect 409104 38972 409110 38984
rect 409782 38972 409788 38984
rect 409840 38972 409846 39024
rect 410058 38972 410064 39024
rect 410116 39012 410122 39024
rect 411070 39012 411076 39024
rect 410116 38984 411076 39012
rect 410116 38972 410122 38984
rect 411070 38972 411076 38984
rect 411128 38972 411134 39024
rect 412082 38972 412088 39024
rect 412140 39012 412146 39024
rect 412542 39012 412548 39024
rect 412140 38984 412548 39012
rect 412140 38972 412146 38984
rect 412542 38972 412548 38984
rect 412600 38972 412606 39024
rect 413094 38972 413100 39024
rect 413152 39012 413158 39024
rect 413922 39012 413928 39024
rect 413152 38984 413928 39012
rect 413152 38972 413158 38984
rect 413922 38972 413928 38984
rect 413980 38972 413986 39024
rect 414106 38972 414112 39024
rect 414164 39012 414170 39024
rect 415302 39012 415308 39024
rect 414164 38984 415308 39012
rect 414164 38972 414170 38984
rect 415302 38972 415308 38984
rect 415360 38972 415366 39024
rect 416130 38972 416136 39024
rect 416188 39012 416194 39024
rect 416682 39012 416688 39024
rect 416188 38984 416688 39012
rect 416188 38972 416194 38984
rect 416682 38972 416688 38984
rect 416740 38972 416746 39024
rect 417142 38972 417148 39024
rect 417200 39012 417206 39024
rect 418062 39012 418068 39024
rect 417200 38984 418068 39012
rect 417200 38972 417206 38984
rect 418062 38972 418068 38984
rect 418120 38972 418126 39024
rect 418154 38972 418160 39024
rect 418212 39012 418218 39024
rect 419350 39012 419356 39024
rect 418212 38984 419356 39012
rect 418212 38972 418218 38984
rect 419350 38972 419356 38984
rect 419408 38972 419414 39024
rect 421190 38972 421196 39024
rect 421248 39012 421254 39024
rect 422202 39012 422208 39024
rect 421248 38984 422208 39012
rect 421248 38972 421254 38984
rect 422202 38972 422208 38984
rect 422260 38972 422266 39024
rect 424318 38972 424324 39024
rect 424376 39012 424382 39024
rect 424962 39012 424968 39024
rect 424376 38984 424968 39012
rect 424376 38972 424382 38984
rect 424962 38972 424968 38984
rect 425020 38972 425026 39024
rect 425330 38972 425336 39024
rect 425388 39012 425394 39024
rect 426250 39012 426256 39024
rect 425388 38984 426256 39012
rect 425388 38972 425394 38984
rect 426250 38972 426256 38984
rect 426308 38972 426314 39024
rect 428366 38972 428372 39024
rect 428424 39012 428430 39024
rect 429102 39012 429108 39024
rect 428424 38984 429108 39012
rect 428424 38972 428430 38984
rect 429102 38972 429108 38984
rect 429160 38972 429166 39024
rect 429378 38972 429384 39024
rect 429436 39012 429442 39024
rect 430482 39012 430488 39024
rect 429436 38984 430488 39012
rect 429436 38972 429442 38984
rect 430482 38972 430488 38984
rect 430540 38972 430546 39024
rect 431402 38972 431408 39024
rect 431460 39012 431466 39024
rect 431862 39012 431868 39024
rect 431460 38984 431868 39012
rect 431460 38972 431466 38984
rect 431862 38972 431868 38984
rect 431920 38972 431926 39024
rect 432414 38972 432420 39024
rect 432472 39012 432478 39024
rect 433242 39012 433248 39024
rect 432472 38984 433248 39012
rect 432472 38972 432478 38984
rect 433242 38972 433248 38984
rect 433300 38972 433306 39024
rect 433426 38972 433432 39024
rect 433484 39012 433490 39024
rect 434622 39012 434628 39024
rect 433484 38984 434628 39012
rect 433484 38972 433490 38984
rect 434622 38972 434628 38984
rect 434680 38972 434686 39024
rect 435450 38972 435456 39024
rect 435508 39012 435514 39024
rect 436002 39012 436008 39024
rect 435508 38984 436008 39012
rect 435508 38972 435514 38984
rect 436002 38972 436008 38984
rect 436060 38972 436066 39024
rect 436462 38972 436468 39024
rect 436520 39012 436526 39024
rect 437382 39012 437388 39024
rect 436520 38984 437388 39012
rect 436520 38972 436526 38984
rect 437382 38972 437388 38984
rect 437440 38972 437446 39024
rect 439590 38972 439596 39024
rect 439648 39012 439654 39024
rect 440142 39012 440148 39024
rect 439648 38984 440148 39012
rect 439648 38972 439654 38984
rect 440142 38972 440148 38984
rect 440200 38972 440206 39024
rect 440602 38972 440608 39024
rect 440660 39012 440666 39024
rect 441522 39012 441528 39024
rect 440660 38984 441528 39012
rect 440660 38972 440666 38984
rect 441522 38972 441528 38984
rect 441580 38972 441586 39024
rect 441614 38972 441620 39024
rect 441672 39012 441678 39024
rect 442902 39012 442908 39024
rect 441672 38984 442908 39012
rect 441672 38972 441678 38984
rect 442902 38972 442908 38984
rect 442960 38972 442966 39024
rect 443638 38972 443644 39024
rect 443696 39012 443702 39024
rect 444282 39012 444288 39024
rect 443696 38984 444288 39012
rect 443696 38972 443702 38984
rect 444282 38972 444288 38984
rect 444340 38972 444346 39024
rect 447686 38972 447692 39024
rect 447744 39012 447750 39024
rect 448422 39012 448428 39024
rect 447744 38984 448428 39012
rect 447744 38972 447750 38984
rect 448422 38972 448428 38984
rect 448480 38972 448486 39024
rect 448698 38972 448704 39024
rect 448756 39012 448762 39024
rect 449802 39012 449808 39024
rect 448756 38984 449808 39012
rect 448756 38972 448762 38984
rect 449802 38972 449808 38984
rect 449860 38972 449866 39024
rect 450722 38972 450728 39024
rect 450780 39012 450786 39024
rect 451182 39012 451188 39024
rect 450780 38984 451188 39012
rect 450780 38972 450786 38984
rect 451182 38972 451188 38984
rect 451240 38972 451246 39024
rect 451734 38972 451740 39024
rect 451792 39012 451798 39024
rect 452562 39012 452568 39024
rect 451792 38984 452568 39012
rect 451792 38972 451798 38984
rect 452562 38972 452568 38984
rect 452620 38972 452626 39024
rect 452746 38972 452752 39024
rect 452804 39012 452810 39024
rect 453850 39012 453856 39024
rect 452804 38984 453856 39012
rect 452804 38972 452810 38984
rect 453850 38972 453856 38984
rect 453908 38972 453914 39024
rect 454862 38972 454868 39024
rect 454920 39012 454926 39024
rect 455322 39012 455328 39024
rect 454920 38984 455328 39012
rect 454920 38972 454926 38984
rect 455322 38972 455328 38984
rect 455380 38972 455386 39024
rect 456886 38972 456892 39024
rect 456944 39012 456950 39024
rect 457990 39012 457996 39024
rect 456944 38984 457996 39012
rect 456944 38972 456950 38984
rect 457990 38972 457996 38984
rect 458048 38972 458054 39024
rect 459922 38972 459928 39024
rect 459980 39012 459986 39024
rect 460842 39012 460848 39024
rect 459980 38984 460848 39012
rect 459980 38972 459986 38984
rect 460842 38972 460848 38984
rect 460900 38972 460906 39024
rect 460934 38972 460940 39024
rect 460992 39012 460998 39024
rect 462222 39012 462228 39024
rect 460992 38984 462228 39012
rect 460992 38972 460998 38984
rect 462222 38972 462228 38984
rect 462280 38972 462286 39024
rect 462958 38972 462964 39024
rect 463016 39012 463022 39024
rect 463602 39012 463608 39024
rect 463016 38984 463608 39012
rect 463016 38972 463022 38984
rect 463602 38972 463608 38984
rect 463660 38972 463666 39024
rect 467006 38972 467012 39024
rect 467064 39012 467070 39024
rect 467742 39012 467748 39024
rect 467064 38984 467748 39012
rect 467064 38972 467070 38984
rect 467742 38972 467748 38984
rect 467800 38972 467806 39024
rect 468018 38972 468024 39024
rect 468076 39012 468082 39024
rect 469030 39012 469036 39024
rect 468076 38984 469036 39012
rect 468076 38972 468082 38984
rect 469030 38972 469036 38984
rect 469088 38972 469094 39024
rect 471146 38972 471152 39024
rect 471204 39012 471210 39024
rect 471882 39012 471888 39024
rect 471204 38984 471888 39012
rect 471204 38972 471210 38984
rect 471882 38972 471888 38984
rect 471940 38972 471946 39024
rect 475194 38972 475200 39024
rect 475252 39012 475258 39024
rect 476022 39012 476028 39024
rect 475252 38984 476028 39012
rect 475252 38972 475258 38984
rect 476022 38972 476028 38984
rect 476080 38972 476086 39024
rect 476206 38972 476212 39024
rect 476264 39012 476270 39024
rect 477402 39012 477408 39024
rect 476264 38984 477408 39012
rect 476264 38972 476270 38984
rect 477402 38972 477408 38984
rect 477460 38972 477466 39024
rect 478230 38972 478236 39024
rect 478288 39012 478294 39024
rect 478782 39012 478788 39024
rect 478288 38984 478788 39012
rect 478288 38972 478294 38984
rect 478782 38972 478788 38984
rect 478840 38972 478846 39024
rect 479242 38972 479248 39024
rect 479300 39012 479306 39024
rect 480162 39012 480168 39024
rect 479300 38984 480168 39012
rect 479300 38972 479306 38984
rect 480162 38972 480168 38984
rect 480220 38972 480226 39024
rect 482278 38972 482284 39024
rect 482336 39012 482342 39024
rect 482922 39012 482928 39024
rect 482336 38984 482928 39012
rect 482336 38972 482342 38984
rect 482922 38972 482928 38984
rect 482980 38972 482986 39024
rect 484394 38972 484400 39024
rect 484452 39012 484458 39024
rect 485590 39012 485596 39024
rect 484452 38984 485596 39012
rect 484452 38972 484458 38984
rect 485590 38972 485596 38984
rect 485648 38972 485654 39024
rect 486418 38972 486424 39024
rect 486476 39012 486482 39024
rect 487062 39012 487068 39024
rect 486476 38984 487068 39012
rect 486476 38972 486482 38984
rect 487062 38972 487068 38984
rect 487120 38972 487126 39024
rect 487430 38972 487436 39024
rect 487488 39012 487494 39024
rect 488442 39012 488448 39024
rect 487488 38984 488448 39012
rect 487488 38972 487494 38984
rect 488442 38972 488448 38984
rect 488500 38972 488506 39024
rect 492490 38972 492496 39024
rect 492548 39012 492554 39024
rect 493318 39012 493324 39024
rect 492548 38984 493324 39012
rect 492548 38972 492554 38984
rect 493318 38972 493324 38984
rect 493376 38972 493382 39024
rect 494514 38972 494520 39024
rect 494572 39012 494578 39024
rect 495342 39012 495348 39024
rect 494572 38984 495348 39012
rect 494572 38972 494578 38984
rect 495342 38972 495348 38984
rect 495400 38972 495406 39024
rect 497550 38972 497556 39024
rect 497608 39012 497614 39024
rect 498102 39012 498108 39024
rect 497608 38984 498108 39012
rect 497608 38972 497614 38984
rect 498102 38972 498108 38984
rect 498160 38972 498166 39024
rect 502702 38972 502708 39024
rect 502760 39012 502766 39024
rect 503622 39012 503628 39024
rect 502760 38984 503628 39012
rect 502760 38972 502766 38984
rect 503622 38972 503628 38984
rect 503680 38972 503686 39024
rect 505738 38972 505744 39024
rect 505796 39012 505802 39024
rect 506382 39012 506388 39024
rect 505796 38984 506388 39012
rect 505796 38972 505802 38984
rect 506382 38972 506388 38984
rect 506440 38972 506446 39024
rect 506750 38972 506756 39024
rect 506808 39012 506814 39024
rect 507762 39012 507768 39024
rect 506808 38984 507768 39012
rect 506808 38972 506814 38984
rect 507762 38972 507768 38984
rect 507820 38972 507826 39024
rect 514938 38972 514944 39024
rect 514996 39012 515002 39024
rect 516042 39012 516048 39024
rect 514996 38984 516048 39012
rect 514996 38972 515002 38984
rect 516042 38972 516048 38984
rect 516100 38972 516106 39024
rect 517974 38972 517980 39024
rect 518032 39012 518038 39024
rect 518802 39012 518808 39024
rect 518032 38984 518808 39012
rect 518032 38972 518038 38984
rect 518802 38972 518808 38984
rect 518860 38972 518866 39024
rect 518986 38972 518992 39024
rect 519044 39012 519050 39024
rect 520182 39012 520188 39024
rect 519044 38984 520188 39012
rect 519044 38972 519050 38984
rect 520182 38972 520188 38984
rect 520240 38972 520246 39024
rect 522022 38972 522028 39024
rect 522080 39012 522086 39024
rect 522942 39012 522948 39024
rect 522080 38984 522948 39012
rect 522080 38972 522086 38984
rect 522942 38972 522948 38984
rect 523000 38972 523006 39024
rect 525058 38972 525064 39024
rect 525116 39012 525122 39024
rect 525702 39012 525708 39024
rect 525116 38984 525708 39012
rect 525116 38972 525122 38984
rect 525702 38972 525708 38984
rect 525760 38972 525766 39024
rect 529106 38972 529112 39024
rect 529164 39012 529170 39024
rect 529842 39012 529848 39024
rect 529164 38984 529848 39012
rect 529164 38972 529170 38984
rect 529842 38972 529848 38984
rect 529900 38972 529906 39024
rect 530210 38972 530216 39024
rect 530268 39012 530274 39024
rect 531222 39012 531228 39024
rect 530268 38984 531228 39012
rect 530268 38972 530274 38984
rect 531222 38972 531228 38984
rect 531280 38972 531286 39024
rect 533246 38972 533252 39024
rect 533304 39012 533310 39024
rect 533982 39012 533988 39024
rect 533304 38984 533988 39012
rect 533304 38972 533310 38984
rect 533982 38972 533988 38984
rect 534040 38972 534046 39024
rect 537294 38972 537300 39024
rect 537352 39012 537358 39024
rect 538122 39012 538128 39024
rect 537352 38984 538128 39012
rect 537352 38972 537358 38984
rect 538122 38972 538128 38984
rect 538180 38972 538186 39024
rect 540330 38972 540336 39024
rect 540388 39012 540394 39024
rect 545758 39012 545764 39024
rect 540388 38984 545764 39012
rect 540388 38972 540394 38984
rect 545758 38972 545764 38984
rect 545816 38972 545822 39024
rect 45462 38904 45468 38956
rect 45520 38944 45526 38956
rect 80054 38944 80060 38956
rect 45520 38916 80060 38944
rect 45520 38904 45526 38916
rect 80054 38904 80060 38916
rect 80112 38904 80118 38956
rect 88978 38904 88984 38956
rect 89036 38944 89042 38956
rect 115658 38944 115664 38956
rect 89036 38916 115664 38944
rect 89036 38904 89042 38916
rect 115658 38904 115664 38916
rect 115716 38904 115722 38956
rect 118602 38904 118608 38956
rect 118660 38944 118666 38956
rect 143166 38944 143172 38956
rect 118660 38916 143172 38944
rect 118660 38904 118666 38916
rect 143166 38904 143172 38916
rect 143224 38904 143230 38956
rect 154482 38904 154488 38956
rect 154540 38944 154546 38956
rect 174722 38944 174728 38956
rect 154540 38916 174728 38944
rect 154540 38904 154546 38916
rect 174722 38904 174728 38916
rect 174780 38904 174786 38956
rect 182082 38904 182088 38956
rect 182140 38944 182146 38956
rect 198182 38944 198188 38956
rect 182140 38916 198188 38944
rect 182140 38904 182146 38916
rect 198182 38904 198188 38916
rect 198240 38904 198246 38956
rect 252462 38904 252468 38956
rect 252520 38944 252526 38956
rect 258258 38944 258264 38956
rect 252520 38916 258264 38944
rect 252520 38904 252526 38916
rect 258258 38904 258264 38916
rect 258316 38904 258322 38956
rect 263502 38904 263508 38956
rect 263560 38944 263566 38956
rect 268378 38944 268384 38956
rect 263560 38916 268384 38944
rect 263560 38904 263566 38916
rect 268378 38904 268384 38916
rect 268436 38904 268442 38956
rect 270402 38904 270408 38956
rect 270460 38944 270466 38956
rect 274634 38944 274640 38956
rect 270460 38916 274640 38944
rect 270460 38904 270466 38916
rect 274634 38904 274640 38916
rect 274692 38904 274698 38956
rect 281442 38904 281448 38956
rect 281500 38944 281506 38956
rect 283650 38944 283656 38956
rect 281500 38916 283656 38944
rect 281500 38904 281506 38916
rect 283650 38904 283656 38916
rect 283708 38904 283714 38956
rect 288342 38904 288348 38956
rect 288400 38944 288406 38956
rect 289814 38944 289820 38956
rect 288400 38916 289820 38944
rect 288400 38904 288406 38916
rect 289814 38904 289820 38916
rect 289872 38904 289878 38956
rect 319438 38904 319444 38956
rect 319496 38944 319502 38956
rect 321646 38944 321652 38956
rect 319496 38916 321652 38944
rect 319496 38904 319502 38916
rect 321646 38904 321652 38916
rect 321704 38904 321710 38956
rect 394786 38904 394792 38956
rect 394844 38944 394850 38956
rect 395890 38944 395896 38956
rect 394844 38916 395896 38944
rect 394844 38904 394850 38916
rect 395890 38904 395896 38916
rect 395948 38904 395954 38956
rect 444650 38904 444656 38956
rect 444708 38944 444714 38956
rect 445662 38944 445668 38956
rect 444708 38916 445668 38944
rect 444708 38904 444714 38916
rect 445662 38904 445668 38916
rect 445720 38904 445726 38956
rect 463970 38904 463976 38956
rect 464028 38944 464034 38956
rect 464982 38944 464988 38956
rect 464028 38916 464988 38944
rect 464028 38904 464034 38916
rect 464982 38904 464988 38916
rect 465040 38904 465046 38956
rect 499666 38904 499672 38956
rect 499724 38944 499730 38956
rect 500770 38944 500776 38956
rect 499724 38916 500776 38944
rect 499724 38904 499730 38916
rect 500770 38904 500776 38916
rect 500828 38904 500834 38956
rect 32398 38836 32404 38888
rect 32456 38876 32462 38888
rect 66806 38876 66812 38888
rect 32456 38848 66812 38876
rect 32456 38836 32462 38848
rect 66806 38836 66812 38848
rect 66864 38836 66870 38888
rect 71038 38836 71044 38888
rect 71096 38876 71102 38888
rect 72970 38876 72976 38888
rect 71096 38848 72976 38876
rect 71096 38836 71102 38848
rect 72970 38836 72976 38848
rect 73028 38836 73034 38888
rect 73062 38836 73068 38888
rect 73120 38876 73126 38888
rect 94314 38876 94320 38888
rect 73120 38848 94320 38876
rect 73120 38836 73126 38848
rect 94314 38836 94320 38848
rect 94372 38836 94378 38888
rect 95878 38836 95884 38888
rect 95936 38876 95942 38888
rect 121822 38876 121828 38888
rect 95936 38848 121828 38876
rect 95936 38836 95942 38848
rect 121822 38836 121828 38848
rect 121880 38836 121886 38888
rect 125502 38836 125508 38888
rect 125560 38876 125566 38888
rect 149330 38876 149336 38888
rect 125560 38848 149336 38876
rect 125560 38836 125566 38848
rect 149330 38836 149336 38848
rect 149388 38836 149394 38888
rect 151722 38836 151728 38888
rect 151780 38876 151786 38888
rect 171686 38876 171692 38888
rect 151780 38848 171692 38876
rect 151780 38836 151786 38848
rect 171686 38836 171692 38848
rect 171744 38836 171750 38888
rect 186222 38836 186228 38888
rect 186280 38876 186286 38888
rect 201218 38876 201224 38888
rect 186280 38848 201224 38876
rect 186280 38836 186286 38848
rect 201218 38836 201224 38848
rect 201276 38836 201282 38888
rect 249702 38836 249708 38888
rect 249760 38876 249766 38888
rect 256234 38876 256240 38888
rect 249760 38848 256240 38876
rect 249760 38836 249766 38848
rect 256234 38836 256240 38848
rect 256292 38836 256298 38888
rect 262122 38836 262128 38888
rect 262180 38876 262186 38888
rect 267366 38876 267372 38888
rect 262180 38848 267372 38876
rect 262180 38836 262186 38848
rect 267366 38836 267372 38848
rect 267424 38836 267430 38888
rect 268930 38836 268936 38888
rect 268988 38876 268994 38888
rect 272518 38876 272524 38888
rect 268988 38848 272524 38876
rect 268988 38836 268994 38848
rect 272518 38836 272524 38848
rect 272576 38836 272582 38888
rect 273162 38836 273168 38888
rect 273220 38876 273226 38888
rect 276566 38876 276572 38888
rect 273220 38848 276572 38876
rect 273220 38836 273226 38848
rect 276566 38836 276572 38848
rect 276624 38836 276630 38888
rect 336734 38836 336740 38888
rect 336792 38876 336798 38888
rect 338758 38876 338764 38888
rect 336792 38848 338764 38876
rect 336792 38836 336798 38848
rect 338758 38836 338764 38848
rect 338816 38836 338822 38888
rect 536282 38836 536288 38888
rect 536340 38876 536346 38888
rect 536742 38876 536748 38888
rect 536340 38848 536748 38876
rect 536340 38836 536346 38848
rect 536742 38836 536748 38848
rect 536800 38836 536806 38888
rect 50338 38768 50344 38820
rect 50396 38808 50402 38820
rect 78030 38808 78036 38820
rect 50396 38780 78036 38808
rect 50396 38768 50402 38780
rect 78030 38768 78036 38780
rect 78088 38768 78094 38820
rect 80698 38768 80704 38820
rect 80756 38808 80762 38820
rect 103514 38808 103520 38820
rect 80756 38780 103520 38808
rect 80756 38768 80762 38780
rect 103514 38768 103520 38780
rect 103572 38768 103578 38820
rect 122742 38768 122748 38820
rect 122800 38808 122806 38820
rect 147214 38808 147220 38820
rect 122800 38780 147220 38808
rect 122800 38768 122806 38780
rect 147214 38768 147220 38780
rect 147272 38768 147278 38820
rect 157242 38768 157248 38820
rect 157300 38808 157306 38820
rect 176746 38808 176752 38820
rect 157300 38780 176752 38808
rect 157300 38768 157306 38780
rect 176746 38768 176752 38780
rect 176804 38768 176810 38820
rect 260650 38768 260656 38820
rect 260708 38808 260714 38820
rect 266354 38808 266360 38820
rect 260708 38780 266360 38808
rect 260708 38768 260714 38780
rect 266354 38768 266360 38780
rect 266412 38768 266418 38820
rect 362218 38768 362224 38820
rect 362276 38808 362282 38820
rect 362862 38808 362868 38820
rect 362276 38780 362868 38808
rect 362276 38768 362282 38780
rect 362862 38768 362868 38780
rect 362920 38768 362926 38820
rect 375374 38768 375380 38820
rect 375432 38808 375438 38820
rect 376570 38808 376576 38820
rect 375432 38780 376576 38808
rect 375432 38768 375438 38780
rect 376570 38768 376576 38780
rect 376628 38768 376634 38820
rect 381538 38768 381544 38820
rect 381596 38808 381602 38820
rect 382182 38808 382188 38820
rect 381596 38780 382188 38808
rect 381596 38768 381602 38780
rect 382182 38768 382188 38780
rect 382240 38768 382246 38820
rect 400858 38768 400864 38820
rect 400916 38808 400922 38820
rect 401502 38808 401508 38820
rect 400916 38780 401508 38808
rect 400916 38768 400922 38780
rect 401502 38768 401508 38780
rect 401560 38768 401566 38820
rect 420178 38768 420184 38820
rect 420236 38808 420242 38820
rect 420822 38808 420828 38820
rect 420236 38780 420828 38808
rect 420236 38768 420242 38780
rect 420822 38768 420828 38780
rect 420880 38768 420886 38820
rect 490466 38768 490472 38820
rect 490524 38808 490530 38820
rect 491202 38808 491208 38820
rect 490524 38780 491208 38808
rect 490524 38768 490530 38780
rect 491202 38768 491208 38780
rect 491260 38768 491266 38820
rect 521010 38768 521016 38820
rect 521068 38808 521074 38820
rect 521562 38808 521568 38820
rect 521068 38780 521568 38808
rect 521068 38768 521074 38780
rect 521562 38768 521568 38780
rect 521620 38768 521626 38820
rect 42058 38700 42064 38752
rect 42116 38740 42122 38752
rect 42116 38712 45554 38740
rect 42116 38700 42122 38712
rect 45526 38672 45554 38712
rect 46198 38700 46204 38752
rect 46256 38740 46262 38752
rect 59722 38740 59728 38752
rect 46256 38712 59728 38740
rect 46256 38700 46262 38712
rect 59722 38700 59728 38712
rect 59780 38700 59786 38752
rect 61378 38700 61384 38752
rect 61436 38740 61442 38752
rect 62758 38740 62764 38752
rect 61436 38712 62764 38740
rect 61436 38700 61442 38712
rect 62758 38700 62764 38712
rect 62816 38700 62822 38752
rect 81066 38740 81072 38752
rect 64846 38712 81072 38740
rect 54570 38672 54576 38684
rect 45526 38644 54576 38672
rect 54570 38632 54576 38644
rect 54628 38632 54634 38684
rect 57238 38632 57244 38684
rect 57296 38672 57302 38684
rect 64846 38672 64874 38712
rect 81066 38700 81072 38712
rect 81124 38700 81130 38752
rect 89070 38700 89076 38752
rect 89128 38740 89134 38752
rect 97350 38740 97356 38752
rect 89128 38712 97356 38740
rect 89128 38700 89134 38712
rect 97350 38700 97356 38712
rect 97408 38700 97414 38752
rect 106918 38700 106924 38752
rect 106976 38740 106982 38752
rect 124858 38740 124864 38752
rect 106976 38712 124864 38740
rect 106976 38700 106982 38712
rect 124858 38700 124864 38712
rect 124916 38700 124922 38752
rect 129734 38700 129740 38752
rect 129792 38740 129798 38752
rect 131942 38740 131948 38752
rect 129792 38712 131948 38740
rect 129792 38700 129798 38712
rect 131942 38700 131948 38712
rect 132000 38700 132006 38752
rect 146202 38700 146208 38752
rect 146260 38740 146266 38752
rect 155129 38743 155187 38749
rect 155129 38740 155141 38743
rect 146260 38712 155141 38740
rect 146260 38700 146266 38712
rect 155129 38709 155141 38712
rect 155175 38709 155187 38743
rect 155129 38703 155187 38709
rect 161382 38700 161388 38752
rect 161440 38740 161446 38752
rect 179874 38740 179880 38752
rect 161440 38712 179880 38740
rect 161440 38700 161446 38712
rect 179874 38700 179880 38712
rect 179932 38700 179938 38752
rect 280062 38700 280068 38752
rect 280120 38740 280126 38752
rect 282638 38740 282644 38752
rect 280120 38712 282644 38740
rect 280120 38700 280126 38712
rect 282638 38700 282644 38712
rect 282696 38700 282702 38752
rect 312262 38700 312268 38752
rect 312320 38740 312326 38752
rect 313458 38740 313464 38752
rect 312320 38712 313464 38740
rect 312320 38700 312326 38712
rect 313458 38700 313464 38712
rect 313516 38700 313522 38752
rect 472158 38700 472164 38752
rect 472216 38740 472222 38752
rect 473170 38740 473176 38752
rect 472216 38712 473176 38740
rect 472216 38700 472222 38712
rect 473170 38700 473176 38712
rect 473228 38700 473234 38752
rect 493502 38700 493508 38752
rect 493560 38740 493566 38752
rect 493962 38740 493968 38752
rect 493560 38712 493968 38740
rect 493560 38700 493566 38712
rect 493962 38700 493968 38712
rect 494020 38700 494026 38752
rect 57296 38644 64874 38672
rect 57296 38632 57302 38644
rect 71130 38632 71136 38684
rect 71188 38672 71194 38684
rect 88334 38672 88340 38684
rect 71188 38644 88340 38672
rect 71188 38632 71194 38644
rect 88334 38632 88340 38644
rect 88392 38632 88398 38684
rect 278682 38632 278688 38684
rect 278740 38672 278746 38684
rect 281626 38672 281632 38684
rect 278740 38644 281632 38672
rect 278740 38632 278746 38644
rect 281626 38632 281632 38644
rect 281684 38632 281690 38684
rect 41322 38360 41328 38412
rect 41380 38400 41386 38412
rect 77018 38400 77024 38412
rect 41380 38372 77024 38400
rect 41380 38360 41386 38372
rect 77018 38360 77024 38372
rect 77076 38360 77082 38412
rect 34422 38292 34428 38344
rect 34480 38332 34486 38344
rect 70854 38332 70860 38344
rect 34480 38304 70860 38332
rect 34480 38292 34486 38304
rect 70854 38292 70860 38304
rect 70912 38292 70918 38344
rect 4798 38224 4804 38276
rect 4856 38264 4862 38276
rect 42150 38264 42156 38276
rect 4856 38236 42156 38264
rect 4856 38224 4862 38236
rect 42150 38224 42156 38236
rect 42208 38224 42214 38276
rect 55122 38224 55128 38276
rect 55180 38264 55186 38276
rect 89254 38264 89260 38276
rect 55180 38236 89260 38264
rect 55180 38224 55186 38236
rect 89254 38224 89260 38236
rect 89312 38224 89318 38276
rect 91002 38224 91008 38276
rect 91060 38264 91066 38276
rect 119798 38264 119804 38276
rect 91060 38236 119804 38264
rect 91060 38224 91066 38236
rect 119798 38224 119804 38236
rect 119856 38224 119862 38276
rect 7558 38156 7564 38208
rect 7616 38196 7622 38208
rect 44450 38196 44456 38208
rect 7616 38168 44456 38196
rect 7616 38156 7622 38168
rect 44450 38156 44456 38168
rect 44508 38156 44514 38208
rect 48222 38156 48228 38208
rect 48280 38196 48286 38208
rect 83090 38196 83096 38208
rect 48280 38168 83096 38196
rect 48280 38156 48286 38168
rect 83090 38156 83096 38168
rect 83148 38156 83154 38208
rect 84102 38156 84108 38208
rect 84160 38196 84166 38208
rect 113634 38196 113640 38208
rect 84160 38168 113640 38196
rect 84160 38156 84166 38168
rect 113634 38156 113640 38168
rect 113692 38156 113698 38208
rect 30282 38088 30288 38140
rect 30340 38128 30346 38140
rect 67818 38128 67824 38140
rect 30340 38100 67824 38128
rect 30340 38088 30346 38100
rect 67818 38088 67824 38100
rect 67876 38088 67882 38140
rect 79962 38088 79968 38140
rect 80020 38128 80026 38140
rect 110598 38128 110604 38140
rect 80020 38100 110604 38128
rect 80020 38088 80026 38100
rect 110598 38088 110604 38100
rect 110656 38088 110662 38140
rect 130378 38088 130384 38140
rect 130436 38128 130442 38140
rect 152366 38128 152372 38140
rect 130436 38100 152372 38128
rect 130436 38088 130442 38100
rect 152366 38088 152372 38100
rect 152424 38088 152430 38140
rect 17862 38020 17868 38072
rect 17920 38060 17926 38072
rect 56594 38060 56600 38072
rect 17920 38032 56600 38060
rect 17920 38020 17926 38032
rect 56594 38020 56600 38032
rect 56652 38020 56658 38072
rect 59262 38020 59268 38072
rect 59320 38060 59326 38072
rect 92290 38060 92296 38072
rect 59320 38032 92296 38060
rect 59320 38020 59326 38032
rect 92290 38020 92296 38032
rect 92348 38020 92354 38072
rect 133782 38020 133788 38072
rect 133840 38060 133846 38072
rect 156414 38060 156420 38072
rect 133840 38032 156420 38060
rect 133840 38020 133846 38032
rect 156414 38020 156420 38032
rect 156472 38020 156478 38072
rect 22002 37952 22008 38004
rect 22060 37992 22066 38004
rect 60734 37992 60740 38004
rect 22060 37964 60740 37992
rect 22060 37952 22066 37964
rect 60734 37952 60740 37964
rect 60792 37952 60798 38004
rect 66162 37952 66168 38004
rect 66220 37992 66226 38004
rect 98362 37992 98368 38004
rect 66220 37964 98368 37992
rect 66220 37952 66226 37964
rect 98362 37952 98368 37964
rect 98420 37952 98426 38004
rect 129642 37952 129648 38004
rect 129700 37992 129706 38004
rect 153378 37992 153384 38004
rect 129700 37964 153384 37992
rect 129700 37952 129706 37964
rect 153378 37952 153384 37964
rect 153436 37952 153442 38004
rect 8202 37884 8208 37936
rect 8260 37924 8266 37936
rect 48498 37924 48504 37936
rect 8260 37896 48504 37924
rect 8260 37884 8266 37896
rect 48498 37884 48504 37896
rect 48556 37884 48562 37936
rect 52362 37884 52368 37936
rect 52420 37924 52426 37936
rect 86126 37924 86132 37936
rect 52420 37896 86132 37924
rect 52420 37884 52426 37896
rect 86126 37884 86132 37896
rect 86184 37884 86190 37936
rect 86862 37884 86868 37936
rect 86920 37924 86926 37936
rect 116670 37924 116676 37936
rect 86920 37896 116676 37924
rect 86920 37884 86926 37896
rect 116670 37884 116676 37896
rect 116728 37884 116734 37936
rect 126882 37884 126888 37936
rect 126940 37924 126946 37936
rect 150434 37924 150440 37936
rect 126940 37896 150440 37924
rect 126940 37884 126946 37896
rect 150434 37884 150440 37896
rect 150492 37884 150498 37936
rect 93118 37272 93124 37324
rect 93176 37312 93182 37324
rect 95326 37312 95332 37324
rect 93176 37284 95332 37312
rect 93176 37272 93182 37284
rect 95326 37272 95332 37284
rect 95384 37272 95390 37324
rect 104802 36592 104808 36644
rect 104860 36632 104866 36644
rect 129734 36632 129740 36644
rect 104860 36604 129740 36632
rect 104860 36592 104866 36604
rect 129734 36592 129740 36604
rect 129792 36592 129798 36644
rect 37182 36524 37188 36576
rect 37240 36564 37246 36576
rect 71774 36564 71780 36576
rect 37240 36536 71780 36564
rect 37240 36524 37246 36536
rect 71774 36524 71780 36536
rect 71832 36524 71838 36576
rect 97902 36524 97908 36576
rect 97960 36564 97966 36576
rect 125870 36564 125876 36576
rect 97960 36536 125876 36564
rect 97960 36524 97966 36536
rect 125870 36524 125876 36536
rect 125928 36524 125934 36576
rect 131022 36524 131028 36576
rect 131080 36564 131086 36576
rect 146938 36564 146944 36576
rect 131080 36536 146944 36564
rect 131080 36524 131086 36536
rect 146938 36524 146944 36536
rect 146996 36524 147002 36576
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 14458 33096 14464 33108
rect 3568 33068 14464 33096
rect 3568 33056 3574 33068
rect 14458 33056 14464 33068
rect 14516 33056 14522 33108
rect 555418 33056 555424 33108
rect 555476 33096 555482 33108
rect 580166 33096 580172 33108
rect 555476 33068 580172 33096
rect 555476 33056 555482 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 14550 32376 14556 32428
rect 14608 32416 14614 32428
rect 42794 32416 42800 32428
rect 14608 32388 42800 32416
rect 14608 32376 14614 32388
rect 42794 32376 42800 32388
rect 42852 32376 42858 32428
rect 51718 30268 51724 30320
rect 51776 30308 51782 30320
rect 52546 30308 52552 30320
rect 51776 30280 52552 30308
rect 51776 30268 51782 30280
rect 52546 30268 52552 30280
rect 52604 30268 52610 30320
rect 102042 26868 102048 26920
rect 102100 26908 102106 26920
rect 128354 26908 128360 26920
rect 102100 26880 128360 26908
rect 102100 26868 102106 26880
rect 128354 26868 128360 26880
rect 128412 26868 128418 26920
rect 551278 20612 551284 20664
rect 551336 20652 551342 20664
rect 579982 20652 579988 20664
rect 551336 20624 579988 20652
rect 551336 20612 551342 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 129458 8916 129464 8968
rect 129516 8956 129522 8968
rect 150618 8956 150624 8968
rect 129516 8928 150624 8956
rect 129516 8916 129522 8928
rect 150618 8916 150624 8928
rect 150676 8916 150682 8968
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 15838 6848 15844 6860
rect 3476 6820 15844 6848
rect 3476 6808 3482 6820
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 547138 6808 547144 6860
rect 547196 6848 547202 6860
rect 580166 6848 580172 6860
rect 547196 6820 580172 6848
rect 547196 6808 547202 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 562318 6196 562324 6248
rect 562376 6236 562382 6248
rect 572714 6236 572720 6248
rect 562376 6208 572720 6236
rect 562376 6196 562382 6208
rect 572714 6196 572720 6208
rect 572772 6196 572778 6248
rect 529842 6128 529848 6180
rect 529900 6168 529906 6180
rect 529900 6140 547874 6168
rect 529900 6128 529906 6140
rect 547846 6100 547874 6140
rect 565078 6128 565084 6180
rect 565136 6168 565142 6180
rect 576302 6168 576308 6180
rect 565136 6140 576308 6168
rect 565136 6128 565142 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 565630 6100 565636 6112
rect 547846 6072 565636 6100
rect 565630 6060 565636 6072
rect 565688 6060 565694 6112
rect 556798 5584 556804 5636
rect 556856 5624 556862 5636
rect 558546 5624 558552 5636
rect 556856 5596 558552 5624
rect 556856 5584 556862 5596
rect 558546 5584 558552 5596
rect 558604 5584 558610 5636
rect 560938 5584 560944 5636
rect 560996 5624 561002 5636
rect 569126 5624 569132 5636
rect 560996 5596 569132 5624
rect 560996 5584 561002 5596
rect 569126 5584 569132 5596
rect 569184 5584 569190 5636
rect 454678 5516 454684 5568
rect 454736 5556 454742 5568
rect 459186 5556 459192 5568
rect 454736 5528 459192 5556
rect 454736 5516 454742 5528
rect 459186 5516 459192 5528
rect 459244 5516 459250 5568
rect 558178 5516 558184 5568
rect 558236 5556 558242 5568
rect 562042 5556 562048 5568
rect 558236 5528 562048 5556
rect 558236 5516 558242 5528
rect 562042 5516 562048 5528
rect 562100 5516 562106 5568
rect 515398 5108 515404 5160
rect 515456 5148 515462 5160
rect 526622 5148 526628 5160
rect 515456 5120 526628 5148
rect 515456 5108 515462 5120
rect 526622 5108 526628 5120
rect 526680 5108 526686 5160
rect 487062 5040 487068 5092
rect 487120 5080 487126 5092
rect 515950 5080 515956 5092
rect 487120 5052 515956 5080
rect 487120 5040 487126 5052
rect 515950 5040 515956 5052
rect 516008 5040 516014 5092
rect 518158 5040 518164 5092
rect 518216 5080 518222 5092
rect 530118 5080 530124 5092
rect 518216 5052 530124 5080
rect 518216 5040 518222 5052
rect 530118 5040 530124 5052
rect 530176 5040 530182 5092
rect 465718 4972 465724 5024
rect 465776 5012 465782 5024
rect 480530 5012 480536 5024
rect 465776 4984 480536 5012
rect 465776 4972 465782 4984
rect 480530 4972 480536 4984
rect 480588 4972 480594 5024
rect 489822 4972 489828 5024
rect 489880 5012 489886 5024
rect 519538 5012 519544 5024
rect 489880 4984 519544 5012
rect 489880 4972 489886 4984
rect 519538 4972 519544 4984
rect 519596 4972 519602 5024
rect 443638 4904 443644 4956
rect 443696 4944 443702 4956
rect 455690 4944 455696 4956
rect 443696 4916 455696 4944
rect 443696 4904 443702 4916
rect 455690 4904 455696 4916
rect 455748 4904 455754 4956
rect 462130 4904 462136 4956
rect 462188 4944 462194 4956
rect 487614 4944 487620 4956
rect 462188 4916 487620 4944
rect 462188 4904 462194 4916
rect 487614 4904 487620 4916
rect 487672 4904 487678 4956
rect 493318 4904 493324 4956
rect 493376 4944 493382 4956
rect 523034 4944 523040 4956
rect 493376 4916 523040 4944
rect 493376 4904 493382 4916
rect 523034 4904 523040 4916
rect 523092 4904 523098 4956
rect 525058 4904 525064 4956
rect 525116 4944 525122 4956
rect 547874 4944 547880 4956
rect 525116 4916 547880 4944
rect 525116 4904 525122 4916
rect 547874 4904 547880 4916
rect 547932 4904 547938 4956
rect 429102 4836 429108 4888
rect 429160 4876 429166 4888
rect 448606 4876 448612 4888
rect 429160 4848 448612 4876
rect 429160 4836 429166 4848
rect 448606 4836 448612 4848
rect 448664 4836 448670 4888
rect 469030 4836 469036 4888
rect 469088 4876 469094 4888
rect 494698 4876 494704 4888
rect 469088 4848 494704 4876
rect 469088 4836 469094 4848
rect 494698 4836 494704 4848
rect 494756 4836 494762 4888
rect 505002 4836 505008 4888
rect 505060 4876 505066 4888
rect 537202 4876 537208 4888
rect 505060 4848 537208 4876
rect 505060 4836 505066 4848
rect 537202 4836 537208 4848
rect 537260 4836 537266 4888
rect 72602 4768 72608 4820
rect 72660 4808 72666 4820
rect 103698 4808 103704 4820
rect 72660 4780 103704 4808
rect 72660 4768 72666 4780
rect 103698 4768 103704 4780
rect 103756 4768 103762 4820
rect 139394 4768 139400 4820
rect 139452 4808 139458 4820
rect 158714 4808 158720 4820
rect 139452 4780 158720 4808
rect 139452 4768 139458 4780
rect 158714 4768 158720 4780
rect 158772 4768 158778 4820
rect 431862 4768 431868 4820
rect 431920 4808 431926 4820
rect 452102 4808 452108 4820
rect 431920 4780 452108 4808
rect 431920 4768 431926 4780
rect 452102 4768 452108 4780
rect 452160 4768 452166 4820
rect 471882 4768 471888 4820
rect 471940 4808 471946 4820
rect 498194 4808 498200 4820
rect 471940 4780 498200 4808
rect 471940 4768 471946 4780
rect 498194 4768 498200 4780
rect 498252 4768 498258 4820
rect 507670 4768 507676 4820
rect 507728 4808 507734 4820
rect 540790 4808 540796 4820
rect 507728 4780 540796 4808
rect 507728 4768 507734 4780
rect 540790 4768 540796 4780
rect 540848 4768 540854 4820
rect 62114 4632 62120 4684
rect 62172 4672 62178 4684
rect 64874 4672 64880 4684
rect 62172 4644 64880 4672
rect 62172 4632 62178 4644
rect 64874 4632 64880 4644
rect 64932 4632 64938 4684
rect 128354 4496 128360 4548
rect 128412 4536 128418 4548
rect 133966 4536 133972 4548
rect 128412 4508 133972 4536
rect 128412 4496 128418 4508
rect 133966 4496 133972 4508
rect 134024 4496 134030 4548
rect 502978 4156 502984 4208
rect 503036 4196 503042 4208
rect 505370 4196 505376 4208
rect 503036 4168 505376 4196
rect 503036 4156 503042 4168
rect 505370 4156 505376 4168
rect 505428 4156 505434 4208
rect 542998 4156 543004 4208
rect 543056 4196 543062 4208
rect 544378 4196 544384 4208
rect 543056 4168 544384 4196
rect 543056 4156 543062 4168
rect 544378 4156 544384 4168
rect 544436 4156 544442 4208
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 7558 4128 7564 4140
rect 2924 4100 7564 4128
rect 2924 4088 2930 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 50154 4088 50160 4140
rect 50212 4128 50218 4140
rect 50212 4100 55214 4128
rect 50212 4088 50218 4100
rect 41874 4020 41880 4072
rect 41932 4060 41938 4072
rect 50338 4060 50344 4072
rect 41932 4032 50344 4060
rect 41932 4020 41938 4032
rect 50338 4020 50344 4032
rect 50396 4020 50402 4072
rect 55186 4060 55214 4100
rect 348970 4088 348976 4140
rect 349028 4128 349034 4140
rect 355226 4128 355232 4140
rect 349028 4100 355232 4128
rect 349028 4088 349034 4100
rect 355226 4088 355232 4100
rect 355284 4088 355290 4140
rect 358722 4088 358728 4140
rect 358780 4128 358786 4140
rect 367002 4128 367008 4140
rect 358780 4100 367008 4128
rect 358780 4088 358786 4100
rect 367002 4088 367008 4100
rect 367060 4088 367066 4140
rect 380710 4088 380716 4140
rect 380768 4128 380774 4140
rect 391658 4128 391664 4140
rect 380768 4100 391664 4128
rect 380768 4088 380774 4100
rect 391658 4088 391664 4100
rect 391716 4088 391722 4140
rect 398742 4088 398748 4140
rect 398800 4128 398806 4140
rect 413094 4128 413100 4140
rect 398800 4100 413100 4128
rect 398800 4088 398806 4100
rect 413094 4088 413100 4100
rect 413152 4088 413158 4140
rect 413922 4088 413928 4140
rect 413980 4128 413986 4140
rect 430850 4128 430856 4140
rect 413980 4100 430856 4128
rect 413980 4088 413986 4100
rect 430850 4088 430856 4100
rect 430908 4088 430914 4140
rect 433242 4088 433248 4140
rect 433300 4128 433306 4140
rect 453298 4128 453304 4140
rect 433300 4100 453304 4128
rect 433300 4088 433306 4100
rect 453298 4088 453304 4100
rect 453356 4088 453362 4140
rect 455322 4088 455328 4140
rect 455380 4128 455386 4140
rect 479334 4128 479340 4140
rect 455380 4100 479340 4128
rect 455380 4088 455386 4100
rect 479334 4088 479340 4100
rect 479392 4088 479398 4140
rect 481542 4088 481548 4140
rect 481600 4128 481606 4140
rect 510062 4128 510068 4140
rect 481600 4100 510068 4128
rect 481600 4088 481606 4100
rect 510062 4088 510068 4100
rect 510120 4088 510126 4140
rect 518802 4088 518808 4140
rect 518860 4128 518866 4140
rect 552658 4128 552664 4140
rect 518860 4100 552664 4128
rect 518860 4088 518866 4100
rect 552658 4088 552664 4100
rect 552716 4088 552722 4140
rect 55186 4032 60044 4060
rect 20530 3952 20536 4004
rect 20588 3992 20594 4004
rect 46198 3992 46204 4004
rect 20588 3964 46204 3992
rect 20588 3952 20594 3964
rect 46198 3952 46204 3964
rect 46256 3952 46262 4004
rect 57146 3992 57152 4004
rect 50356 3964 57152 3992
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 42058 3924 42064 3936
rect 14792 3896 42064 3924
rect 14792 3884 14798 3896
rect 42058 3884 42064 3896
rect 42116 3884 42122 3936
rect 45370 3884 45376 3936
rect 45428 3924 45434 3936
rect 50356 3924 50384 3964
rect 57146 3952 57152 3964
rect 57204 3952 57210 4004
rect 60016 3992 60044 4032
rect 60826 4020 60832 4072
rect 60884 4060 60890 4072
rect 72418 4060 72424 4072
rect 60884 4032 72424 4060
rect 60884 4020 60890 4032
rect 72418 4020 72424 4032
rect 72476 4020 72482 4072
rect 82078 4020 82084 4072
rect 82136 4060 82142 4072
rect 84838 4060 84844 4072
rect 82136 4032 84844 4060
rect 82136 4020 82142 4032
rect 84838 4020 84844 4032
rect 84896 4020 84902 4072
rect 340690 4020 340696 4072
rect 340748 4060 340754 4072
rect 346946 4060 346952 4072
rect 340748 4032 346952 4060
rect 340748 4020 340754 4032
rect 346946 4020 346952 4032
rect 347004 4020 347010 4072
rect 361482 4020 361488 4072
rect 361540 4060 361546 4072
rect 370590 4060 370596 4072
rect 361540 4032 370596 4060
rect 361540 4020 361546 4032
rect 370590 4020 370596 4032
rect 370648 4020 370654 4072
rect 380802 4020 380808 4072
rect 380860 4060 380866 4072
rect 393038 4060 393044 4072
rect 380860 4032 393044 4060
rect 380860 4020 380866 4032
rect 393038 4020 393044 4032
rect 393096 4020 393102 4072
rect 395890 4020 395896 4072
rect 395948 4060 395954 4072
rect 409598 4060 409604 4072
rect 395948 4032 409604 4060
rect 395948 4020 395954 4032
rect 409598 4020 409604 4032
rect 409656 4020 409662 4072
rect 411162 4020 411168 4072
rect 411220 4060 411226 4072
rect 428458 4060 428464 4072
rect 411220 4032 428464 4060
rect 411220 4020 411226 4032
rect 428458 4020 428464 4032
rect 428516 4020 428522 4072
rect 430390 4020 430396 4072
rect 430448 4060 430454 4072
rect 450906 4060 450912 4072
rect 430448 4032 450912 4060
rect 430448 4020 430454 4032
rect 450906 4020 450912 4032
rect 450964 4020 450970 4072
rect 453942 4020 453948 4072
rect 454000 4060 454006 4072
rect 478138 4060 478144 4072
rect 454000 4032 478144 4060
rect 454000 4020 454006 4032
rect 478138 4020 478144 4032
rect 478196 4020 478202 4072
rect 485590 4020 485596 4072
rect 485648 4060 485654 4072
rect 513558 4060 513564 4072
rect 485648 4032 513564 4060
rect 485648 4020 485654 4032
rect 513558 4020 513564 4032
rect 513616 4020 513622 4072
rect 525702 4020 525708 4072
rect 525760 4060 525766 4072
rect 560846 4060 560852 4072
rect 525760 4032 560852 4060
rect 525760 4020 525766 4032
rect 560846 4020 560852 4032
rect 560904 4020 560910 4072
rect 68278 3992 68284 4004
rect 60016 3964 68284 3992
rect 68278 3952 68284 3964
rect 68336 3952 68342 4004
rect 92750 3952 92756 4004
rect 92808 3992 92814 4004
rect 95878 3992 95884 4004
rect 92808 3964 95884 3992
rect 92808 3952 92814 3964
rect 95878 3952 95884 3964
rect 95936 3952 95942 4004
rect 368290 3952 368296 4004
rect 368348 3992 368354 4004
rect 377674 3992 377680 4004
rect 368348 3964 377680 3992
rect 368348 3952 368354 3964
rect 377674 3952 377680 3964
rect 377732 3952 377738 4004
rect 379422 3952 379428 4004
rect 379480 3992 379486 4004
rect 390646 3992 390652 4004
rect 379480 3964 390652 3992
rect 379480 3952 379486 3964
rect 390646 3952 390652 3964
rect 390704 3952 390710 4004
rect 391750 3952 391756 4004
rect 391808 3992 391814 4004
rect 404814 3992 404820 4004
rect 391808 3964 404820 3992
rect 391808 3952 391814 3964
rect 404814 3952 404820 3964
rect 404872 3952 404878 4004
rect 405642 3952 405648 4004
rect 405700 3992 405706 4004
rect 421374 3992 421380 4004
rect 405700 3964 421380 3992
rect 405700 3952 405706 3964
rect 421374 3952 421380 3964
rect 421432 3952 421438 4004
rect 422202 3952 422208 4004
rect 422260 3992 422266 4004
rect 440326 3992 440332 4004
rect 422260 3964 440332 3992
rect 422260 3952 422266 3964
rect 440326 3952 440332 3964
rect 440384 3952 440390 4004
rect 441522 3952 441528 4004
rect 441580 3992 441586 4004
rect 462774 3992 462780 4004
rect 441580 3964 462780 3992
rect 441580 3952 441586 3964
rect 462774 3952 462780 3964
rect 462832 3952 462838 4004
rect 463602 3952 463608 4004
rect 463660 3992 463666 4004
rect 488810 3992 488816 4004
rect 463660 3964 488816 3992
rect 463660 3952 463666 3964
rect 488810 3952 488816 3964
rect 488868 3952 488874 4004
rect 491202 3952 491208 4004
rect 491260 3992 491266 4004
rect 520734 3992 520740 4004
rect 491260 3964 520740 3992
rect 491260 3952 491266 3964
rect 520734 3952 520740 3964
rect 520792 3952 520798 4004
rect 521562 3952 521568 4004
rect 521620 3992 521626 4004
rect 556154 3992 556160 4004
rect 521620 3964 556160 3992
rect 521620 3952 521626 3964
rect 556154 3952 556160 3964
rect 556212 3952 556218 4004
rect 45428 3896 50384 3924
rect 45428 3884 45434 3896
rect 52546 3884 52552 3936
rect 52604 3924 52610 3936
rect 53742 3924 53748 3936
rect 52604 3896 53748 3924
rect 52604 3884 52610 3896
rect 53742 3884 53748 3896
rect 53800 3884 53806 3936
rect 53837 3927 53895 3933
rect 53837 3893 53849 3927
rect 53883 3924 53895 3927
rect 75178 3924 75184 3936
rect 53883 3896 75184 3924
rect 53883 3893 53895 3896
rect 53837 3887 53895 3893
rect 75178 3884 75184 3896
rect 75236 3884 75242 3936
rect 343542 3884 343548 3936
rect 343600 3924 343606 3936
rect 349246 3924 349252 3936
rect 343600 3896 349252 3924
rect 343600 3884 343606 3896
rect 349246 3884 349252 3896
rect 349304 3884 349310 3936
rect 357342 3884 357348 3936
rect 357400 3924 357406 3936
rect 364610 3924 364616 3936
rect 357400 3896 364616 3924
rect 357400 3884 357406 3896
rect 364610 3884 364616 3896
rect 364668 3884 364674 3936
rect 369762 3884 369768 3936
rect 369820 3924 369826 3936
rect 379974 3924 379980 3936
rect 369820 3896 379980 3924
rect 369820 3884 369826 3896
rect 379974 3884 379980 3896
rect 380032 3884 380038 3936
rect 382182 3884 382188 3936
rect 382240 3924 382246 3936
rect 394234 3924 394240 3936
rect 382240 3896 394240 3924
rect 382240 3884 382246 3896
rect 394234 3884 394240 3896
rect 394292 3884 394298 3936
rect 397362 3884 397368 3936
rect 397420 3924 397426 3936
rect 411898 3924 411904 3936
rect 397420 3896 411904 3924
rect 397420 3884 397426 3896
rect 411898 3884 411904 3896
rect 411956 3884 411962 3936
rect 419350 3884 419356 3936
rect 419408 3924 419414 3936
rect 436738 3924 436744 3936
rect 419408 3896 436744 3924
rect 419408 3884 419414 3896
rect 436738 3884 436744 3896
rect 436796 3884 436802 3936
rect 438762 3884 438768 3936
rect 438820 3924 438826 3936
rect 460382 3924 460388 3936
rect 438820 3896 460388 3924
rect 438820 3884 438826 3896
rect 460382 3884 460388 3896
rect 460440 3884 460446 3936
rect 464982 3884 464988 3936
rect 465040 3924 465046 3936
rect 489914 3924 489920 3936
rect 465040 3896 489920 3924
rect 465040 3884 465046 3896
rect 489914 3884 489920 3896
rect 489972 3884 489978 3936
rect 493962 3884 493968 3936
rect 494020 3924 494026 3936
rect 524230 3924 524236 3936
rect 494020 3896 524236 3924
rect 494020 3884 494026 3896
rect 524230 3884 524236 3896
rect 524288 3884 524294 3936
rect 524322 3884 524328 3936
rect 524380 3924 524386 3936
rect 559742 3924 559748 3936
rect 524380 3896 559748 3924
rect 524380 3884 524386 3896
rect 559742 3884 559748 3896
rect 559800 3884 559806 3936
rect 32398 3816 32404 3868
rect 32456 3856 32462 3868
rect 64138 3856 64144 3868
rect 32456 3828 64144 3856
rect 32456 3816 32462 3828
rect 64138 3816 64144 3828
rect 64196 3816 64202 3868
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 80698 3856 80704 3868
rect 71556 3828 80704 3856
rect 71556 3816 71562 3828
rect 80698 3816 80704 3828
rect 80756 3816 80762 3868
rect 344922 3816 344928 3868
rect 344980 3856 344986 3868
rect 351638 3856 351644 3868
rect 344980 3828 351644 3856
rect 344980 3816 344986 3828
rect 351638 3816 351644 3828
rect 351696 3816 351702 3868
rect 351822 3816 351828 3868
rect 351880 3856 351886 3868
rect 358722 3856 358728 3868
rect 351880 3828 358728 3856
rect 351880 3816 351886 3828
rect 358722 3816 358728 3828
rect 358780 3816 358786 3868
rect 362862 3816 362868 3868
rect 362920 3856 362926 3868
rect 371694 3856 371700 3868
rect 362920 3828 371700 3856
rect 362920 3816 362926 3828
rect 371694 3816 371700 3828
rect 371752 3816 371758 3868
rect 372522 3816 372528 3868
rect 372580 3856 372586 3868
rect 382366 3856 382372 3868
rect 372580 3828 382372 3856
rect 372580 3816 372586 3828
rect 382366 3816 382372 3828
rect 382424 3816 382430 3868
rect 383562 3816 383568 3868
rect 383620 3856 383626 3868
rect 396534 3856 396540 3868
rect 383620 3828 396540 3856
rect 383620 3816 383626 3828
rect 396534 3816 396540 3828
rect 396592 3816 396598 3868
rect 401502 3816 401508 3868
rect 401560 3856 401566 3868
rect 416682 3856 416688 3868
rect 401560 3828 416688 3856
rect 401560 3816 401566 3828
rect 416682 3816 416688 3828
rect 416740 3816 416746 3868
rect 420822 3816 420828 3868
rect 420880 3856 420886 3868
rect 439130 3856 439136 3868
rect 420880 3828 439136 3856
rect 420880 3816 420886 3828
rect 439130 3816 439136 3828
rect 439188 3816 439194 3868
rect 442902 3816 442908 3868
rect 442960 3856 442966 3868
rect 463970 3856 463976 3868
rect 442960 3828 463976 3856
rect 442960 3816 442966 3828
rect 463970 3816 463976 3828
rect 464028 3816 464034 3868
rect 467742 3816 467748 3868
rect 467800 3856 467806 3868
rect 493502 3856 493508 3868
rect 467800 3828 493508 3856
rect 467800 3816 467806 3828
rect 493502 3816 493508 3828
rect 493560 3816 493566 3868
rect 495342 3816 495348 3868
rect 495400 3856 495406 3868
rect 525426 3856 525432 3868
rect 495400 3828 525432 3856
rect 495400 3816 495406 3828
rect 525426 3816 525432 3828
rect 525484 3816 525490 3868
rect 531222 3816 531228 3868
rect 531280 3856 531286 3868
rect 566826 3856 566832 3868
rect 531280 3828 566832 3856
rect 531280 3816 531286 3828
rect 566826 3816 566832 3828
rect 566884 3816 566890 3868
rect 35986 3748 35992 3800
rect 36044 3788 36050 3800
rect 71038 3788 71044 3800
rect 36044 3760 71044 3788
rect 36044 3748 36050 3760
rect 71038 3748 71044 3760
rect 71096 3748 71102 3800
rect 353202 3748 353208 3800
rect 353260 3788 353266 3800
rect 359918 3788 359924 3800
rect 353260 3760 359924 3788
rect 353260 3748 353266 3760
rect 359918 3748 359924 3760
rect 359976 3748 359982 3800
rect 360102 3748 360108 3800
rect 360160 3788 360166 3800
rect 368198 3788 368204 3800
rect 360160 3760 368204 3788
rect 360160 3748 360166 3760
rect 368198 3748 368204 3760
rect 368256 3748 368262 3800
rect 368382 3748 368388 3800
rect 368440 3788 368446 3800
rect 378870 3788 378876 3800
rect 368440 3760 378876 3788
rect 368440 3748 368446 3760
rect 378870 3748 378876 3760
rect 378928 3748 378934 3800
rect 383470 3748 383476 3800
rect 383528 3788 383534 3800
rect 395338 3788 395344 3800
rect 383528 3760 395344 3788
rect 383528 3748 383534 3760
rect 395338 3748 395344 3760
rect 395396 3748 395402 3800
rect 395982 3748 395988 3800
rect 396040 3788 396046 3800
rect 410794 3788 410800 3800
rect 396040 3760 410800 3788
rect 396040 3748 396046 3760
rect 410794 3748 410800 3760
rect 410852 3748 410858 3800
rect 415210 3748 415216 3800
rect 415268 3788 415274 3800
rect 433242 3788 433248 3800
rect 415268 3760 433248 3788
rect 415268 3748 415274 3760
rect 433242 3748 433248 3760
rect 433300 3748 433306 3800
rect 436002 3748 436008 3800
rect 436060 3788 436066 3800
rect 456886 3788 456892 3800
rect 436060 3760 456892 3788
rect 436060 3748 436066 3760
rect 456886 3748 456892 3760
rect 456944 3748 456950 3800
rect 457990 3748 457996 3800
rect 458048 3788 458054 3800
rect 481726 3788 481732 3800
rect 458048 3760 481732 3788
rect 458048 3748 458054 3760
rect 481726 3748 481732 3760
rect 481784 3748 481790 3800
rect 485682 3748 485688 3800
rect 485740 3788 485746 3800
rect 514754 3788 514760 3800
rect 485740 3760 514760 3788
rect 485740 3748 485746 3760
rect 514754 3748 514760 3760
rect 514812 3748 514818 3800
rect 527082 3748 527088 3800
rect 527140 3788 527146 3800
rect 563238 3788 563244 3800
rect 527140 3760 563244 3788
rect 527140 3748 527146 3760
rect 563238 3748 563244 3760
rect 563296 3748 563302 3800
rect 26510 3680 26516 3732
rect 26568 3720 26574 3732
rect 62114 3720 62120 3732
rect 26568 3692 62120 3720
rect 26568 3680 26574 3692
rect 62114 3680 62120 3692
rect 62172 3680 62178 3732
rect 64322 3680 64328 3732
rect 64380 3720 64386 3732
rect 89070 3720 89076 3732
rect 64380 3692 89076 3720
rect 64380 3680 64386 3692
rect 89070 3680 89076 3692
rect 89128 3680 89134 3732
rect 354582 3680 354588 3732
rect 354640 3720 354646 3732
rect 362310 3720 362316 3732
rect 354640 3692 362316 3720
rect 354640 3680 354646 3692
rect 362310 3680 362316 3692
rect 362368 3680 362374 3732
rect 365622 3680 365628 3732
rect 365680 3720 365686 3732
rect 375282 3720 375288 3732
rect 365680 3692 375288 3720
rect 365680 3680 365686 3692
rect 375282 3680 375288 3692
rect 375340 3680 375346 3732
rect 376662 3680 376668 3732
rect 376720 3720 376726 3732
rect 388254 3720 388260 3732
rect 376720 3692 388260 3720
rect 376720 3680 376726 3692
rect 388254 3680 388260 3692
rect 388312 3680 388318 3732
rect 393222 3680 393228 3732
rect 393280 3720 393286 3732
rect 407206 3720 407212 3732
rect 393280 3692 407212 3720
rect 393280 3680 393286 3692
rect 407206 3680 407212 3692
rect 407264 3680 407270 3732
rect 411070 3680 411076 3732
rect 411128 3720 411134 3732
rect 427262 3720 427268 3732
rect 411128 3692 427268 3720
rect 411128 3680 411134 3692
rect 427262 3680 427268 3692
rect 427320 3680 427326 3732
rect 427722 3680 427728 3732
rect 427780 3720 427786 3732
rect 447410 3720 447416 3732
rect 427780 3692 447416 3720
rect 427780 3680 427786 3692
rect 447410 3680 447416 3692
rect 447468 3680 447474 3732
rect 448422 3680 448428 3732
rect 448480 3720 448486 3732
rect 471054 3720 471060 3732
rect 448480 3692 471060 3720
rect 448480 3680 448486 3692
rect 471054 3680 471060 3692
rect 471112 3680 471118 3732
rect 473170 3680 473176 3732
rect 473228 3720 473234 3732
rect 499390 3720 499396 3732
rect 473228 3692 499396 3720
rect 473228 3680 473234 3692
rect 499390 3680 499396 3692
rect 499448 3680 499454 3732
rect 500862 3680 500868 3732
rect 500920 3720 500926 3732
rect 532510 3720 532516 3732
rect 500920 3692 532516 3720
rect 500920 3680 500926 3692
rect 532510 3680 532516 3692
rect 532568 3680 532574 3732
rect 533982 3680 533988 3732
rect 534040 3720 534046 3732
rect 570322 3720 570328 3732
rect 534040 3692 570328 3720
rect 534040 3680 534046 3692
rect 570322 3680 570328 3692
rect 570380 3680 570386 3732
rect 14550 3652 14556 3664
rect 6886 3624 14556 3652
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 6886 3584 6914 3624
rect 14550 3612 14556 3624
rect 14608 3612 14614 3664
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 75914 3652 75920 3664
rect 39632 3624 75920 3652
rect 39632 3612 39638 3624
rect 75914 3612 75920 3624
rect 75972 3612 75978 3664
rect 96246 3612 96252 3664
rect 96304 3652 96310 3664
rect 106918 3652 106924 3664
rect 96304 3624 106924 3652
rect 96304 3612 96310 3624
rect 106918 3612 106924 3624
rect 106976 3612 106982 3664
rect 108114 3612 108120 3664
rect 108172 3652 108178 3664
rect 128354 3652 128360 3664
rect 108172 3624 113174 3652
rect 108172 3612 108178 3624
rect 1728 3556 6914 3584
rect 1728 3544 1734 3556
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12308 3556 12572 3584
rect 12308 3544 12314 3556
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 4798 3516 4804 3528
rect 624 3488 4804 3516
rect 624 3476 630 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12342 3516 12348 3528
rect 11204 3488 12348 3516
rect 11204 3476 11210 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 12544 3516 12572 3556
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 16482 3584 16488 3596
rect 15988 3556 16488 3584
rect 15988 3544 15994 3556
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17862 3584 17868 3596
rect 17092 3556 17868 3584
rect 17092 3544 17098 3556
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 19242 3584 19248 3596
rect 18288 3556 19248 3584
rect 18288 3544 18294 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 20622 3584 20628 3596
rect 19484 3556 20628 3584
rect 19484 3544 19490 3556
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 61378 3584 61384 3596
rect 24268 3556 61384 3584
rect 24268 3544 24274 3556
rect 61378 3544 61384 3556
rect 61436 3544 61442 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 100754 3584 100760 3596
rect 69164 3556 100760 3584
rect 69164 3544 69170 3556
rect 100754 3544 100760 3556
rect 100812 3544 100818 3596
rect 107654 3584 107660 3596
rect 103486 3556 107660 3584
rect 12544 3488 47348 3516
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 45738 3448 45744 3460
rect 5316 3420 45744 3448
rect 5316 3408 5322 3420
rect 45738 3408 45744 3420
rect 45796 3408 45802 3460
rect 47320 3448 47348 3488
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 52362 3516 52368 3528
rect 51408 3488 52368 3516
rect 51408 3476 51414 3488
rect 52362 3476 52368 3488
rect 52420 3476 52426 3528
rect 53742 3476 53748 3528
rect 53800 3516 53806 3528
rect 53800 3488 65472 3516
rect 53800 3476 53806 3488
rect 51718 3448 51724 3460
rect 47320 3420 51724 3448
rect 51718 3408 51724 3420
rect 51776 3408 51782 3460
rect 56042 3408 56048 3460
rect 56100 3448 56106 3460
rect 56502 3448 56508 3460
rect 56100 3420 56508 3448
rect 56100 3408 56106 3420
rect 56502 3408 56508 3420
rect 56560 3408 56566 3460
rect 57238 3408 57244 3460
rect 57296 3448 57302 3460
rect 57882 3448 57888 3460
rect 57296 3420 57888 3448
rect 57296 3408 57302 3420
rect 57882 3408 57888 3420
rect 57940 3408 57946 3460
rect 58434 3408 58440 3460
rect 58492 3448 58498 3460
rect 59262 3448 59268 3460
rect 58492 3420 59268 3448
rect 58492 3408 58498 3420
rect 59262 3408 59268 3420
rect 59320 3408 59326 3460
rect 59630 3408 59636 3460
rect 59688 3448 59694 3460
rect 60642 3448 60648 3460
rect 59688 3420 60648 3448
rect 59688 3408 59694 3420
rect 60642 3408 60648 3420
rect 60700 3408 60706 3460
rect 62022 3408 62028 3460
rect 62080 3448 62086 3460
rect 65444 3448 65472 3488
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 66714 3476 66720 3528
rect 66772 3516 66778 3528
rect 67542 3516 67548 3528
rect 66772 3488 67548 3516
rect 66772 3476 66778 3488
rect 67542 3476 67548 3488
rect 67600 3476 67606 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 73798 3476 73804 3528
rect 73856 3516 73862 3528
rect 74442 3516 74448 3528
rect 73856 3488 74448 3516
rect 73856 3476 73862 3488
rect 74442 3476 74448 3488
rect 74500 3476 74506 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 77386 3476 77392 3528
rect 77444 3516 77450 3528
rect 78582 3516 78588 3528
rect 77444 3488 78588 3516
rect 77444 3476 77450 3488
rect 78582 3476 78588 3488
rect 78640 3476 78646 3528
rect 103486 3516 103514 3556
rect 107654 3544 107660 3556
rect 107712 3544 107718 3596
rect 111610 3544 111616 3596
rect 111668 3584 111674 3596
rect 113146 3584 113174 3624
rect 122806 3624 128360 3652
rect 122806 3584 122834 3624
rect 128354 3612 128360 3624
rect 128412 3612 128418 3664
rect 334618 3612 334624 3664
rect 334676 3652 334682 3664
rect 338666 3652 338672 3664
rect 334676 3624 338672 3652
rect 334676 3612 334682 3624
rect 338666 3612 338672 3624
rect 338724 3612 338730 3664
rect 364242 3612 364248 3664
rect 364300 3652 364306 3664
rect 372890 3652 372896 3664
rect 364300 3624 372896 3652
rect 364300 3612 364306 3624
rect 372890 3612 372896 3624
rect 372948 3612 372954 3664
rect 373902 3612 373908 3664
rect 373960 3652 373966 3664
rect 384758 3652 384764 3664
rect 373960 3624 384764 3652
rect 373960 3612 373966 3624
rect 384758 3612 384764 3624
rect 384816 3612 384822 3664
rect 386322 3612 386328 3664
rect 386380 3652 386386 3664
rect 398926 3652 398932 3664
rect 386380 3624 398932 3652
rect 386380 3612 386386 3624
rect 398926 3612 398932 3624
rect 398984 3612 398990 3664
rect 404262 3612 404268 3664
rect 404320 3652 404326 3664
rect 420178 3652 420184 3664
rect 404320 3624 420184 3652
rect 404320 3612 404326 3624
rect 420178 3612 420184 3624
rect 420236 3612 420242 3664
rect 426250 3612 426256 3664
rect 426308 3652 426314 3664
rect 445018 3652 445024 3664
rect 426308 3624 445024 3652
rect 426308 3612 426314 3624
rect 445018 3612 445024 3624
rect 445076 3612 445082 3664
rect 445662 3612 445668 3664
rect 445720 3652 445726 3664
rect 467466 3652 467472 3664
rect 445720 3624 467472 3652
rect 445720 3612 445726 3624
rect 467466 3612 467472 3624
rect 467524 3612 467530 3664
rect 469122 3612 469128 3664
rect 469180 3652 469186 3664
rect 495894 3652 495900 3664
rect 469180 3624 495900 3652
rect 469180 3612 469186 3624
rect 495894 3612 495900 3624
rect 495952 3612 495958 3664
rect 496722 3612 496728 3664
rect 496780 3652 496786 3664
rect 527818 3652 527824 3664
rect 496780 3624 527824 3652
rect 496780 3612 496786 3624
rect 527818 3612 527824 3624
rect 527876 3612 527882 3664
rect 536742 3612 536748 3664
rect 536800 3652 536806 3664
rect 573910 3652 573916 3664
rect 536800 3624 573916 3652
rect 536800 3612 536806 3624
rect 573910 3612 573916 3624
rect 573968 3612 573974 3664
rect 137278 3584 137284 3596
rect 111668 3556 111840 3584
rect 113146 3556 122834 3584
rect 123404 3556 137284 3584
rect 111668 3544 111674 3556
rect 78692 3488 103514 3516
rect 71130 3448 71136 3460
rect 62080 3420 64874 3448
rect 65444 3420 71136 3448
rect 62080 3408 62086 3420
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 28902 3380 28908 3392
rect 27764 3352 28908 3380
rect 27764 3340 27770 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 34422 3380 34428 3392
rect 33652 3352 34428 3380
rect 33652 3340 33658 3352
rect 34422 3340 34428 3352
rect 34480 3340 34486 3392
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 39298 3380 39304 3392
rect 38436 3352 39304 3380
rect 38436 3340 38442 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 43070 3340 43076 3392
rect 43128 3380 43134 3392
rect 44082 3380 44088 3392
rect 43128 3352 44088 3380
rect 43128 3340 43134 3352
rect 44082 3340 44088 3352
rect 44140 3340 44146 3392
rect 44266 3340 44272 3392
rect 44324 3380 44330 3392
rect 45462 3380 45468 3392
rect 44324 3352 45468 3380
rect 44324 3340 44330 3352
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 46658 3340 46664 3392
rect 46716 3380 46722 3392
rect 53837 3383 53895 3389
rect 53837 3380 53849 3383
rect 46716 3352 53849 3380
rect 46716 3340 46722 3352
rect 53837 3349 53849 3352
rect 53883 3349 53895 3383
rect 53837 3343 53895 3349
rect 64846 3312 64874 3420
rect 71130 3408 71136 3420
rect 71188 3408 71194 3460
rect 76190 3340 76196 3392
rect 76248 3380 76254 3392
rect 78692 3380 78720 3488
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 106182 3516 106188 3528
rect 105780 3488 106188 3516
rect 105780 3476 105786 3488
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 110322 3516 110328 3528
rect 109368 3488 110328 3516
rect 109368 3476 109374 3488
rect 110322 3476 110328 3488
rect 110380 3476 110386 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111702 3516 111708 3528
rect 110564 3488 111708 3516
rect 110564 3476 110570 3488
rect 111702 3476 111708 3488
rect 111760 3476 111766 3528
rect 111812 3516 111840 3556
rect 123404 3516 123432 3556
rect 137278 3544 137284 3556
rect 137336 3544 137342 3596
rect 267734 3544 267740 3596
rect 267792 3584 267798 3596
rect 268930 3584 268936 3596
rect 267792 3556 268936 3584
rect 267792 3544 267798 3556
rect 268930 3544 268936 3556
rect 268988 3544 268994 3596
rect 307754 3544 307760 3596
rect 307812 3584 307818 3596
rect 309042 3584 309048 3596
rect 307812 3556 309048 3584
rect 307812 3544 307818 3556
rect 309042 3544 309048 3556
rect 309100 3544 309106 3596
rect 328362 3544 328368 3596
rect 328420 3584 328426 3596
rect 331582 3584 331588 3596
rect 328420 3556 331588 3584
rect 328420 3544 328426 3556
rect 331582 3544 331588 3556
rect 331640 3544 331646 3596
rect 336642 3544 336648 3596
rect 336700 3584 336706 3596
rect 340966 3584 340972 3596
rect 336700 3556 340972 3584
rect 336700 3544 336706 3556
rect 340966 3544 340972 3556
rect 341024 3544 341030 3596
rect 357250 3544 357256 3596
rect 357308 3584 357314 3596
rect 365806 3584 365812 3596
rect 357308 3556 365812 3584
rect 357308 3544 357314 3556
rect 365806 3544 365812 3556
rect 365864 3544 365870 3596
rect 366910 3544 366916 3596
rect 366968 3584 366974 3596
rect 376478 3584 376484 3596
rect 366968 3556 376484 3584
rect 366968 3544 366974 3556
rect 376478 3544 376484 3556
rect 376536 3544 376542 3596
rect 376570 3544 376576 3596
rect 376628 3584 376634 3596
rect 387150 3584 387156 3596
rect 376628 3556 387156 3584
rect 376628 3544 376634 3556
rect 387150 3544 387156 3556
rect 387208 3544 387214 3596
rect 387610 3544 387616 3596
rect 387668 3584 387674 3596
rect 401318 3584 401324 3596
rect 387668 3556 401324 3584
rect 387668 3544 387674 3556
rect 401318 3544 401324 3556
rect 401376 3544 401382 3596
rect 402790 3544 402796 3596
rect 402848 3584 402854 3596
rect 418982 3584 418988 3596
rect 402848 3556 418988 3584
rect 402848 3544 402854 3556
rect 418982 3544 418988 3556
rect 419040 3544 419046 3596
rect 419442 3544 419448 3596
rect 419500 3584 419506 3596
rect 437934 3584 437940 3596
rect 419500 3556 437940 3584
rect 419500 3544 419506 3556
rect 437934 3544 437940 3556
rect 437992 3544 437998 3596
rect 442810 3544 442816 3596
rect 442868 3584 442874 3596
rect 465166 3584 465172 3596
rect 442868 3556 465172 3584
rect 442868 3544 442874 3556
rect 465166 3544 465172 3556
rect 465224 3544 465230 3596
rect 473262 3544 473268 3596
rect 473320 3584 473326 3596
rect 500586 3584 500592 3596
rect 473320 3556 500592 3584
rect 473320 3544 473326 3556
rect 500586 3544 500592 3556
rect 500644 3544 500650 3596
rect 500770 3544 500776 3596
rect 500828 3584 500834 3596
rect 531314 3584 531320 3596
rect 500828 3556 531320 3584
rect 500828 3544 500834 3556
rect 531314 3544 531320 3556
rect 531372 3544 531378 3596
rect 538122 3544 538128 3596
rect 538180 3584 538186 3596
rect 575106 3584 575112 3596
rect 538180 3556 575112 3584
rect 538180 3544 538186 3556
rect 575106 3544 575112 3556
rect 575164 3544 575170 3596
rect 111812 3488 123432 3516
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126882 3516 126888 3528
rect 125928 3488 126888 3516
rect 125928 3476 125934 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
rect 128170 3476 128176 3528
rect 128228 3516 128234 3528
rect 130378 3516 130384 3528
rect 128228 3488 130384 3516
rect 128228 3476 128234 3488
rect 130378 3476 130384 3488
rect 130436 3476 130442 3528
rect 130562 3476 130568 3528
rect 130620 3516 130626 3528
rect 131022 3516 131028 3528
rect 130620 3488 131028 3516
rect 130620 3476 130626 3488
rect 131022 3476 131028 3488
rect 131080 3476 131086 3528
rect 131758 3476 131764 3528
rect 131816 3516 131822 3528
rect 132402 3516 132408 3528
rect 131816 3488 132408 3516
rect 131816 3476 131822 3488
rect 132402 3476 132408 3488
rect 132460 3476 132466 3528
rect 132954 3476 132960 3528
rect 133012 3516 133018 3528
rect 133782 3516 133788 3528
rect 133012 3488 133788 3516
rect 133012 3476 133018 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
rect 134150 3476 134156 3528
rect 134208 3516 134214 3528
rect 135162 3516 135168 3528
rect 134208 3488 135168 3516
rect 134208 3476 134214 3488
rect 135162 3476 135168 3488
rect 135220 3476 135226 3528
rect 135254 3476 135260 3528
rect 135312 3516 135318 3528
rect 136542 3516 136548 3528
rect 135312 3488 136548 3516
rect 135312 3476 135318 3488
rect 136542 3476 136548 3488
rect 136600 3476 136606 3528
rect 138842 3476 138848 3528
rect 138900 3516 138906 3528
rect 139302 3516 139308 3528
rect 138900 3488 139308 3516
rect 138900 3476 138906 3488
rect 139302 3476 139308 3488
rect 139360 3476 139366 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 140682 3516 140688 3528
rect 140096 3488 140688 3516
rect 140096 3476 140102 3488
rect 140682 3476 140688 3488
rect 140740 3476 140746 3528
rect 141234 3476 141240 3528
rect 141292 3516 141298 3528
rect 142062 3516 142068 3528
rect 141292 3488 142068 3516
rect 141292 3476 141298 3488
rect 142062 3476 142068 3488
rect 142120 3476 142126 3528
rect 142430 3476 142436 3528
rect 142488 3516 142494 3528
rect 143442 3516 143448 3528
rect 142488 3488 143448 3516
rect 142488 3476 142494 3488
rect 143442 3476 143448 3488
rect 143500 3476 143506 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
rect 150342 3516 150348 3528
rect 149572 3488 150348 3516
rect 149572 3476 149578 3488
rect 150342 3476 150348 3488
rect 150400 3476 150406 3528
rect 150618 3476 150624 3528
rect 150676 3516 150682 3528
rect 151722 3516 151728 3528
rect 150676 3488 151728 3516
rect 150676 3476 150682 3488
rect 151722 3476 151728 3488
rect 151780 3476 151786 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 153102 3516 153108 3528
rect 151872 3488 153108 3516
rect 151872 3476 151878 3488
rect 153102 3476 153108 3488
rect 153160 3476 153166 3528
rect 155402 3476 155408 3528
rect 155460 3516 155466 3528
rect 155862 3516 155868 3528
rect 155460 3488 155868 3516
rect 155460 3476 155466 3488
rect 155862 3476 155868 3488
rect 155920 3476 155926 3528
rect 156598 3476 156604 3528
rect 156656 3516 156662 3528
rect 157242 3516 157248 3528
rect 156656 3488 157248 3516
rect 156656 3476 156662 3488
rect 157242 3476 157248 3488
rect 157300 3476 157306 3528
rect 157794 3476 157800 3528
rect 157852 3516 157858 3528
rect 158622 3516 158628 3528
rect 157852 3488 158628 3516
rect 157852 3476 157858 3488
rect 158622 3476 158628 3488
rect 158680 3476 158686 3528
rect 158898 3476 158904 3528
rect 158956 3516 158962 3528
rect 160002 3516 160008 3528
rect 158956 3488 160008 3516
rect 158956 3476 158962 3488
rect 160002 3476 160008 3488
rect 160060 3476 160066 3528
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161382 3516 161388 3528
rect 160152 3488 161388 3516
rect 160152 3476 160158 3488
rect 161382 3476 161388 3488
rect 161440 3476 161446 3528
rect 163682 3476 163688 3528
rect 163740 3516 163746 3528
rect 164142 3516 164148 3528
rect 163740 3488 164148 3516
rect 163740 3476 163746 3488
rect 164142 3476 164148 3488
rect 164200 3476 164206 3528
rect 166074 3476 166080 3528
rect 166132 3516 166138 3528
rect 166902 3516 166908 3528
rect 166132 3488 166908 3516
rect 166132 3476 166138 3488
rect 166902 3476 166908 3488
rect 166960 3476 166966 3528
rect 167178 3476 167184 3528
rect 167236 3516 167242 3528
rect 168282 3516 168288 3528
rect 167236 3488 168288 3516
rect 167236 3476 167242 3488
rect 168282 3476 168288 3488
rect 168340 3476 168346 3528
rect 168374 3476 168380 3528
rect 168432 3516 168438 3528
rect 169478 3516 169484 3528
rect 168432 3488 169484 3516
rect 168432 3476 168438 3488
rect 169478 3476 169484 3488
rect 169536 3476 169542 3528
rect 171962 3476 171968 3528
rect 172020 3516 172026 3528
rect 172422 3516 172428 3528
rect 172020 3488 172428 3516
rect 172020 3476 172026 3488
rect 172422 3476 172428 3488
rect 172480 3476 172486 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173802 3516 173808 3528
rect 173216 3488 173808 3516
rect 173216 3476 173222 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 174262 3476 174268 3528
rect 174320 3516 174326 3528
rect 175182 3516 175188 3528
rect 174320 3488 175188 3516
rect 174320 3476 174326 3488
rect 175182 3476 175188 3488
rect 175240 3476 175246 3528
rect 175458 3476 175464 3528
rect 175516 3516 175522 3528
rect 176562 3516 176568 3528
rect 175516 3488 176568 3516
rect 175516 3476 175522 3488
rect 176562 3476 176568 3488
rect 176620 3476 176626 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177758 3516 177764 3528
rect 176712 3488 177764 3516
rect 176712 3476 176718 3488
rect 177758 3476 177764 3488
rect 177816 3476 177822 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180702 3516 180708 3528
rect 180300 3488 180708 3516
rect 180300 3476 180306 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 181438 3476 181444 3528
rect 181496 3516 181502 3528
rect 182082 3516 182088 3528
rect 181496 3488 182088 3516
rect 181496 3476 181502 3488
rect 182082 3476 182088 3488
rect 182140 3476 182146 3528
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 184934 3476 184940 3528
rect 184992 3516 184998 3528
rect 186222 3516 186228 3528
rect 184992 3488 186228 3516
rect 184992 3476 184998 3488
rect 186222 3476 186228 3488
rect 186280 3476 186286 3528
rect 188522 3476 188528 3528
rect 188580 3516 188586 3528
rect 188982 3516 188988 3528
rect 188580 3488 188988 3516
rect 188580 3476 188586 3488
rect 188982 3476 188988 3488
rect 189040 3476 189046 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 191742 3516 191748 3528
rect 190880 3488 191748 3516
rect 190880 3476 190886 3488
rect 191742 3476 191748 3488
rect 191800 3476 191806 3528
rect 192018 3476 192024 3528
rect 192076 3516 192082 3528
rect 193122 3516 193128 3528
rect 192076 3488 193128 3516
rect 192076 3476 192082 3488
rect 193122 3476 193128 3488
rect 193180 3476 193186 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194318 3516 194324 3528
rect 193272 3488 194324 3516
rect 193272 3476 193278 3488
rect 194318 3476 194324 3488
rect 194376 3476 194382 3528
rect 197906 3476 197912 3528
rect 197964 3516 197970 3528
rect 198642 3516 198648 3528
rect 197964 3488 198648 3516
rect 197964 3476 197970 3488
rect 198642 3476 198648 3488
rect 198700 3476 198706 3528
rect 199102 3476 199108 3528
rect 199160 3516 199166 3528
rect 200022 3516 200028 3528
rect 199160 3488 200028 3516
rect 199160 3476 199166 3488
rect 200022 3476 200028 3488
rect 200080 3476 200086 3528
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 202782 3516 202788 3528
rect 201552 3488 202788 3516
rect 201552 3476 201558 3488
rect 202782 3476 202788 3488
rect 202840 3476 202846 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 205542 3516 205548 3528
rect 205140 3488 205548 3516
rect 205140 3476 205146 3488
rect 205542 3476 205548 3488
rect 205600 3476 205606 3528
rect 206186 3476 206192 3528
rect 206244 3516 206250 3528
rect 206922 3516 206928 3528
rect 206244 3488 206928 3516
rect 206244 3476 206250 3488
rect 206922 3476 206928 3488
rect 206980 3476 206986 3528
rect 207382 3476 207388 3528
rect 207440 3516 207446 3528
rect 208302 3516 208308 3528
rect 207440 3488 208308 3516
rect 207440 3476 207446 3488
rect 208302 3476 208308 3488
rect 208360 3476 208366 3528
rect 209774 3476 209780 3528
rect 209832 3516 209838 3528
rect 211062 3516 211068 3528
rect 209832 3488 211068 3516
rect 209832 3476 209838 3488
rect 211062 3476 211068 3488
rect 211120 3476 211126 3528
rect 213362 3476 213368 3528
rect 213420 3516 213426 3528
rect 213822 3516 213828 3528
rect 213420 3488 213828 3516
rect 213420 3476 213426 3488
rect 213822 3476 213828 3488
rect 213880 3476 213886 3528
rect 214466 3476 214472 3528
rect 214524 3516 214530 3528
rect 215202 3516 215208 3528
rect 214524 3488 215208 3516
rect 214524 3476 214530 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 216582 3516 216588 3528
rect 215720 3488 216588 3516
rect 215720 3476 215726 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 216858 3476 216864 3528
rect 216916 3516 216922 3528
rect 217962 3516 217968 3528
rect 216916 3488 217968 3516
rect 216916 3476 216922 3488
rect 217962 3476 217968 3488
rect 218020 3476 218026 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 219158 3516 219164 3528
rect 218112 3488 219164 3516
rect 218112 3476 218118 3488
rect 219158 3476 219164 3488
rect 219216 3476 219222 3528
rect 222746 3476 222752 3528
rect 222804 3516 222810 3528
rect 223482 3516 223488 3528
rect 222804 3488 223488 3516
rect 222804 3476 222810 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 224862 3516 224868 3528
rect 224000 3488 224868 3516
rect 224000 3476 224006 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 227622 3516 227628 3528
rect 226392 3488 227628 3516
rect 226392 3476 226398 3488
rect 227622 3476 227628 3488
rect 227680 3476 227686 3528
rect 229830 3476 229836 3528
rect 229888 3516 229894 3528
rect 230382 3516 230388 3528
rect 229888 3488 230388 3516
rect 229888 3476 229894 3488
rect 230382 3476 230388 3488
rect 230440 3476 230446 3528
rect 231026 3476 231032 3528
rect 231084 3516 231090 3528
rect 231762 3516 231768 3528
rect 231084 3488 231768 3516
rect 231084 3476 231090 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 234614 3476 234620 3528
rect 234672 3516 234678 3528
rect 235902 3516 235908 3528
rect 234672 3488 235908 3516
rect 234672 3476 234678 3488
rect 235902 3476 235908 3488
rect 235960 3476 235966 3528
rect 238110 3476 238116 3528
rect 238168 3516 238174 3528
rect 238662 3516 238668 3528
rect 238168 3488 238668 3516
rect 238168 3476 238174 3488
rect 238662 3476 238668 3488
rect 238720 3476 238726 3528
rect 239306 3476 239312 3528
rect 239364 3516 239370 3528
rect 240042 3516 240048 3528
rect 239364 3488 240048 3516
rect 239364 3476 239370 3488
rect 240042 3476 240048 3488
rect 240100 3476 240106 3528
rect 240502 3476 240508 3528
rect 240560 3516 240566 3528
rect 241422 3516 241428 3528
rect 240560 3488 241428 3516
rect 240560 3476 240566 3488
rect 241422 3476 241428 3488
rect 241480 3476 241486 3528
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 243998 3516 244004 3528
rect 242952 3488 244004 3516
rect 242952 3476 242958 3488
rect 243998 3476 244004 3488
rect 244056 3476 244062 3528
rect 247586 3476 247592 3528
rect 247644 3516 247650 3528
rect 248322 3516 248328 3528
rect 247644 3488 248328 3516
rect 247644 3476 247650 3488
rect 248322 3476 248328 3488
rect 248380 3476 248386 3528
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 251082 3516 251088 3528
rect 250036 3488 251088 3516
rect 250036 3476 250042 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 251174 3476 251180 3528
rect 251232 3516 251238 3528
rect 252462 3516 252468 3528
rect 251232 3488 252468 3516
rect 251232 3476 251238 3488
rect 252462 3476 252468 3488
rect 252520 3476 252526 3528
rect 254670 3476 254676 3528
rect 254728 3516 254734 3528
rect 255222 3516 255228 3528
rect 254728 3488 255228 3516
rect 254728 3476 254734 3488
rect 255222 3476 255228 3488
rect 255280 3476 255286 3528
rect 255866 3476 255872 3528
rect 255924 3516 255930 3528
rect 256602 3516 256608 3528
rect 255924 3488 256608 3516
rect 255924 3476 255930 3488
rect 256602 3476 256608 3488
rect 256660 3476 256666 3528
rect 257062 3476 257068 3528
rect 257120 3516 257126 3528
rect 257982 3516 257988 3528
rect 257120 3488 257988 3516
rect 257120 3476 257126 3488
rect 257982 3476 257988 3488
rect 258040 3476 258046 3528
rect 258258 3476 258264 3528
rect 258316 3516 258322 3528
rect 259362 3516 259368 3528
rect 258316 3488 259368 3516
rect 258316 3476 258322 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 259454 3476 259460 3528
rect 259512 3516 259518 3528
rect 260742 3516 260748 3528
rect 259512 3488 260748 3516
rect 259512 3476 259518 3488
rect 260742 3476 260748 3488
rect 260800 3476 260806 3528
rect 262950 3476 262956 3528
rect 263008 3516 263014 3528
rect 263502 3516 263508 3528
rect 263008 3488 263508 3516
rect 263008 3476 263014 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 264882 3516 264888 3528
rect 264204 3488 264888 3516
rect 264204 3476 264210 3488
rect 264882 3476 264888 3488
rect 264940 3476 264946 3528
rect 266538 3476 266544 3528
rect 266596 3516 266602 3528
rect 267642 3516 267648 3528
rect 266596 3488 267648 3516
rect 266596 3476 266602 3488
rect 267642 3476 267648 3488
rect 267700 3476 267706 3528
rect 272426 3476 272432 3528
rect 272484 3516 272490 3528
rect 273162 3516 273168 3528
rect 272484 3488 273168 3516
rect 272484 3476 272490 3488
rect 273162 3476 273168 3488
rect 273220 3476 273226 3528
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 274542 3516 274548 3528
rect 273680 3488 274548 3516
rect 273680 3476 273686 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 274818 3476 274824 3528
rect 274876 3516 274882 3528
rect 275922 3516 275928 3528
rect 274876 3488 275928 3516
rect 274876 3476 274882 3488
rect 275922 3476 275928 3488
rect 275980 3476 275986 3528
rect 280706 3476 280712 3528
rect 280764 3516 280770 3528
rect 281442 3516 281448 3528
rect 280764 3488 281448 3516
rect 280764 3476 280770 3488
rect 281442 3476 281448 3488
rect 281500 3476 281506 3528
rect 281902 3476 281908 3528
rect 281960 3516 281966 3528
rect 282822 3516 282828 3528
rect 281960 3488 282828 3516
rect 281960 3476 281966 3488
rect 282822 3476 282828 3488
rect 282880 3476 282886 3528
rect 287790 3476 287796 3528
rect 287848 3516 287854 3528
rect 288342 3516 288348 3528
rect 287848 3488 288348 3516
rect 287848 3476 287854 3488
rect 288342 3476 288348 3488
rect 288400 3476 288406 3528
rect 288986 3476 288992 3528
rect 289044 3516 289050 3528
rect 289722 3516 289728 3528
rect 289044 3488 289728 3516
rect 289044 3476 289050 3488
rect 289722 3476 289728 3488
rect 289780 3476 289786 3528
rect 290182 3476 290188 3528
rect 290240 3516 290246 3528
rect 291286 3516 291292 3528
rect 290240 3488 291292 3516
rect 290240 3476 290246 3488
rect 291286 3476 291292 3488
rect 291344 3476 291350 3528
rect 291378 3476 291384 3528
rect 291436 3516 291442 3528
rect 292482 3516 292488 3528
rect 291436 3488 292488 3516
rect 291436 3476 291442 3488
rect 292482 3476 292488 3488
rect 292540 3476 292546 3528
rect 293678 3476 293684 3528
rect 293736 3516 293742 3528
rect 294230 3516 294236 3528
rect 293736 3488 294236 3516
rect 293736 3476 293742 3488
rect 294230 3476 294236 3488
rect 294288 3476 294294 3528
rect 296070 3476 296076 3528
rect 296128 3516 296134 3528
rect 296622 3516 296628 3528
rect 296128 3488 296628 3516
rect 296128 3476 296134 3488
rect 296622 3476 296628 3488
rect 296680 3476 296686 3528
rect 300946 3476 300952 3528
rect 301004 3516 301010 3528
rect 301958 3516 301964 3528
rect 301004 3488 301964 3516
rect 301004 3476 301010 3488
rect 301958 3476 301964 3488
rect 302016 3476 302022 3528
rect 302234 3476 302240 3528
rect 302292 3516 302298 3528
rect 303154 3516 303160 3528
rect 302292 3488 303160 3516
rect 302292 3476 302298 3488
rect 303154 3476 303160 3488
rect 303212 3476 303218 3528
rect 309134 3476 309140 3528
rect 309192 3516 309198 3528
rect 310238 3516 310244 3528
rect 309192 3488 310244 3516
rect 309192 3476 309198 3488
rect 310238 3476 310244 3488
rect 310296 3476 310302 3528
rect 310422 3476 310428 3528
rect 310480 3516 310486 3528
rect 311434 3516 311440 3528
rect 310480 3488 311440 3516
rect 310480 3476 310486 3488
rect 311434 3476 311440 3488
rect 311492 3476 311498 3528
rect 311802 3476 311808 3528
rect 311860 3516 311866 3528
rect 312630 3516 312636 3528
rect 311860 3488 312636 3516
rect 311860 3476 311866 3488
rect 312630 3476 312636 3488
rect 312688 3476 312694 3528
rect 314562 3476 314568 3528
rect 314620 3516 314626 3528
rect 315022 3516 315028 3528
rect 314620 3488 315028 3516
rect 314620 3476 314626 3488
rect 315022 3476 315028 3488
rect 315080 3476 315086 3528
rect 317322 3476 317328 3528
rect 317380 3516 317386 3528
rect 318518 3516 318524 3528
rect 317380 3488 318524 3516
rect 317380 3476 317386 3488
rect 318518 3476 318524 3488
rect 318576 3476 318582 3528
rect 318702 3476 318708 3528
rect 318760 3516 318766 3528
rect 319714 3516 319720 3528
rect 318760 3488 319720 3516
rect 318760 3476 318766 3488
rect 319714 3476 319720 3488
rect 319772 3476 319778 3528
rect 329742 3476 329748 3528
rect 329800 3516 329806 3528
rect 332686 3516 332692 3528
rect 329800 3488 332692 3516
rect 329800 3476 329806 3488
rect 332686 3476 332692 3488
rect 332744 3476 332750 3528
rect 335998 3476 336004 3528
rect 336056 3516 336062 3528
rect 337470 3516 337476 3528
rect 336056 3488 337476 3516
rect 336056 3476 336062 3488
rect 337470 3476 337476 3488
rect 337528 3476 337534 3528
rect 342070 3476 342076 3528
rect 342128 3516 342134 3528
rect 348050 3516 348056 3528
rect 342128 3488 348056 3516
rect 342128 3476 342134 3488
rect 348050 3476 348056 3488
rect 348108 3476 348114 3528
rect 350442 3476 350448 3528
rect 350500 3516 350506 3528
rect 357526 3516 357532 3528
rect 350500 3488 357532 3516
rect 350500 3476 350506 3488
rect 357526 3476 357532 3488
rect 357584 3476 357590 3528
rect 360010 3476 360016 3528
rect 360068 3516 360074 3528
rect 369394 3516 369400 3528
rect 360068 3488 369400 3516
rect 360068 3476 360074 3488
rect 369394 3476 369400 3488
rect 369452 3476 369458 3528
rect 372430 3476 372436 3528
rect 372488 3516 372494 3528
rect 383562 3516 383568 3528
rect 372488 3488 383568 3516
rect 372488 3476 372494 3488
rect 383562 3476 383568 3488
rect 383620 3476 383626 3528
rect 384942 3476 384948 3528
rect 385000 3516 385006 3528
rect 397730 3516 397736 3528
rect 385000 3488 397736 3516
rect 385000 3476 385006 3488
rect 397730 3476 397736 3488
rect 397788 3476 397794 3528
rect 400030 3476 400036 3528
rect 400088 3516 400094 3528
rect 415486 3516 415492 3528
rect 400088 3488 415492 3516
rect 400088 3476 400094 3488
rect 415486 3476 415492 3488
rect 415544 3476 415550 3528
rect 422110 3476 422116 3528
rect 422168 3516 422174 3528
rect 441522 3516 441528 3528
rect 422168 3488 441528 3516
rect 422168 3476 422174 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 445570 3476 445576 3528
rect 445628 3516 445634 3528
rect 468662 3516 468668 3528
rect 445628 3488 468668 3516
rect 445628 3476 445634 3488
rect 468662 3476 468668 3488
rect 468720 3476 468726 3528
rect 470502 3476 470508 3528
rect 470560 3516 470566 3528
rect 497090 3516 497096 3528
rect 470560 3488 497096 3516
rect 470560 3476 470566 3488
rect 497090 3476 497096 3488
rect 497148 3476 497154 3528
rect 498102 3476 498108 3528
rect 498160 3516 498166 3528
rect 529014 3516 529020 3528
rect 498160 3488 529020 3516
rect 498160 3476 498166 3488
rect 529014 3476 529020 3488
rect 529072 3476 529078 3528
rect 531130 3476 531136 3528
rect 531188 3516 531194 3528
rect 568022 3516 568028 3528
rect 531188 3488 568028 3516
rect 531188 3476 531194 3488
rect 568022 3476 568028 3488
rect 568080 3476 568086 3528
rect 76248 3352 78720 3380
rect 78784 3420 85620 3448
rect 76248 3340 76254 3352
rect 78784 3312 78812 3420
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 83274 3340 83280 3392
rect 83332 3380 83338 3392
rect 84102 3380 84108 3392
rect 83332 3352 84108 3380
rect 83332 3340 83338 3352
rect 84102 3340 84108 3352
rect 84160 3340 84166 3392
rect 64846 3284 78812 3312
rect 85592 3312 85620 3420
rect 85666 3408 85672 3460
rect 85724 3448 85730 3460
rect 88978 3448 88984 3460
rect 85724 3420 88984 3448
rect 85724 3408 85730 3420
rect 88978 3408 88984 3420
rect 89036 3408 89042 3460
rect 90358 3408 90364 3460
rect 90416 3448 90422 3460
rect 91002 3448 91008 3460
rect 90416 3420 91008 3448
rect 90416 3408 90422 3420
rect 91002 3408 91008 3420
rect 91060 3408 91066 3460
rect 91554 3408 91560 3460
rect 91612 3448 91618 3460
rect 92382 3448 92388 3460
rect 91612 3420 92388 3448
rect 91612 3408 91618 3420
rect 92382 3408 92388 3420
rect 92440 3408 92446 3460
rect 97442 3408 97448 3460
rect 97500 3448 97506 3460
rect 97902 3448 97908 3460
rect 97500 3420 97908 3448
rect 97500 3408 97506 3420
rect 97902 3408 97908 3420
rect 97960 3408 97966 3460
rect 98638 3408 98644 3460
rect 98696 3448 98702 3460
rect 99282 3448 99288 3460
rect 98696 3420 99288 3448
rect 98696 3408 98702 3420
rect 99282 3408 99288 3420
rect 99340 3408 99346 3460
rect 99834 3408 99840 3460
rect 99892 3448 99898 3460
rect 100662 3448 100668 3460
rect 99892 3420 100668 3448
rect 99892 3408 99898 3420
rect 100662 3408 100668 3420
rect 100720 3408 100726 3460
rect 101030 3408 101036 3460
rect 101088 3448 101094 3460
rect 102042 3448 102048 3460
rect 101088 3420 102048 3448
rect 101088 3408 101094 3420
rect 102042 3408 102048 3420
rect 102100 3408 102106 3460
rect 122926 3448 122932 3460
rect 103486 3420 122932 3448
rect 89162 3340 89168 3392
rect 89220 3380 89226 3392
rect 91738 3380 91744 3392
rect 89220 3352 91744 3380
rect 89220 3340 89226 3352
rect 91738 3340 91744 3352
rect 91796 3340 91802 3392
rect 93946 3340 93952 3392
rect 94004 3380 94010 3392
rect 103486 3380 103514 3420
rect 122926 3408 122932 3420
rect 122984 3408 122990 3460
rect 161290 3408 161296 3460
rect 161348 3448 161354 3460
rect 180058 3448 180064 3460
rect 161348 3420 180064 3448
rect 161348 3408 161354 3420
rect 180058 3408 180064 3420
rect 180116 3408 180122 3460
rect 189718 3408 189724 3460
rect 189776 3448 189782 3460
rect 190362 3448 190368 3460
rect 189776 3420 190368 3448
rect 189776 3408 189782 3420
rect 190362 3408 190368 3420
rect 190420 3408 190426 3460
rect 265342 3408 265348 3460
rect 265400 3448 265406 3460
rect 266998 3448 267004 3460
rect 265400 3420 267004 3448
rect 265400 3408 265406 3420
rect 266998 3408 267004 3420
rect 267056 3408 267062 3460
rect 325602 3408 325608 3460
rect 325660 3448 325666 3460
rect 329190 3448 329196 3460
rect 325660 3420 329196 3448
rect 325660 3408 325666 3420
rect 329190 3408 329196 3420
rect 329248 3408 329254 3460
rect 331122 3408 331128 3460
rect 331180 3448 331186 3460
rect 335078 3448 335084 3460
rect 331180 3420 335084 3448
rect 331180 3408 331186 3420
rect 335078 3408 335084 3420
rect 335136 3408 335142 3460
rect 335262 3408 335268 3460
rect 335320 3448 335326 3460
rect 339862 3448 339868 3460
rect 335320 3420 339868 3448
rect 335320 3408 335326 3420
rect 339862 3408 339868 3420
rect 339920 3408 339926 3460
rect 353110 3408 353116 3460
rect 353168 3448 353174 3460
rect 361114 3448 361120 3460
rect 353168 3420 361120 3448
rect 353168 3408 353174 3420
rect 361114 3408 361120 3420
rect 361172 3408 361178 3460
rect 364150 3408 364156 3460
rect 364208 3448 364214 3460
rect 374086 3448 374092 3460
rect 364208 3420 374092 3448
rect 364208 3408 364214 3420
rect 374086 3408 374092 3420
rect 374144 3408 374150 3460
rect 378042 3408 378048 3460
rect 378100 3448 378106 3460
rect 389450 3448 389456 3460
rect 378100 3420 389456 3448
rect 378100 3408 378106 3420
rect 389450 3408 389456 3420
rect 389508 3408 389514 3460
rect 391842 3408 391848 3460
rect 391900 3448 391906 3460
rect 406010 3448 406016 3460
rect 391900 3420 406016 3448
rect 391900 3408 391906 3420
rect 406010 3408 406016 3420
rect 406068 3408 406074 3460
rect 406930 3408 406936 3460
rect 406988 3448 406994 3460
rect 423766 3448 423772 3460
rect 406988 3420 423772 3448
rect 406988 3408 406994 3420
rect 423766 3408 423772 3420
rect 423824 3408 423830 3460
rect 426342 3408 426348 3460
rect 426400 3448 426406 3460
rect 446214 3448 446220 3460
rect 426400 3420 446220 3448
rect 426400 3408 426406 3420
rect 446214 3408 446220 3420
rect 446272 3408 446278 3460
rect 449710 3408 449716 3460
rect 449768 3448 449774 3460
rect 473446 3448 473452 3460
rect 449768 3420 473452 3448
rect 449768 3408 449774 3420
rect 473446 3408 473452 3420
rect 473504 3408 473510 3460
rect 477402 3408 477408 3460
rect 477460 3448 477466 3460
rect 504174 3448 504180 3460
rect 477460 3420 504180 3448
rect 477460 3408 477466 3420
rect 504174 3408 504180 3420
rect 504232 3408 504238 3460
rect 506382 3408 506388 3460
rect 506440 3448 506446 3460
rect 538398 3448 538404 3460
rect 506440 3420 538404 3448
rect 506440 3408 506446 3420
rect 538398 3408 538404 3420
rect 538456 3408 538462 3460
rect 540330 3408 540336 3460
rect 540388 3448 540394 3460
rect 543182 3448 543188 3460
rect 540388 3420 543188 3448
rect 540388 3408 540394 3420
rect 543182 3408 543188 3420
rect 543240 3408 543246 3460
rect 544470 3408 544476 3460
rect 544528 3448 544534 3460
rect 546678 3448 546684 3460
rect 544528 3420 546684 3448
rect 544528 3408 544534 3420
rect 546678 3408 546684 3420
rect 546736 3408 546742 3460
rect 546773 3451 546831 3457
rect 546773 3417 546785 3451
rect 546819 3448 546831 3451
rect 577406 3448 577412 3460
rect 546819 3420 577412 3448
rect 546819 3417 546831 3420
rect 546773 3411 546831 3417
rect 577406 3408 577412 3420
rect 577464 3408 577470 3460
rect 94004 3352 103514 3380
rect 94004 3340 94010 3352
rect 114002 3340 114008 3392
rect 114060 3380 114066 3392
rect 114462 3380 114468 3392
rect 114060 3352 114468 3380
rect 114060 3340 114066 3352
rect 114462 3340 114468 3352
rect 114520 3340 114526 3392
rect 115198 3340 115204 3392
rect 115256 3380 115262 3392
rect 115842 3380 115848 3392
rect 115256 3352 115848 3380
rect 115256 3340 115262 3352
rect 115842 3340 115848 3352
rect 115900 3340 115906 3392
rect 116394 3340 116400 3392
rect 116452 3380 116458 3392
rect 117222 3380 117228 3392
rect 116452 3352 117228 3380
rect 116452 3340 116458 3352
rect 117222 3340 117228 3352
rect 117280 3340 117286 3392
rect 117590 3340 117596 3392
rect 117648 3380 117654 3392
rect 118602 3380 118608 3392
rect 117648 3352 118608 3380
rect 117648 3340 117654 3352
rect 118602 3340 118608 3352
rect 118660 3340 118666 3392
rect 118786 3340 118792 3392
rect 118844 3380 118850 3392
rect 119798 3380 119804 3392
rect 118844 3352 119804 3380
rect 118844 3340 118850 3352
rect 119798 3340 119804 3352
rect 119856 3340 119862 3392
rect 122282 3340 122288 3392
rect 122340 3380 122346 3392
rect 122742 3380 122748 3392
rect 122340 3352 122748 3380
rect 122340 3340 122346 3352
rect 122742 3340 122748 3352
rect 122800 3340 122806 3392
rect 329650 3340 329656 3392
rect 329708 3380 329714 3392
rect 333882 3380 333888 3392
rect 329708 3352 333888 3380
rect 329708 3340 329714 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 339402 3340 339408 3392
rect 339460 3380 339466 3392
rect 344554 3380 344560 3392
rect 339460 3352 344560 3380
rect 339460 3340 339466 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 347682 3340 347688 3392
rect 347740 3380 347746 3392
rect 354030 3380 354036 3392
rect 347740 3352 354036 3380
rect 347740 3340 347746 3352
rect 354030 3340 354036 3352
rect 354088 3340 354094 3392
rect 371142 3340 371148 3392
rect 371200 3380 371206 3392
rect 381170 3380 381176 3392
rect 371200 3352 381176 3380
rect 371200 3340 371206 3352
rect 381170 3340 381176 3352
rect 381228 3340 381234 3392
rect 387702 3340 387708 3392
rect 387760 3380 387766 3392
rect 400122 3380 400128 3392
rect 387760 3352 400128 3380
rect 387760 3340 387766 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 400214 3340 400220 3392
rect 400272 3380 400278 3392
rect 414290 3380 414296 3392
rect 400272 3352 414296 3380
rect 400272 3340 400278 3352
rect 414290 3340 414296 3352
rect 414348 3340 414354 3392
rect 415302 3340 415308 3392
rect 415360 3380 415366 3392
rect 432046 3380 432052 3392
rect 415360 3352 432052 3380
rect 415360 3340 415366 3352
rect 432046 3340 432052 3352
rect 432104 3340 432110 3392
rect 437382 3340 437388 3392
rect 437440 3380 437446 3392
rect 457990 3380 457996 3392
rect 437440 3352 457996 3380
rect 437440 3340 437446 3352
rect 457990 3340 457996 3352
rect 458048 3340 458054 3392
rect 458082 3340 458088 3392
rect 458140 3380 458146 3392
rect 482830 3380 482836 3392
rect 458140 3352 482836 3380
rect 458140 3340 458146 3352
rect 482830 3340 482836 3352
rect 482888 3340 482894 3392
rect 482922 3340 482928 3392
rect 482980 3380 482986 3392
rect 511258 3380 511264 3392
rect 482980 3352 511264 3380
rect 482980 3340 482986 3352
rect 511258 3340 511264 3352
rect 511316 3340 511322 3392
rect 511902 3340 511908 3392
rect 511960 3380 511966 3392
rect 545482 3380 545488 3392
rect 511960 3352 545488 3380
rect 511960 3340 511966 3352
rect 545482 3340 545488 3352
rect 545540 3340 545546 3392
rect 547230 3340 547236 3392
rect 547288 3380 547294 3392
rect 550266 3380 550272 3392
rect 547288 3352 550272 3380
rect 547288 3340 547294 3352
rect 550266 3340 550272 3352
rect 550324 3340 550330 3392
rect 552661 3383 552719 3389
rect 552661 3349 552673 3383
rect 552707 3380 552719 3383
rect 578602 3380 578608 3392
rect 552707 3352 578608 3380
rect 552707 3349 552719 3352
rect 552661 3343 552719 3349
rect 578602 3340 578608 3352
rect 578660 3340 578666 3392
rect 93118 3312 93124 3324
rect 85592 3284 93124 3312
rect 93118 3272 93124 3284
rect 93176 3272 93182 3324
rect 196802 3272 196808 3324
rect 196860 3312 196866 3324
rect 197262 3312 197268 3324
rect 196860 3284 197268 3312
rect 196860 3272 196866 3284
rect 197262 3272 197268 3284
rect 197320 3272 197326 3324
rect 221550 3272 221556 3324
rect 221608 3312 221614 3324
rect 222102 3312 222108 3324
rect 221608 3284 222108 3312
rect 221608 3272 221614 3284
rect 222102 3272 222108 3284
rect 222160 3272 222166 3324
rect 271230 3272 271236 3324
rect 271288 3312 271294 3324
rect 271782 3312 271788 3324
rect 271288 3284 271788 3312
rect 271288 3272 271294 3284
rect 271782 3272 271788 3284
rect 271840 3272 271846 3324
rect 276014 3272 276020 3324
rect 276072 3312 276078 3324
rect 277302 3312 277308 3324
rect 276072 3284 277308 3312
rect 276072 3272 276078 3284
rect 277302 3272 277308 3284
rect 277360 3272 277366 3324
rect 279510 3272 279516 3324
rect 279568 3312 279574 3324
rect 280062 3312 280068 3324
rect 279568 3284 280068 3312
rect 279568 3272 279574 3284
rect 280062 3272 280068 3284
rect 280120 3272 280126 3324
rect 304994 3272 305000 3324
rect 305052 3312 305058 3324
rect 305546 3312 305552 3324
rect 305052 3284 305552 3312
rect 305052 3272 305058 3284
rect 305546 3272 305552 3284
rect 305604 3272 305610 3324
rect 325510 3272 325516 3324
rect 325568 3312 325574 3324
rect 327994 3312 328000 3324
rect 325568 3284 328000 3312
rect 325568 3272 325574 3284
rect 327994 3272 328000 3284
rect 328052 3272 328058 3324
rect 338022 3272 338028 3324
rect 338080 3312 338086 3324
rect 343358 3312 343364 3324
rect 338080 3284 343364 3312
rect 338080 3272 338086 3284
rect 343358 3272 343364 3284
rect 343416 3272 343422 3324
rect 375190 3272 375196 3324
rect 375248 3312 375254 3324
rect 385954 3312 385960 3324
rect 375248 3284 385960 3312
rect 375248 3272 375254 3284
rect 385954 3272 385960 3284
rect 386012 3272 386018 3324
rect 389082 3272 389088 3324
rect 389140 3312 389146 3324
rect 402514 3312 402520 3324
rect 389140 3284 402520 3312
rect 389140 3272 389146 3284
rect 402514 3272 402520 3284
rect 402572 3272 402578 3324
rect 402882 3272 402888 3324
rect 402940 3312 402946 3324
rect 417878 3312 417884 3324
rect 402940 3284 417884 3312
rect 402940 3272 402946 3284
rect 417878 3272 417884 3284
rect 417936 3272 417942 3324
rect 418062 3272 418068 3324
rect 418120 3312 418126 3324
rect 435542 3312 435548 3324
rect 418120 3284 435548 3312
rect 418120 3272 418126 3284
rect 435542 3272 435548 3284
rect 435600 3272 435606 3324
rect 440142 3272 440148 3324
rect 440200 3312 440206 3324
rect 461578 3312 461584 3324
rect 440200 3284 461584 3312
rect 440200 3272 440206 3284
rect 461578 3272 461584 3284
rect 461636 3272 461642 3324
rect 462222 3272 462228 3324
rect 462280 3312 462286 3324
rect 486418 3312 486424 3324
rect 462280 3284 486424 3312
rect 462280 3272 462286 3284
rect 486418 3272 486424 3284
rect 486476 3272 486482 3324
rect 488442 3272 488448 3324
rect 488500 3312 488506 3324
rect 517146 3312 517152 3324
rect 488500 3284 517152 3312
rect 488500 3272 488506 3284
rect 517146 3272 517152 3284
rect 517204 3272 517210 3324
rect 520182 3272 520188 3324
rect 520240 3312 520246 3324
rect 553762 3312 553768 3324
rect 520240 3284 553768 3312
rect 520240 3272 520246 3284
rect 553762 3272 553768 3284
rect 553820 3272 553826 3324
rect 28902 3204 28908 3256
rect 28960 3244 28966 3256
rect 32306 3244 32312 3256
rect 28960 3216 32312 3244
rect 28960 3204 28966 3216
rect 32306 3204 32312 3216
rect 32364 3204 32370 3256
rect 183738 3204 183744 3256
rect 183796 3244 183802 3256
rect 184842 3244 184848 3256
rect 183796 3216 184848 3244
rect 183796 3204 183802 3216
rect 184842 3204 184848 3216
rect 184900 3204 184906 3256
rect 200298 3204 200304 3256
rect 200356 3244 200362 3256
rect 201402 3244 201408 3256
rect 200356 3216 201408 3244
rect 200356 3204 200362 3216
rect 201402 3204 201408 3216
rect 201460 3204 201466 3256
rect 225138 3204 225144 3256
rect 225196 3244 225202 3256
rect 226242 3244 226248 3256
rect 225196 3216 226248 3244
rect 225196 3204 225202 3216
rect 226242 3204 226248 3216
rect 226300 3204 226306 3256
rect 322842 3204 322848 3256
rect 322900 3244 322906 3256
rect 325602 3244 325608 3256
rect 322900 3216 325608 3244
rect 322900 3204 322906 3216
rect 325602 3204 325608 3216
rect 325660 3204 325666 3256
rect 338758 3204 338764 3256
rect 338816 3244 338822 3256
rect 342162 3244 342168 3256
rect 338816 3216 342168 3244
rect 338816 3204 338822 3216
rect 342162 3204 342168 3216
rect 342220 3204 342226 3256
rect 390462 3204 390468 3256
rect 390520 3244 390526 3256
rect 403618 3244 403624 3256
rect 390520 3216 403624 3244
rect 390520 3204 390526 3216
rect 403618 3204 403624 3216
rect 403676 3204 403682 3256
rect 412542 3204 412548 3256
rect 412600 3244 412606 3256
rect 429654 3244 429660 3256
rect 412600 3216 429660 3244
rect 412600 3204 412606 3216
rect 429654 3204 429660 3216
rect 429712 3204 429718 3256
rect 430482 3204 430488 3256
rect 430540 3244 430546 3256
rect 449802 3244 449808 3256
rect 430540 3216 449808 3244
rect 430540 3204 430546 3216
rect 449802 3204 449808 3216
rect 449860 3204 449866 3256
rect 453850 3204 453856 3256
rect 453908 3244 453914 3256
rect 476942 3244 476948 3256
rect 453908 3216 476948 3244
rect 453908 3204 453914 3216
rect 476942 3204 476948 3216
rect 477000 3204 477006 3256
rect 478782 3204 478788 3256
rect 478840 3244 478846 3256
rect 506474 3244 506480 3256
rect 478840 3216 506480 3244
rect 478840 3204 478846 3216
rect 506474 3204 506480 3216
rect 506532 3204 506538 3256
rect 512638 3204 512644 3256
rect 512696 3244 512702 3256
rect 521838 3244 521844 3256
rect 512696 3216 521844 3244
rect 512696 3204 512702 3216
rect 521838 3204 521844 3216
rect 521896 3204 521902 3256
rect 522942 3204 522948 3256
rect 523000 3244 523006 3256
rect 523000 3216 552612 3244
rect 523000 3204 523006 3216
rect 78582 3136 78588 3188
rect 78640 3176 78646 3188
rect 81986 3176 81992 3188
rect 78640 3148 81992 3176
rect 78640 3136 78646 3148
rect 81986 3136 81992 3148
rect 82044 3136 82050 3188
rect 241698 3136 241704 3188
rect 241756 3176 241762 3188
rect 242802 3176 242808 3188
rect 241756 3148 242808 3176
rect 241756 3136 241762 3148
rect 242802 3136 242808 3148
rect 242860 3136 242866 3188
rect 321370 3136 321376 3188
rect 321428 3176 321434 3188
rect 324406 3176 324412 3188
rect 321428 3148 324412 3176
rect 321428 3136 321434 3148
rect 324406 3136 324412 3148
rect 324464 3136 324470 3188
rect 326982 3136 326988 3188
rect 327040 3176 327046 3188
rect 330386 3176 330392 3188
rect 327040 3148 330392 3176
rect 327040 3136 327046 3148
rect 330386 3136 330392 3148
rect 330444 3136 330450 3188
rect 332502 3136 332508 3188
rect 332560 3176 332566 3188
rect 336274 3176 336280 3188
rect 332560 3148 336280 3176
rect 332560 3136 332566 3148
rect 336274 3136 336280 3148
rect 336332 3136 336338 3188
rect 407022 3136 407028 3188
rect 407080 3176 407086 3188
rect 422570 3176 422576 3188
rect 407080 3148 422576 3176
rect 407080 3136 407086 3148
rect 422570 3136 422576 3148
rect 422628 3136 422634 3188
rect 424962 3136 424968 3188
rect 425020 3176 425026 3188
rect 443822 3176 443828 3188
rect 425020 3148 443828 3176
rect 425020 3136 425026 3148
rect 443822 3136 443828 3148
rect 443880 3136 443886 3188
rect 451182 3136 451188 3188
rect 451240 3176 451246 3188
rect 474550 3176 474556 3188
rect 451240 3148 474556 3176
rect 451240 3136 451246 3148
rect 474550 3136 474556 3148
rect 474608 3136 474614 3188
rect 476022 3136 476028 3188
rect 476080 3176 476086 3188
rect 502978 3176 502984 3188
rect 476080 3148 502984 3176
rect 476080 3136 476086 3148
rect 502978 3136 502984 3148
rect 503036 3136 503042 3188
rect 507762 3136 507768 3188
rect 507820 3176 507826 3188
rect 539594 3176 539600 3188
rect 507820 3148 539600 3176
rect 507820 3136 507826 3148
rect 539594 3136 539600 3148
rect 539652 3136 539658 3188
rect 548518 3136 548524 3188
rect 548576 3176 548582 3188
rect 552584 3176 552612 3216
rect 557350 3176 557356 3188
rect 548576 3148 549208 3176
rect 552584 3148 557356 3176
rect 548576 3136 548582 3148
rect 102226 3068 102232 3120
rect 102284 3108 102290 3120
rect 103422 3108 103428 3120
rect 102284 3080 103428 3108
rect 102284 3068 102290 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 126974 3068 126980 3120
rect 127032 3108 127038 3120
rect 129458 3108 129464 3120
rect 127032 3080 129464 3108
rect 127032 3068 127038 3080
rect 129458 3068 129464 3080
rect 129516 3068 129522 3120
rect 246390 3068 246396 3120
rect 246448 3108 246454 3120
rect 246942 3108 246948 3120
rect 246448 3080 246948 3108
rect 246448 3068 246454 3080
rect 246942 3068 246948 3080
rect 247000 3068 247006 3120
rect 349062 3068 349068 3120
rect 349120 3108 349126 3120
rect 356330 3108 356336 3120
rect 349120 3080 356336 3108
rect 349120 3068 349126 3080
rect 356330 3068 356336 3080
rect 356388 3068 356394 3120
rect 394602 3068 394608 3120
rect 394660 3108 394666 3120
rect 408402 3108 408408 3120
rect 394660 3080 408408 3108
rect 394660 3068 394666 3080
rect 408402 3068 408408 3080
rect 408460 3068 408466 3120
rect 423582 3068 423588 3120
rect 423640 3108 423646 3120
rect 442626 3108 442632 3120
rect 423640 3080 442632 3108
rect 423640 3068 423646 3080
rect 442626 3068 442632 3080
rect 442684 3068 442690 3120
rect 449710 3068 449716 3120
rect 449768 3108 449774 3120
rect 472250 3108 472256 3120
rect 449768 3080 472256 3108
rect 449768 3068 449774 3080
rect 472250 3068 472256 3080
rect 472308 3068 472314 3120
rect 480162 3068 480168 3120
rect 480220 3108 480226 3120
rect 507670 3108 507676 3120
rect 480220 3080 507676 3108
rect 480220 3068 480226 3080
rect 507670 3068 507676 3080
rect 507728 3068 507734 3120
rect 516042 3068 516048 3120
rect 516100 3108 516106 3120
rect 549070 3108 549076 3120
rect 516100 3080 549076 3108
rect 516100 3068 516106 3080
rect 549070 3068 549076 3080
rect 549128 3068 549134 3120
rect 549180 3108 549208 3148
rect 557350 3136 557356 3148
rect 557408 3136 557414 3188
rect 580994 3176 581000 3188
rect 557506 3148 581000 3176
rect 557506 3108 557534 3148
rect 580994 3136 581000 3148
rect 581052 3136 581058 3188
rect 549180 3080 557534 3108
rect 25314 3000 25320 3052
rect 25372 3040 25378 3052
rect 26142 3040 26148 3052
rect 25372 3012 26148 3040
rect 25372 3000 25378 3012
rect 26142 3000 26148 3012
rect 26200 3000 26206 3052
rect 143534 3000 143540 3052
rect 143592 3040 143598 3052
rect 144638 3040 144644 3052
rect 143592 3012 144644 3040
rect 143592 3000 143598 3012
rect 144638 3000 144644 3012
rect 144696 3000 144702 3052
rect 164878 3000 164884 3052
rect 164936 3040 164942 3052
rect 165522 3040 165528 3052
rect 164936 3012 165528 3040
rect 164936 3000 164942 3012
rect 165522 3000 165528 3012
rect 165580 3000 165586 3052
rect 208578 3000 208584 3052
rect 208636 3040 208642 3052
rect 209682 3040 209688 3052
rect 208636 3012 209688 3040
rect 208636 3000 208642 3012
rect 209682 3000 209688 3012
rect 209740 3000 209746 3052
rect 248782 3000 248788 3052
rect 248840 3040 248846 3052
rect 249702 3040 249708 3052
rect 248840 3012 249708 3040
rect 248840 3000 248846 3012
rect 249702 3000 249708 3012
rect 249760 3000 249766 3052
rect 283098 3000 283104 3052
rect 283156 3040 283162 3052
rect 284938 3040 284944 3052
rect 283156 3012 284944 3040
rect 283156 3000 283162 3012
rect 284938 3000 284944 3012
rect 284996 3000 285002 3052
rect 318610 3000 318616 3052
rect 318668 3040 318674 3052
rect 320910 3040 320916 3052
rect 318668 3012 320916 3040
rect 318668 3000 318674 3012
rect 320910 3000 320916 3012
rect 320968 3000 320974 3052
rect 340782 3000 340788 3052
rect 340840 3040 340846 3052
rect 345750 3040 345756 3052
rect 340840 3012 345756 3040
rect 340840 3000 340846 3012
rect 345750 3000 345756 3012
rect 345808 3000 345814 3052
rect 346302 3000 346308 3052
rect 346360 3040 346366 3052
rect 352834 3040 352840 3052
rect 346360 3012 352840 3040
rect 346360 3000 346366 3012
rect 352834 3000 352840 3012
rect 352892 3000 352898 3052
rect 355962 3000 355968 3052
rect 356020 3040 356026 3052
rect 363506 3040 363512 3052
rect 356020 3012 363512 3040
rect 356020 3000 356026 3012
rect 363506 3000 363512 3012
rect 363564 3000 363570 3052
rect 416590 3000 416596 3052
rect 416648 3040 416654 3052
rect 434438 3040 434444 3052
rect 416648 3012 434444 3040
rect 416648 3000 416654 3012
rect 434438 3000 434444 3012
rect 434496 3000 434502 3052
rect 444282 3000 444288 3052
rect 444340 3040 444346 3052
rect 466270 3040 466276 3052
rect 444340 3012 466276 3040
rect 444340 3000 444346 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 466362 3000 466368 3052
rect 466420 3040 466426 3052
rect 492306 3040 492312 3052
rect 466420 3012 492312 3040
rect 466420 3000 466426 3012
rect 492306 3000 492312 3012
rect 492364 3000 492370 3052
rect 509142 3000 509148 3052
rect 509200 3040 509206 3052
rect 541986 3040 541992 3052
rect 509200 3012 541992 3040
rect 509200 3000 509206 3012
rect 541986 3000 541992 3012
rect 542044 3000 542050 3052
rect 546773 3043 546831 3049
rect 546773 3040 546785 3043
rect 542096 3012 546785 3040
rect 284294 2932 284300 2984
rect 284352 2972 284358 2984
rect 285858 2972 285864 2984
rect 284352 2944 285864 2972
rect 284352 2932 284358 2944
rect 285858 2932 285864 2944
rect 285916 2932 285922 2984
rect 314470 2932 314476 2984
rect 314528 2972 314534 2984
rect 316218 2972 316224 2984
rect 314528 2944 316224 2972
rect 314528 2932 314534 2944
rect 316218 2932 316224 2944
rect 316276 2932 316282 2984
rect 321462 2932 321468 2984
rect 321520 2972 321526 2984
rect 323302 2972 323308 2984
rect 321520 2944 323308 2972
rect 321520 2932 321526 2944
rect 323302 2932 323308 2944
rect 323360 2932 323366 2984
rect 409782 2932 409788 2984
rect 409840 2972 409846 2984
rect 426158 2972 426164 2984
rect 409840 2944 426164 2972
rect 409840 2932 409846 2944
rect 426158 2932 426164 2944
rect 426216 2932 426222 2984
rect 434622 2932 434628 2984
rect 434680 2972 434686 2984
rect 454494 2972 454500 2984
rect 434680 2944 454500 2972
rect 434680 2932 434686 2944
rect 454494 2932 454500 2944
rect 454552 2932 454558 2984
rect 460842 2932 460848 2984
rect 460900 2972 460906 2984
rect 485222 2972 485228 2984
rect 460900 2944 485228 2972
rect 460900 2932 460906 2944
rect 485222 2932 485228 2944
rect 485280 2932 485286 2984
rect 503622 2932 503628 2984
rect 503680 2972 503686 2984
rect 534902 2972 534908 2984
rect 503680 2944 534908 2972
rect 503680 2932 503686 2944
rect 534902 2932 534908 2944
rect 534960 2932 534966 2984
rect 539502 2932 539508 2984
rect 539560 2972 539566 2984
rect 542096 2972 542124 3012
rect 546773 3009 546785 3012
rect 546819 3009 546831 3043
rect 546773 3003 546831 3009
rect 548610 3000 548616 3052
rect 548668 3040 548674 3052
rect 582190 3040 582196 3052
rect 548668 3012 582196 3040
rect 548668 3000 548674 3012
rect 582190 3000 582196 3012
rect 582248 3000 582254 3052
rect 582377 3043 582435 3049
rect 582377 3009 582389 3043
rect 582423 3040 582435 3043
rect 583386 3040 583392 3052
rect 582423 3012 583392 3040
rect 582423 3009 582435 3012
rect 582377 3003 582435 3009
rect 583386 3000 583392 3012
rect 583444 3000 583450 3052
rect 539560 2944 542124 2972
rect 539560 2932 539566 2944
rect 545758 2932 545764 2984
rect 545816 2972 545822 2984
rect 552661 2975 552719 2981
rect 552661 2972 552673 2975
rect 545816 2944 552673 2972
rect 545816 2932 545822 2944
rect 552661 2941 552673 2944
rect 552707 2941 552719 2975
rect 552661 2935 552719 2941
rect 552753 2975 552811 2981
rect 552753 2941 552765 2975
rect 552799 2972 552811 2975
rect 571518 2972 571524 2984
rect 552799 2944 571524 2972
rect 552799 2941 552811 2944
rect 552753 2935 552811 2941
rect 571518 2932 571524 2944
rect 571576 2932 571582 2984
rect 48958 2864 48964 2916
rect 49016 2904 49022 2916
rect 49602 2904 49608 2916
rect 49016 2876 49608 2904
rect 49016 2864 49022 2876
rect 49602 2864 49608 2876
rect 49660 2864 49666 2916
rect 84470 2864 84476 2916
rect 84528 2904 84534 2916
rect 85482 2904 85488 2916
rect 84528 2876 85488 2904
rect 84528 2864 84534 2876
rect 85482 2864 85488 2876
rect 85540 2864 85546 2916
rect 292574 2864 292580 2916
rect 292632 2904 292638 2916
rect 293954 2904 293960 2916
rect 292632 2876 293960 2904
rect 292632 2864 292638 2876
rect 293954 2864 293960 2876
rect 294012 2864 294018 2916
rect 324222 2864 324228 2916
rect 324280 2904 324286 2916
rect 326798 2904 326804 2916
rect 324280 2876 326804 2904
rect 324280 2864 324286 2876
rect 326798 2864 326804 2876
rect 326856 2864 326862 2916
rect 408310 2864 408316 2916
rect 408368 2904 408374 2916
rect 424962 2904 424968 2916
rect 408368 2876 424968 2904
rect 408368 2864 408374 2876
rect 424962 2864 424968 2876
rect 425020 2864 425026 2916
rect 452562 2864 452568 2916
rect 452620 2904 452626 2916
rect 475746 2904 475752 2916
rect 452620 2876 475752 2904
rect 452620 2864 452626 2876
rect 475746 2864 475752 2876
rect 475804 2864 475810 2916
rect 497458 2864 497464 2916
rect 497516 2904 497522 2916
rect 518342 2904 518348 2916
rect 497516 2876 518348 2904
rect 497516 2864 497522 2876
rect 518342 2864 518348 2876
rect 518400 2864 518406 2916
rect 522298 2864 522304 2916
rect 522356 2904 522362 2916
rect 536098 2904 536104 2916
rect 522356 2876 536104 2904
rect 522356 2864 522362 2876
rect 536098 2864 536104 2876
rect 536156 2864 536162 2916
rect 540238 2864 540244 2916
rect 540296 2904 540302 2916
rect 564434 2904 564440 2916
rect 540296 2876 552704 2904
rect 540296 2864 540302 2876
rect 136450 2796 136456 2848
rect 136508 2836 136514 2848
rect 139394 2836 139400 2848
rect 136508 2808 139400 2836
rect 136508 2796 136514 2808
rect 139394 2796 139400 2808
rect 139452 2796 139458 2848
rect 294874 2796 294880 2848
rect 294932 2836 294938 2848
rect 295426 2836 295432 2848
rect 294932 2808 295432 2836
rect 294932 2796 294938 2808
rect 295426 2796 295432 2808
rect 295484 2796 295490 2848
rect 447042 2796 447048 2848
rect 447100 2836 447106 2848
rect 469858 2836 469864 2848
rect 447100 2808 469864 2836
rect 447100 2796 447106 2808
rect 469858 2796 469864 2808
rect 469916 2796 469922 2848
rect 541618 2796 541624 2848
rect 541676 2836 541682 2848
rect 552569 2839 552627 2845
rect 552569 2836 552581 2839
rect 541676 2808 552581 2836
rect 541676 2796 541682 2808
rect 552569 2805 552581 2808
rect 552615 2805 552627 2839
rect 552569 2799 552627 2805
rect 552676 2768 552704 2876
rect 557506 2876 564440 2904
rect 557506 2836 557534 2876
rect 564434 2864 564440 2876
rect 564492 2864 564498 2916
rect 552860 2808 557534 2836
rect 552860 2768 552888 2808
rect 552676 2740 552888 2768
<< via1 >>
rect 273168 700952 273220 701004
rect 397460 700952 397512 701004
rect 154120 700884 154172 700936
rect 268384 700884 268436 700936
rect 278688 700884 278740 700936
rect 413652 700884 413704 700936
rect 137836 700816 137888 700868
rect 325700 700816 325752 700868
rect 331864 700816 331916 700868
rect 494796 700816 494848 700868
rect 89168 700748 89220 700800
rect 93124 700748 93176 700800
rect 260748 700748 260800 700800
rect 462320 700748 462372 700800
rect 218980 700680 219032 700732
rect 255964 700680 256016 700732
rect 264888 700680 264940 700732
rect 478512 700680 478564 700732
rect 105452 700612 105504 700664
rect 333980 700612 334032 700664
rect 72976 700544 73028 700596
rect 338120 700544 338172 700596
rect 246948 700476 247000 700528
rect 527180 700476 527232 700528
rect 24308 700408 24360 700460
rect 65524 700408 65576 700460
rect 170312 700408 170364 700460
rect 180064 700408 180116 700460
rect 235172 700408 235224 700460
rect 242164 700408 242216 700460
rect 251088 700408 251140 700460
rect 543464 700408 543516 700460
rect 40500 700340 40552 700392
rect 347780 700340 347832 700392
rect 8116 700272 8168 700324
rect 351920 700272 351972 700324
rect 400864 700272 400916 700324
rect 429844 700272 429896 700324
rect 538864 700272 538916 700324
rect 559656 700272 559708 700324
rect 202788 700204 202840 700256
rect 311900 700204 311952 700256
rect 324964 700204 325016 700256
rect 364984 700204 365036 700256
rect 291108 700136 291160 700188
rect 348792 700136 348844 700188
rect 286968 700068 287020 700120
rect 332508 700068 332560 700120
rect 267648 700000 267700 700052
rect 299480 700000 299532 700052
rect 283840 699932 283892 699984
rect 303620 699932 303672 699984
rect 234528 696940 234580 696992
rect 580172 696940 580224 696992
rect 238668 683204 238720 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 360200 683136 360252 683188
rect 3516 670692 3568 670744
rect 61384 670692 61436 670744
rect 230388 670692 230440 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 364340 656888 364392 656940
rect 220728 643084 220780 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 374000 632068 374052 632120
rect 224868 630640 224920 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 68284 618264 68336 618316
rect 216588 616836 216640 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 378140 605820 378192 605872
rect 208308 590656 208360 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 386420 579640 386472 579692
rect 212448 576852 212500 576904
rect 580172 576852 580224 576904
rect 202788 563048 202840 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 391940 553392 391992 553444
rect 282276 551284 282328 551336
rect 324964 551284 325016 551336
rect 268384 550536 268436 550588
rect 329932 550536 329984 550588
rect 242164 550468 242216 550520
rect 307944 550468 307996 550520
rect 255780 550400 255832 550452
rect 331864 550400 331916 550452
rect 268936 550332 268988 550384
rect 400864 550332 400916 550384
rect 180064 550264 180116 550316
rect 321560 550264 321612 550316
rect 93124 550196 93176 550248
rect 343180 550196 343232 550248
rect 65524 550128 65576 550180
rect 356428 550128 356480 550180
rect 242532 550060 242584 550112
rect 538864 550060 538916 550112
rect 61384 549992 61436 550044
rect 370044 549992 370096 550044
rect 68284 549924 68336 549976
rect 382832 549924 382884 549976
rect 3516 549856 3568 549908
rect 396172 549856 396224 549908
rect 255964 549788 256016 549840
rect 316776 549788 316828 549840
rect 295248 549720 295300 549772
rect 299572 549720 299624 549772
rect 172060 549176 172112 549228
rect 431316 549176 431368 549228
rect 198556 549108 198608 549160
rect 554044 549108 554096 549160
rect 40868 549040 40920 549092
rect 404820 549040 404872 549092
rect 180708 548972 180760 549024
rect 565176 548972 565228 549024
rect 132408 548904 132460 548956
rect 180800 548904 180852 548956
rect 185308 548904 185360 548956
rect 576216 548904 576268 548956
rect 11796 548836 11848 548888
rect 409236 548836 409288 548888
rect 167736 548768 167788 548820
rect 574836 548768 574888 548820
rect 150072 548700 150124 548752
rect 561036 548700 561088 548752
rect 154304 548632 154356 548684
rect 573456 548632 573508 548684
rect 40684 548564 40736 548616
rect 462504 548564 462556 548616
rect 17316 548496 17368 548548
rect 448888 548496 448940 548548
rect 22744 548428 22796 548480
rect 470876 548428 470928 548480
rect 471520 548428 471572 548480
rect 541348 548428 541400 548480
rect 25596 548360 25648 548412
rect 475292 548360 475344 548412
rect 29644 548292 29696 548344
rect 488540 548292 488592 548344
rect 101680 548224 101732 548276
rect 562324 548224 562376 548276
rect 15936 548156 15988 548208
rect 484400 548156 484452 548208
rect 32404 548088 32456 548140
rect 501696 548088 501748 548140
rect 17224 548020 17276 548072
rect 497280 548020 497332 548072
rect 75276 547952 75328 548004
rect 558184 547952 558236 548004
rect 25504 547884 25556 547936
rect 514852 547884 514904 547936
rect 189724 547748 189776 547800
rect 548616 547748 548668 547800
rect 35256 547680 35308 547732
rect 414112 547680 414164 547732
rect 36636 547612 36688 547664
rect 426808 547612 426860 547664
rect 35164 547544 35216 547596
rect 431224 547544 431276 547596
rect 431316 547544 431368 547596
rect 580448 547544 580500 547596
rect 39396 547476 39448 547528
rect 440240 547476 440292 547528
rect 39304 547408 39356 547460
rect 457628 547408 457680 547460
rect 33784 547340 33836 547392
rect 453212 547340 453264 547392
rect 136916 547272 136968 547324
rect 558276 547272 558328 547324
rect 123668 547204 123720 547256
rect 556896 547204 556948 547256
rect 110328 547136 110380 547188
rect 555516 547136 555568 547188
rect 97264 547068 97316 547120
rect 551376 547068 551428 547120
rect 83924 547000 83976 547052
rect 544384 547000 544436 547052
rect 4896 546932 4948 546984
rect 466460 546932 466512 546984
rect 7656 546864 7708 546916
rect 479708 546864 479760 546916
rect 88248 546796 88300 546848
rect 560944 546796 560996 546848
rect 70860 546728 70912 546780
rect 548524 546728 548576 546780
rect 11704 546660 11756 546712
rect 492864 546660 492916 546712
rect 21364 546592 21416 546644
rect 506572 546592 506624 546644
rect 62028 546524 62080 546576
rect 556804 546524 556856 546576
rect 4804 546456 4856 546508
rect 519268 546456 519320 546508
rect 180800 546388 180852 546440
rect 580264 546388 580316 546440
rect 194140 546320 194192 546372
rect 544476 546320 544528 546372
rect 33876 546252 33928 546304
rect 400404 546252 400456 546304
rect 176154 546184 176206 546236
rect 545856 546184 545908 546236
rect 40776 546116 40828 546168
rect 418160 546116 418212 546168
rect 163320 546048 163372 546100
rect 562416 546048 562468 546100
rect 145656 545980 145708 546032
rect 547236 545980 547288 546032
rect 36544 545912 36596 545964
rect 444472 545912 444524 545964
rect 10324 545844 10376 545896
rect 422484 545844 422536 545896
rect 14556 545776 14608 545828
rect 435640 545776 435692 545828
rect 158720 545708 158772 545760
rect 580356 545708 580408 545760
rect 141240 545640 141292 545692
rect 569316 545640 569368 545692
rect 128084 545572 128136 545624
rect 566556 545572 566608 545624
rect 114836 545504 114888 545556
rect 565084 545504 565136 545556
rect 57612 545368 57664 545420
rect 66260 545368 66312 545420
rect 119252 545436 119304 545488
rect 576124 545436 576176 545488
rect 79600 545368 79652 545420
rect 92848 545368 92900 545420
rect 106096 545368 106148 545420
rect 574744 545368 574796 545420
rect 573364 545300 573416 545352
rect 545764 545232 545816 545284
rect 569224 545164 569276 545216
rect 566464 545096 566516 545148
rect 544476 538160 544528 538212
rect 580172 538160 580224 538212
rect 3332 528504 3384 528556
rect 33876 528504 33928 528556
rect 554044 525716 554096 525768
rect 580172 525716 580224 525768
rect 3148 516060 3200 516112
rect 11796 516060 11848 516112
rect 548616 511912 548668 511964
rect 580172 511912 580224 511964
rect 2964 502256 3016 502308
rect 40868 502256 40920 502308
rect 565176 485732 565228 485784
rect 580172 485732 580224 485784
rect 3240 476008 3292 476060
rect 35256 476008 35308 476060
rect 576216 471928 576268 471980
rect 580172 471928 580224 471980
rect 3056 463632 3108 463684
rect 10324 463632 10376 463684
rect 545856 458124 545908 458176
rect 580172 458124 580224 458176
rect 3332 449828 3384 449880
rect 40776 449828 40828 449880
rect 574836 431876 574888 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 36636 423580 36688 423632
rect 2964 411204 3016 411256
rect 14556 411204 14608 411256
rect 562416 405628 562468 405680
rect 580172 405628 580224 405680
rect 3332 398760 3384 398812
rect 35164 398760 35216 398812
rect 573456 379448 573508 379500
rect 580172 379448 580224 379500
rect 3332 372512 3384 372564
rect 39396 372512 39448 372564
rect 3332 358708 3384 358760
rect 17316 358708 17368 358760
rect 561036 353200 561088 353252
rect 580172 353200 580224 353252
rect 3332 346332 3384 346384
rect 36544 346332 36596 346384
rect 569316 325592 569368 325644
rect 579896 325592 579948 325644
rect 3332 320084 3384 320136
rect 33784 320084 33836 320136
rect 547236 313216 547288 313268
rect 580172 313216 580224 313268
rect 3332 306280 3384 306332
rect 40684 306280 40736 306332
rect 558276 299412 558328 299464
rect 579620 299412 579672 299464
rect 3332 293904 3384 293956
rect 39304 293904 39356 293956
rect 566556 273164 566608 273216
rect 579896 273164 579948 273216
rect 2780 267248 2832 267300
rect 4896 267248 4948 267300
rect 3148 255212 3200 255264
rect 25596 255212 25648 255264
rect 556896 245556 556948 245608
rect 580172 245556 580224 245608
rect 3240 241408 3292 241460
rect 22744 241408 22796 241460
rect 565084 233180 565136 233232
rect 579988 233180 580040 233232
rect 576124 219376 576176 219428
rect 580172 219376 580224 219428
rect 3332 214956 3384 215008
rect 7656 214956 7708 215008
rect 555516 206932 555568 206984
rect 579804 206932 579856 206984
rect 3056 202784 3108 202836
rect 29644 202784 29696 202836
rect 562324 193128 562376 193180
rect 580172 193128 580224 193180
rect 3148 188980 3200 189032
rect 15936 188980 15988 189032
rect 574744 179324 574796 179376
rect 580172 179324 580224 179376
rect 551376 166948 551428 167000
rect 580172 166948 580224 167000
rect 3332 164160 3384 164212
rect 11704 164160 11756 164212
rect 560944 153144 560996 153196
rect 580172 153144 580224 153196
rect 3608 150356 3660 150408
rect 32404 150356 32456 150408
rect 573364 139340 573416 139392
rect 580172 139340 580224 139392
rect 3332 137912 3384 137964
rect 17224 137912 17276 137964
rect 544384 126896 544436 126948
rect 580172 126896 580224 126948
rect 558184 113092 558236 113144
rect 579804 113092 579856 113144
rect 3148 111732 3200 111784
rect 21364 111732 21416 111784
rect 569224 100648 569276 100700
rect 580172 100648 580224 100700
rect 3240 97928 3292 97980
rect 25504 97928 25556 97980
rect 548524 86912 548576 86964
rect 580172 86912 580224 86964
rect 3332 85484 3384 85536
rect 18604 85484 18656 85536
rect 556804 73108 556856 73160
rect 580172 73108 580224 73160
rect 2780 71612 2832 71664
rect 4804 71612 4856 71664
rect 566464 60664 566516 60716
rect 580172 60664 580224 60716
rect 545764 46860 545816 46912
rect 580172 46860 580224 46912
rect 3516 45500 3568 45552
rect 7564 45500 7616 45552
rect 133972 41828 134024 41880
rect 135122 41828 135174 41880
rect 20628 39992 20680 40044
rect 58716 39992 58768 40044
rect 75828 39992 75880 40044
rect 106556 39992 106608 40044
rect 110328 39992 110380 40044
rect 136088 39992 136140 40044
rect 136548 39992 136600 40044
rect 158444 39992 158496 40044
rect 158628 39992 158680 40044
rect 177764 39992 177816 40044
rect 177948 39992 178000 40044
rect 180064 39992 180116 40044
rect 180892 39992 180944 40044
rect 195152 39992 195204 40044
rect 200028 39992 200080 40044
rect 213460 39992 213512 40044
rect 223488 39992 223540 40044
rect 233792 39992 233844 40044
rect 242808 39992 242860 40044
rect 250076 39992 250128 40044
rect 253848 39992 253900 40044
rect 260288 39992 260340 40044
rect 277308 39992 277360 40044
rect 279608 39992 279660 40044
rect 286968 39992 287020 40044
rect 288808 39992 288860 40044
rect 315304 39992 315356 40044
rect 316132 39992 316184 40044
rect 509792 39992 509844 40044
rect 538312 39992 538364 40044
rect 565084 39992 565136 40044
rect 26148 39924 26200 39976
rect 63776 39924 63828 39976
rect 74448 39924 74500 39976
rect 105544 39924 105596 39976
rect 107568 39924 107620 39976
rect 134064 39924 134116 39976
rect 144828 39924 144880 39976
rect 166632 39924 166684 39976
rect 169576 39924 169628 39976
rect 186964 39924 187016 39976
rect 190368 39924 190420 39976
rect 205272 39924 205324 39976
rect 205548 39924 205600 39976
rect 218520 39924 218572 39976
rect 222108 39924 222160 39976
rect 232780 39924 232832 39976
rect 275928 39924 275980 39976
rect 278596 39924 278648 39976
rect 285588 39924 285640 39976
rect 287796 39924 287848 39976
rect 495532 39924 495584 39976
rect 23388 39856 23440 39908
rect 61752 39856 61804 39908
rect 68928 39856 68980 39908
rect 100392 39856 100444 39908
rect 103428 39856 103480 39908
rect 129924 39856 129976 39908
rect 142068 39856 142120 39908
rect 163504 39856 163556 39908
rect 165528 39856 165580 39908
rect 183928 39856 183980 39908
rect 187608 39856 187660 39908
rect 203248 39856 203300 39908
rect 204168 39856 204220 39908
rect 217508 39856 217560 39908
rect 217968 39856 218020 39908
rect 228732 39856 228784 39908
rect 235908 39856 235960 39908
rect 244004 39856 244056 39908
rect 513840 39924 513892 39976
rect 524972 39924 525024 39976
rect 532240 39924 532292 39976
rect 560944 39924 560996 39976
rect 515404 39856 515456 39908
rect 540428 39856 540480 39908
rect 542360 39856 542412 39908
rect 548616 39856 548668 39908
rect 19248 39788 19300 39840
rect 57704 39788 57756 39840
rect 60648 39788 60700 39840
rect 93308 39788 93360 39840
rect 95148 39788 95200 39840
rect 123852 39788 123904 39840
rect 124128 39788 124180 39840
rect 148232 39788 148284 39840
rect 153016 39788 153068 39840
rect 173716 39788 173768 39840
rect 173808 39788 173860 39840
rect 191012 39788 191064 39840
rect 195888 39788 195940 39840
rect 210424 39788 210476 39840
rect 211068 39788 211120 39840
rect 222568 39788 222620 39840
rect 224868 39788 224920 39840
rect 234804 39788 234856 39840
rect 237288 39788 237340 39840
rect 246028 39788 246080 39840
rect 248328 39788 248380 39840
rect 255136 39788 255188 39840
rect 501696 39788 501748 39840
rect 532700 39788 532752 39840
rect 535276 39788 535328 39840
rect 562324 39788 562376 39840
rect 9588 39720 9640 39772
rect 49516 39720 49568 39772
rect 63408 39720 63460 39772
rect 96344 39720 96396 39772
rect 106188 39720 106240 39772
rect 132960 39720 133012 39772
rect 139308 39720 139360 39772
rect 161480 39720 161532 39772
rect 162768 39720 162820 39772
rect 181904 39720 181956 39772
rect 184848 39720 184900 39772
rect 200212 39720 200264 39772
rect 201408 39720 201460 39772
rect 214472 39720 214524 39772
rect 219256 39720 219308 39772
rect 229744 39720 229796 39772
rect 230388 39720 230440 39772
rect 239864 39720 239916 39772
rect 241428 39720 241480 39772
rect 249064 39720 249116 39772
rect 257988 39720 258040 39772
rect 263324 39720 263376 39772
rect 498568 39720 498620 39772
rect 518164 39720 518216 39772
rect 526076 39720 526128 39772
rect 558184 39720 558236 39772
rect 10968 39652 11020 39704
rect 50528 39652 50580 39704
rect 67548 39652 67600 39704
rect 99380 39652 99432 39704
rect 100668 39652 100720 39704
rect 127900 39652 127952 39704
rect 135168 39652 135220 39704
rect 157432 39652 157484 39704
rect 160008 39652 160060 39704
rect 178776 39652 178828 39704
rect 180708 39652 180760 39704
rect 197176 39652 197228 39704
rect 198648 39652 198700 39704
rect 212540 39652 212592 39704
rect 219348 39652 219400 39704
rect 230756 39652 230808 39704
rect 233148 39652 233200 39704
rect 241980 39652 242032 39704
rect 244188 39652 244240 39704
rect 252100 39652 252152 39704
rect 267648 39652 267700 39704
rect 271512 39652 271564 39704
rect 488448 39652 488500 39704
rect 497464 39652 497516 39704
rect 512828 39652 512880 39704
rect 16488 39584 16540 39636
rect 55588 39584 55640 39636
rect 64144 39584 64196 39636
rect 69848 39584 69900 39636
rect 70308 39584 70360 39636
rect 102416 39584 102468 39636
rect 103336 39584 103388 39636
rect 130936 39584 130988 39636
rect 137928 39584 137980 39636
rect 160468 39584 160520 39636
rect 164148 39584 164200 39636
rect 182916 39584 182968 39636
rect 183468 39584 183520 39636
rect 199200 39584 199252 39636
rect 202696 39584 202748 39636
rect 216496 39584 216548 39636
rect 216588 39584 216640 39636
rect 227720 39584 227772 39636
rect 231768 39584 231820 39636
rect 240968 39584 241020 39636
rect 264888 39584 264940 39636
rect 269396 39584 269448 39636
rect 464988 39584 465040 39636
rect 490012 39584 490064 39636
rect 491484 39584 491536 39636
rect 512644 39584 512696 39636
rect 515956 39584 516008 39636
rect 541348 39652 541400 39704
rect 548524 39652 548576 39704
rect 544384 39584 544436 39636
rect 13728 39516 13780 39568
rect 53564 39516 53616 39568
rect 53748 39516 53800 39568
rect 87144 39516 87196 39568
rect 88248 39516 88300 39568
rect 117688 39516 117740 39568
rect 119988 39516 120040 39568
rect 145196 39516 145248 39568
rect 146944 39516 146996 39568
rect 154396 39516 154448 39568
rect 167644 39516 167696 39568
rect 169668 39516 169720 39568
rect 187976 39516 188028 39568
rect 188988 39516 189040 39568
rect 204260 39516 204312 39568
rect 206928 39516 206980 39568
rect 219532 39516 219584 39568
rect 220728 39516 220780 39568
rect 231860 39516 231912 39568
rect 234528 39516 234580 39568
rect 242992 39516 243044 39568
rect 245568 39516 245620 39568
rect 253112 39516 253164 39568
rect 256608 39516 256660 39568
rect 262312 39516 262364 39568
rect 477224 39516 477276 39568
rect 502984 39516 503036 39568
rect 503720 39516 503772 39568
rect 522304 39516 522356 39568
rect 523040 39516 523092 39568
rect 556804 39516 556856 39568
rect 12348 39448 12400 39500
rect 51540 39448 51592 39500
rect 56508 39448 56560 39500
rect 90272 39448 90324 39500
rect 92388 39448 92440 39500
rect 120816 39448 120868 39500
rect 121368 39448 121420 39500
rect 146300 39448 146352 39500
rect 148968 39448 149020 39500
rect 169760 39448 169812 39500
rect 171048 39448 171100 39500
rect 189080 39448 189132 39500
rect 194416 39448 194468 39500
rect 208400 39448 208452 39500
rect 215208 39448 215260 39500
rect 226708 39448 226760 39500
rect 235816 39448 235868 39500
rect 245016 39448 245068 39500
rect 246948 39448 247000 39500
rect 254124 39448 254176 39500
rect 255228 39448 255280 39500
rect 261300 39448 261352 39500
rect 267004 39448 267056 39500
rect 270500 39448 270552 39500
rect 332692 39448 332744 39500
rect 336004 39448 336056 39500
rect 480260 39448 480312 39500
rect 507860 39448 507912 39500
rect 516968 39448 517020 39500
rect 550640 39448 550692 39500
rect 6828 39380 6880 39432
rect 47492 39380 47544 39432
rect 57888 39380 57940 39432
rect 91284 39380 91336 39432
rect 99288 39380 99340 39432
rect 126980 39380 127032 39432
rect 132408 39380 132460 39432
rect 155408 39380 155460 39432
rect 155868 39380 155920 39432
rect 175740 39380 175792 39432
rect 179328 39380 179380 39432
rect 196164 39380 196216 39432
rect 197268 39380 197320 39432
rect 211436 39380 211488 39432
rect 213828 39380 213880 39432
rect 225696 39380 225748 39432
rect 229008 39380 229060 39432
rect 238852 39380 238904 39432
rect 244096 39380 244148 39432
rect 251180 39380 251232 39432
rect 434444 39380 434496 39432
rect 443552 39380 443604 39432
rect 458916 39380 458968 39432
rect 483020 39380 483072 39432
rect 483296 39380 483348 39432
rect 512000 39380 512052 39432
rect 520004 39380 520056 39432
rect 554780 39380 554832 39432
rect 4068 39312 4120 39364
rect 45560 39312 45612 39364
rect 49608 39312 49660 39364
rect 84200 39312 84252 39364
rect 85488 39312 85540 39364
rect 114652 39312 114704 39364
rect 117228 39312 117280 39364
rect 142160 39312 142212 39364
rect 144736 39312 144788 39364
rect 165620 39312 165672 39364
rect 166908 39312 166960 39364
rect 184940 39312 184992 39364
rect 186136 39312 186188 39364
rect 202236 39312 202288 39364
rect 210976 39312 211028 39364
rect 223580 39312 223632 39364
rect 227536 39312 227588 39364
rect 237840 39312 237892 39364
rect 238668 39312 238720 39364
rect 247040 39312 247092 39364
rect 277216 39312 277268 39364
rect 280620 39312 280672 39364
rect 343824 39312 343876 39364
rect 349252 39312 349304 39364
rect 437480 39312 437532 39364
rect 454684 39312 454736 39364
rect 455880 39312 455932 39364
rect 465724 39312 465776 39364
rect 474188 39312 474240 39364
rect 31668 39244 31720 39296
rect 68836 39244 68888 39296
rect 71780 39244 71832 39296
rect 73988 39244 74040 39296
rect 75184 39244 75236 39296
rect 82084 39244 82136 39296
rect 28908 39176 28960 39228
rect 65800 39176 65852 39228
rect 68284 39176 68336 39228
rect 35808 39108 35860 39160
rect 71872 39108 71924 39160
rect 72424 39108 72476 39160
rect 73068 39108 73120 39160
rect 39304 39040 39356 39092
rect 75000 39040 75052 39092
rect 81348 39176 81400 39228
rect 111616 39244 111668 39296
rect 113088 39244 113140 39296
rect 139124 39244 139176 39296
rect 143448 39244 143500 39296
rect 164608 39244 164660 39296
rect 172428 39244 172480 39296
rect 190000 39244 190052 39296
rect 193128 39244 193180 39296
rect 207296 39244 207348 39296
rect 208308 39244 208360 39296
rect 220544 39244 220596 39296
rect 227628 39244 227680 39296
rect 236828 39244 236880 39296
rect 510804 39312 510856 39364
rect 543004 39312 543056 39364
rect 543648 39312 543700 39364
rect 500960 39244 501012 39296
rect 528100 39244 528152 39296
rect 540244 39244 540296 39296
rect 547236 39244 547288 39296
rect 78588 39108 78640 39160
rect 108580 39176 108632 39228
rect 114468 39176 114520 39228
rect 140136 39176 140188 39228
rect 140688 39176 140740 39228
rect 162492 39176 162544 39228
rect 168288 39176 168340 39228
rect 185952 39176 186004 39228
rect 191748 39176 191800 39228
rect 206284 39176 206336 39228
rect 209688 39176 209740 39228
rect 221556 39176 221608 39228
rect 226248 39176 226300 39228
rect 235724 39176 235776 39228
rect 274548 39176 274600 39228
rect 277584 39176 277636 39228
rect 534264 39176 534316 39228
rect 541624 39176 541676 39228
rect 84844 39108 84896 39160
rect 112628 39108 112680 39160
rect 115848 39108 115900 39160
rect 141148 39108 141200 39160
rect 147588 39108 147640 39160
rect 168656 39108 168708 39160
rect 175188 39108 175240 39160
rect 192024 39108 192076 39160
rect 194508 39108 194560 39160
rect 209320 39108 209372 39160
rect 212448 39108 212500 39160
rect 224592 39108 224644 39160
rect 44088 38972 44140 39024
rect 79048 38972 79100 39024
rect 82084 39040 82136 39092
rect 109592 39040 109644 39092
rect 111708 39040 111760 39092
rect 137100 39040 137152 39092
rect 137284 39040 137336 39092
rect 138112 39040 138164 39092
rect 153108 39040 153160 39092
rect 172704 39040 172756 39092
rect 177856 39040 177908 39092
rect 194048 39040 194100 39092
rect 202788 39040 202840 39092
rect 215484 39040 215536 39092
rect 252376 39040 252428 39092
rect 259276 39040 259328 39092
rect 259368 39040 259420 39092
rect 264336 39040 264388 39092
rect 269028 39040 269080 39092
rect 273536 39040 273588 39092
rect 85120 38972 85172 39024
rect 91744 38972 91796 39024
rect 118792 38972 118844 39024
rect 119896 38972 119948 39024
rect 144184 38972 144236 39024
rect 150348 38972 150400 39024
rect 170680 38972 170732 39024
rect 176568 38972 176620 39024
rect 193036 38972 193088 39024
rect 240048 38972 240100 39024
rect 248052 38972 248104 39024
rect 251088 38972 251140 39024
rect 257252 38972 257304 39024
rect 260748 38972 260800 39024
rect 265348 38972 265400 39024
rect 271788 38972 271840 39024
rect 275560 38972 275612 39024
rect 282828 38972 282880 39024
rect 284668 38972 284720 39024
rect 284944 38972 284996 39024
rect 285680 38972 285732 39024
rect 289728 38972 289780 39024
rect 290832 38972 290884 39024
rect 296720 38972 296772 39024
rect 297916 38972 297968 39024
rect 303620 38972 303672 39024
rect 304080 38972 304132 39024
rect 307208 38972 307260 39024
rect 307668 38972 307720 39024
rect 311256 38972 311308 39024
rect 311808 38972 311860 39024
rect 313280 38972 313332 39024
rect 314568 38972 314620 39024
rect 316408 38972 316460 39024
rect 317328 38972 317380 39024
rect 317420 38972 317472 39024
rect 318708 38972 318760 39024
rect 320456 38972 320508 39024
rect 321468 38972 321520 39024
rect 323492 38972 323544 39024
rect 324228 38972 324280 39024
rect 324504 38972 324556 39024
rect 325516 38972 325568 39024
rect 326528 38972 326580 39024
rect 326988 38972 327040 39024
rect 327540 38972 327592 39024
rect 328368 38972 328420 39024
rect 328552 38972 328604 39024
rect 329748 38972 329800 39024
rect 330576 38972 330628 39024
rect 331128 38972 331180 39024
rect 331680 38972 331732 39024
rect 332508 38972 332560 39024
rect 333704 38972 333756 39024
rect 334624 38972 334676 39024
rect 334716 38972 334768 39024
rect 335268 38972 335320 39024
rect 335728 38972 335780 39024
rect 336648 38972 336700 39024
rect 338764 38972 338816 39024
rect 339408 38972 339460 39024
rect 339776 38972 339828 39024
rect 340788 38972 340840 39024
rect 342812 38972 342864 39024
rect 343548 38972 343600 39024
rect 345848 38972 345900 39024
rect 346308 38972 346360 39024
rect 346952 38972 347004 39024
rect 347688 38972 347740 39024
rect 347964 38972 348016 39024
rect 348976 38972 349028 39024
rect 349988 38972 350040 39024
rect 350448 38972 350500 39024
rect 351000 38972 351052 39024
rect 351828 38972 351880 39024
rect 352012 38972 352064 39024
rect 353208 38972 353260 39024
rect 354036 38972 354088 39024
rect 354588 38972 354640 39024
rect 355048 38972 355100 39024
rect 355968 38972 356020 39024
rect 356060 38972 356112 39024
rect 357348 38972 357400 39024
rect 358084 38972 358136 39024
rect 358728 38972 358780 39024
rect 359096 38972 359148 39024
rect 360108 38972 360160 39024
rect 363236 38972 363288 39024
rect 364248 38972 364300 39024
rect 366272 38972 366324 39024
rect 367008 38972 367060 39024
rect 367284 38972 367336 39024
rect 368296 38972 368348 39024
rect 369308 38972 369360 39024
rect 369768 38972 369820 39024
rect 370320 38972 370372 39024
rect 371148 38972 371200 39024
rect 371332 38972 371384 39024
rect 372528 38972 372580 39024
rect 373356 38972 373408 39024
rect 373908 38972 373960 39024
rect 374368 38972 374420 39024
rect 375288 38972 375340 39024
rect 377496 38972 377548 39024
rect 378048 38972 378100 39024
rect 378508 38972 378560 39024
rect 379428 38972 379480 39024
rect 379520 38972 379572 39024
rect 380716 38972 380768 39024
rect 382556 38972 382608 39024
rect 383476 38972 383528 39024
rect 385592 38972 385644 39024
rect 386328 38972 386380 39024
rect 386604 38972 386656 39024
rect 387708 38972 387760 39024
rect 388628 38972 388680 39024
rect 389088 38972 389140 39024
rect 389640 38972 389692 39024
rect 390468 38972 390520 39024
rect 390652 38972 390704 39024
rect 391756 38972 391808 39024
rect 392768 38972 392820 39024
rect 393228 38972 393280 39024
rect 393780 38972 393832 39024
rect 394608 38972 394660 39024
rect 396816 38972 396868 39024
rect 397368 38972 397420 39024
rect 397828 38972 397880 39024
rect 398748 38972 398800 39024
rect 398840 38972 398892 39024
rect 400128 38972 400180 39024
rect 401876 38972 401928 39024
rect 402888 38972 402940 39024
rect 404912 38972 404964 39024
rect 405648 38972 405700 39024
rect 405924 38972 405976 39024
rect 407028 38972 407080 39024
rect 409052 38972 409104 39024
rect 409788 38972 409840 39024
rect 410064 38972 410116 39024
rect 411076 38972 411128 39024
rect 412088 38972 412140 39024
rect 412548 38972 412600 39024
rect 413100 38972 413152 39024
rect 413928 38972 413980 39024
rect 414112 38972 414164 39024
rect 415308 38972 415360 39024
rect 416136 38972 416188 39024
rect 416688 38972 416740 39024
rect 417148 38972 417200 39024
rect 418068 38972 418120 39024
rect 418160 38972 418212 39024
rect 419356 38972 419408 39024
rect 421196 38972 421248 39024
rect 422208 38972 422260 39024
rect 424324 38972 424376 39024
rect 424968 38972 425020 39024
rect 425336 38972 425388 39024
rect 426256 38972 426308 39024
rect 428372 38972 428424 39024
rect 429108 38972 429160 39024
rect 429384 38972 429436 39024
rect 430488 38972 430540 39024
rect 431408 38972 431460 39024
rect 431868 38972 431920 39024
rect 432420 38972 432472 39024
rect 433248 38972 433300 39024
rect 433432 38972 433484 39024
rect 434628 38972 434680 39024
rect 435456 38972 435508 39024
rect 436008 38972 436060 39024
rect 436468 38972 436520 39024
rect 437388 38972 437440 39024
rect 439596 38972 439648 39024
rect 440148 38972 440200 39024
rect 440608 38972 440660 39024
rect 441528 38972 441580 39024
rect 441620 38972 441672 39024
rect 442908 38972 442960 39024
rect 443644 38972 443696 39024
rect 444288 38972 444340 39024
rect 447692 38972 447744 39024
rect 448428 38972 448480 39024
rect 448704 38972 448756 39024
rect 449808 38972 449860 39024
rect 450728 38972 450780 39024
rect 451188 38972 451240 39024
rect 451740 38972 451792 39024
rect 452568 38972 452620 39024
rect 452752 38972 452804 39024
rect 453856 38972 453908 39024
rect 454868 38972 454920 39024
rect 455328 38972 455380 39024
rect 456892 38972 456944 39024
rect 457996 38972 458048 39024
rect 459928 38972 459980 39024
rect 460848 38972 460900 39024
rect 460940 38972 460992 39024
rect 462228 38972 462280 39024
rect 462964 38972 463016 39024
rect 463608 38972 463660 39024
rect 467012 38972 467064 39024
rect 467748 38972 467800 39024
rect 468024 38972 468076 39024
rect 469036 38972 469088 39024
rect 471152 38972 471204 39024
rect 471888 38972 471940 39024
rect 475200 38972 475252 39024
rect 476028 38972 476080 39024
rect 476212 38972 476264 39024
rect 477408 38972 477460 39024
rect 478236 38972 478288 39024
rect 478788 38972 478840 39024
rect 479248 38972 479300 39024
rect 480168 38972 480220 39024
rect 482284 38972 482336 39024
rect 482928 38972 482980 39024
rect 484400 38972 484452 39024
rect 485596 38972 485648 39024
rect 486424 38972 486476 39024
rect 487068 38972 487120 39024
rect 487436 38972 487488 39024
rect 488448 38972 488500 39024
rect 492496 38972 492548 39024
rect 493324 38972 493376 39024
rect 494520 38972 494572 39024
rect 495348 38972 495400 39024
rect 497556 38972 497608 39024
rect 498108 38972 498160 39024
rect 502708 38972 502760 39024
rect 503628 38972 503680 39024
rect 505744 38972 505796 39024
rect 506388 38972 506440 39024
rect 506756 38972 506808 39024
rect 507768 38972 507820 39024
rect 514944 38972 514996 39024
rect 516048 38972 516100 39024
rect 517980 38972 518032 39024
rect 518808 38972 518860 39024
rect 518992 38972 519044 39024
rect 520188 38972 520240 39024
rect 522028 38972 522080 39024
rect 522948 38972 523000 39024
rect 525064 38972 525116 39024
rect 525708 38972 525760 39024
rect 529112 38972 529164 39024
rect 529848 38972 529900 39024
rect 530216 38972 530268 39024
rect 531228 38972 531280 39024
rect 533252 38972 533304 39024
rect 533988 38972 534040 39024
rect 537300 38972 537352 39024
rect 538128 38972 538180 39024
rect 540336 38972 540388 39024
rect 545764 38972 545816 39024
rect 45468 38904 45520 38956
rect 80060 38904 80112 38956
rect 88984 38904 89036 38956
rect 115664 38904 115716 38956
rect 118608 38904 118660 38956
rect 143172 38904 143224 38956
rect 154488 38904 154540 38956
rect 174728 38904 174780 38956
rect 182088 38904 182140 38956
rect 198188 38904 198240 38956
rect 252468 38904 252520 38956
rect 258264 38904 258316 38956
rect 263508 38904 263560 38956
rect 268384 38904 268436 38956
rect 270408 38904 270460 38956
rect 274640 38904 274692 38956
rect 281448 38904 281500 38956
rect 283656 38904 283708 38956
rect 288348 38904 288400 38956
rect 289820 38904 289872 38956
rect 319444 38904 319496 38956
rect 321652 38904 321704 38956
rect 394792 38904 394844 38956
rect 395896 38904 395948 38956
rect 444656 38904 444708 38956
rect 445668 38904 445720 38956
rect 463976 38904 464028 38956
rect 464988 38904 465040 38956
rect 499672 38904 499724 38956
rect 500776 38904 500828 38956
rect 32404 38836 32456 38888
rect 66812 38836 66864 38888
rect 71044 38836 71096 38888
rect 72976 38836 73028 38888
rect 73068 38836 73120 38888
rect 94320 38836 94372 38888
rect 95884 38836 95936 38888
rect 121828 38836 121880 38888
rect 125508 38836 125560 38888
rect 149336 38836 149388 38888
rect 151728 38836 151780 38888
rect 171692 38836 171744 38888
rect 186228 38836 186280 38888
rect 201224 38836 201276 38888
rect 249708 38836 249760 38888
rect 256240 38836 256292 38888
rect 262128 38836 262180 38888
rect 267372 38836 267424 38888
rect 268936 38836 268988 38888
rect 272524 38836 272576 38888
rect 273168 38836 273220 38888
rect 276572 38836 276624 38888
rect 336740 38836 336792 38888
rect 338764 38836 338816 38888
rect 536288 38836 536340 38888
rect 536748 38836 536800 38888
rect 50344 38768 50396 38820
rect 78036 38768 78088 38820
rect 80704 38768 80756 38820
rect 103520 38768 103572 38820
rect 122748 38768 122800 38820
rect 147220 38768 147272 38820
rect 157248 38768 157300 38820
rect 176752 38768 176804 38820
rect 260656 38768 260708 38820
rect 266360 38768 266412 38820
rect 362224 38768 362276 38820
rect 362868 38768 362920 38820
rect 375380 38768 375432 38820
rect 376576 38768 376628 38820
rect 381544 38768 381596 38820
rect 382188 38768 382240 38820
rect 400864 38768 400916 38820
rect 401508 38768 401560 38820
rect 420184 38768 420236 38820
rect 420828 38768 420880 38820
rect 490472 38768 490524 38820
rect 491208 38768 491260 38820
rect 521016 38768 521068 38820
rect 521568 38768 521620 38820
rect 42064 38700 42116 38752
rect 46204 38700 46256 38752
rect 59728 38700 59780 38752
rect 61384 38700 61436 38752
rect 62764 38700 62816 38752
rect 54576 38632 54628 38684
rect 57244 38632 57296 38684
rect 81072 38700 81124 38752
rect 89076 38700 89128 38752
rect 97356 38700 97408 38752
rect 106924 38700 106976 38752
rect 124864 38700 124916 38752
rect 129740 38700 129792 38752
rect 131948 38700 132000 38752
rect 146208 38700 146260 38752
rect 161388 38700 161440 38752
rect 179880 38700 179932 38752
rect 280068 38700 280120 38752
rect 282644 38700 282696 38752
rect 312268 38700 312320 38752
rect 313464 38700 313516 38752
rect 472164 38700 472216 38752
rect 473176 38700 473228 38752
rect 493508 38700 493560 38752
rect 493968 38700 494020 38752
rect 71136 38632 71188 38684
rect 88340 38632 88392 38684
rect 278688 38632 278740 38684
rect 281632 38632 281684 38684
rect 41328 38360 41380 38412
rect 77024 38360 77076 38412
rect 34428 38292 34480 38344
rect 70860 38292 70912 38344
rect 4804 38224 4856 38276
rect 42156 38224 42208 38276
rect 55128 38224 55180 38276
rect 89260 38224 89312 38276
rect 91008 38224 91060 38276
rect 119804 38224 119856 38276
rect 7564 38156 7616 38208
rect 44456 38156 44508 38208
rect 48228 38156 48280 38208
rect 83096 38156 83148 38208
rect 84108 38156 84160 38208
rect 113640 38156 113692 38208
rect 30288 38088 30340 38140
rect 67824 38088 67876 38140
rect 79968 38088 80020 38140
rect 110604 38088 110656 38140
rect 130384 38088 130436 38140
rect 152372 38088 152424 38140
rect 17868 38020 17920 38072
rect 56600 38020 56652 38072
rect 59268 38020 59320 38072
rect 92296 38020 92348 38072
rect 133788 38020 133840 38072
rect 156420 38020 156472 38072
rect 22008 37952 22060 38004
rect 60740 37952 60792 38004
rect 66168 37952 66220 38004
rect 98368 37952 98420 38004
rect 129648 37952 129700 38004
rect 153384 37952 153436 38004
rect 8208 37884 8260 37936
rect 48504 37884 48556 37936
rect 52368 37884 52420 37936
rect 86132 37884 86184 37936
rect 86868 37884 86920 37936
rect 116676 37884 116728 37936
rect 126888 37884 126940 37936
rect 150440 37884 150492 37936
rect 93124 37272 93176 37324
rect 95332 37272 95384 37324
rect 104808 36592 104860 36644
rect 129740 36592 129792 36644
rect 37188 36524 37240 36576
rect 71780 36524 71832 36576
rect 97908 36524 97960 36576
rect 125876 36524 125928 36576
rect 131028 36524 131080 36576
rect 146944 36524 146996 36576
rect 3516 33056 3568 33108
rect 14464 33056 14516 33108
rect 555424 33056 555476 33108
rect 580172 33056 580224 33108
rect 14556 32376 14608 32428
rect 42800 32376 42852 32428
rect 51724 30268 51776 30320
rect 52552 30268 52604 30320
rect 102048 26868 102100 26920
rect 128360 26868 128412 26920
rect 551284 20612 551336 20664
rect 579988 20612 580040 20664
rect 129464 8916 129516 8968
rect 150624 8916 150676 8968
rect 3424 6808 3476 6860
rect 15844 6808 15896 6860
rect 547144 6808 547196 6860
rect 580172 6808 580224 6860
rect 562324 6196 562376 6248
rect 572720 6196 572772 6248
rect 529848 6128 529900 6180
rect 565084 6128 565136 6180
rect 576308 6128 576360 6180
rect 565636 6060 565688 6112
rect 556804 5584 556856 5636
rect 558552 5584 558604 5636
rect 560944 5584 560996 5636
rect 569132 5584 569184 5636
rect 454684 5516 454736 5568
rect 459192 5516 459244 5568
rect 558184 5516 558236 5568
rect 562048 5516 562100 5568
rect 515404 5108 515456 5160
rect 526628 5108 526680 5160
rect 487068 5040 487120 5092
rect 515956 5040 516008 5092
rect 518164 5040 518216 5092
rect 530124 5040 530176 5092
rect 465724 4972 465776 5024
rect 480536 4972 480588 5024
rect 489828 4972 489880 5024
rect 519544 4972 519596 5024
rect 443644 4904 443696 4956
rect 455696 4904 455748 4956
rect 462136 4904 462188 4956
rect 487620 4904 487672 4956
rect 493324 4904 493376 4956
rect 523040 4904 523092 4956
rect 525064 4904 525116 4956
rect 547880 4904 547932 4956
rect 429108 4836 429160 4888
rect 448612 4836 448664 4888
rect 469036 4836 469088 4888
rect 494704 4836 494756 4888
rect 505008 4836 505060 4888
rect 537208 4836 537260 4888
rect 72608 4768 72660 4820
rect 103704 4768 103756 4820
rect 139400 4768 139452 4820
rect 158720 4768 158772 4820
rect 431868 4768 431920 4820
rect 452108 4768 452160 4820
rect 471888 4768 471940 4820
rect 498200 4768 498252 4820
rect 507676 4768 507728 4820
rect 540796 4768 540848 4820
rect 62120 4632 62172 4684
rect 64880 4632 64932 4684
rect 128360 4496 128412 4548
rect 133972 4496 134024 4548
rect 502984 4156 503036 4208
rect 505376 4156 505428 4208
rect 543004 4156 543056 4208
rect 544384 4156 544436 4208
rect 2872 4088 2924 4140
rect 7564 4088 7616 4140
rect 50160 4088 50212 4140
rect 41880 4020 41932 4072
rect 50344 4020 50396 4072
rect 348976 4088 349028 4140
rect 355232 4088 355284 4140
rect 358728 4088 358780 4140
rect 367008 4088 367060 4140
rect 380716 4088 380768 4140
rect 391664 4088 391716 4140
rect 398748 4088 398800 4140
rect 413100 4088 413152 4140
rect 413928 4088 413980 4140
rect 430856 4088 430908 4140
rect 433248 4088 433300 4140
rect 453304 4088 453356 4140
rect 455328 4088 455380 4140
rect 479340 4088 479392 4140
rect 481548 4088 481600 4140
rect 510068 4088 510120 4140
rect 518808 4088 518860 4140
rect 552664 4088 552716 4140
rect 20536 3952 20588 4004
rect 46204 3952 46256 4004
rect 14740 3884 14792 3936
rect 42064 3884 42116 3936
rect 45376 3884 45428 3936
rect 57152 3952 57204 4004
rect 60832 4020 60884 4072
rect 72424 4020 72476 4072
rect 82084 4020 82136 4072
rect 84844 4020 84896 4072
rect 340696 4020 340748 4072
rect 346952 4020 347004 4072
rect 361488 4020 361540 4072
rect 370596 4020 370648 4072
rect 380808 4020 380860 4072
rect 393044 4020 393096 4072
rect 395896 4020 395948 4072
rect 409604 4020 409656 4072
rect 411168 4020 411220 4072
rect 428464 4020 428516 4072
rect 430396 4020 430448 4072
rect 450912 4020 450964 4072
rect 453948 4020 454000 4072
rect 478144 4020 478196 4072
rect 485596 4020 485648 4072
rect 513564 4020 513616 4072
rect 525708 4020 525760 4072
rect 560852 4020 560904 4072
rect 68284 3952 68336 4004
rect 92756 3952 92808 4004
rect 95884 3952 95936 4004
rect 368296 3952 368348 4004
rect 377680 3952 377732 4004
rect 379428 3952 379480 4004
rect 390652 3952 390704 4004
rect 391756 3952 391808 4004
rect 404820 3952 404872 4004
rect 405648 3952 405700 4004
rect 421380 3952 421432 4004
rect 422208 3952 422260 4004
rect 440332 3952 440384 4004
rect 441528 3952 441580 4004
rect 462780 3952 462832 4004
rect 463608 3952 463660 4004
rect 488816 3952 488868 4004
rect 491208 3952 491260 4004
rect 520740 3952 520792 4004
rect 521568 3952 521620 4004
rect 556160 3952 556212 4004
rect 52552 3884 52604 3936
rect 53748 3884 53800 3936
rect 75184 3884 75236 3936
rect 343548 3884 343600 3936
rect 349252 3884 349304 3936
rect 357348 3884 357400 3936
rect 364616 3884 364668 3936
rect 369768 3884 369820 3936
rect 379980 3884 380032 3936
rect 382188 3884 382240 3936
rect 394240 3884 394292 3936
rect 397368 3884 397420 3936
rect 411904 3884 411956 3936
rect 419356 3884 419408 3936
rect 436744 3884 436796 3936
rect 438768 3884 438820 3936
rect 460388 3884 460440 3936
rect 464988 3884 465040 3936
rect 489920 3884 489972 3936
rect 493968 3884 494020 3936
rect 524236 3884 524288 3936
rect 524328 3884 524380 3936
rect 559748 3884 559800 3936
rect 32404 3816 32456 3868
rect 64144 3816 64196 3868
rect 71504 3816 71556 3868
rect 80704 3816 80756 3868
rect 344928 3816 344980 3868
rect 351644 3816 351696 3868
rect 351828 3816 351880 3868
rect 358728 3816 358780 3868
rect 362868 3816 362920 3868
rect 371700 3816 371752 3868
rect 372528 3816 372580 3868
rect 382372 3816 382424 3868
rect 383568 3816 383620 3868
rect 396540 3816 396592 3868
rect 401508 3816 401560 3868
rect 416688 3816 416740 3868
rect 420828 3816 420880 3868
rect 439136 3816 439188 3868
rect 442908 3816 442960 3868
rect 463976 3816 464028 3868
rect 467748 3816 467800 3868
rect 493508 3816 493560 3868
rect 495348 3816 495400 3868
rect 525432 3816 525484 3868
rect 531228 3816 531280 3868
rect 566832 3816 566884 3868
rect 35992 3748 36044 3800
rect 71044 3748 71096 3800
rect 353208 3748 353260 3800
rect 359924 3748 359976 3800
rect 360108 3748 360160 3800
rect 368204 3748 368256 3800
rect 368388 3748 368440 3800
rect 378876 3748 378928 3800
rect 383476 3748 383528 3800
rect 395344 3748 395396 3800
rect 395988 3748 396040 3800
rect 410800 3748 410852 3800
rect 415216 3748 415268 3800
rect 433248 3748 433300 3800
rect 436008 3748 436060 3800
rect 456892 3748 456944 3800
rect 457996 3748 458048 3800
rect 481732 3748 481784 3800
rect 485688 3748 485740 3800
rect 514760 3748 514812 3800
rect 527088 3748 527140 3800
rect 563244 3748 563296 3800
rect 26516 3680 26568 3732
rect 62120 3680 62172 3732
rect 64328 3680 64380 3732
rect 89076 3680 89128 3732
rect 354588 3680 354640 3732
rect 362316 3680 362368 3732
rect 365628 3680 365680 3732
rect 375288 3680 375340 3732
rect 376668 3680 376720 3732
rect 388260 3680 388312 3732
rect 393228 3680 393280 3732
rect 407212 3680 407264 3732
rect 411076 3680 411128 3732
rect 427268 3680 427320 3732
rect 427728 3680 427780 3732
rect 447416 3680 447468 3732
rect 448428 3680 448480 3732
rect 471060 3680 471112 3732
rect 473176 3680 473228 3732
rect 499396 3680 499448 3732
rect 500868 3680 500920 3732
rect 532516 3680 532568 3732
rect 533988 3680 534040 3732
rect 570328 3680 570380 3732
rect 1676 3544 1728 3596
rect 14556 3612 14608 3664
rect 39580 3612 39632 3664
rect 75920 3612 75972 3664
rect 96252 3612 96304 3664
rect 106924 3612 106976 3664
rect 108120 3612 108172 3664
rect 12256 3544 12308 3596
rect 572 3476 624 3528
rect 4804 3476 4856 3528
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12348 3476 12400 3528
rect 15936 3544 15988 3596
rect 16488 3544 16540 3596
rect 17040 3544 17092 3596
rect 17868 3544 17920 3596
rect 18236 3544 18288 3596
rect 19248 3544 19300 3596
rect 19432 3544 19484 3596
rect 20628 3544 20680 3596
rect 24216 3544 24268 3596
rect 61384 3544 61436 3596
rect 69112 3544 69164 3596
rect 100760 3544 100812 3596
rect 5264 3408 5316 3460
rect 45744 3408 45796 3460
rect 51356 3476 51408 3528
rect 52368 3476 52420 3528
rect 53748 3476 53800 3528
rect 51724 3408 51776 3460
rect 56048 3408 56100 3460
rect 56508 3408 56560 3460
rect 57244 3408 57296 3460
rect 57888 3408 57940 3460
rect 58440 3408 58492 3460
rect 59268 3408 59320 3460
rect 59636 3408 59688 3460
rect 60648 3408 60700 3460
rect 62028 3408 62080 3460
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 66720 3476 66772 3528
rect 67548 3476 67600 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 73804 3476 73856 3528
rect 74448 3476 74500 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 77392 3476 77444 3528
rect 78588 3476 78640 3528
rect 107660 3544 107712 3596
rect 111616 3544 111668 3596
rect 128360 3612 128412 3664
rect 334624 3612 334676 3664
rect 338672 3612 338724 3664
rect 364248 3612 364300 3664
rect 372896 3612 372948 3664
rect 373908 3612 373960 3664
rect 384764 3612 384816 3664
rect 386328 3612 386380 3664
rect 398932 3612 398984 3664
rect 404268 3612 404320 3664
rect 420184 3612 420236 3664
rect 426256 3612 426308 3664
rect 445024 3612 445076 3664
rect 445668 3612 445720 3664
rect 467472 3612 467524 3664
rect 469128 3612 469180 3664
rect 495900 3612 495952 3664
rect 496728 3612 496780 3664
rect 527824 3612 527876 3664
rect 536748 3612 536800 3664
rect 573916 3612 573968 3664
rect 27712 3340 27764 3392
rect 28908 3340 28960 3392
rect 33600 3340 33652 3392
rect 34428 3340 34480 3392
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 38384 3340 38436 3392
rect 39304 3340 39356 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 43076 3340 43128 3392
rect 44088 3340 44140 3392
rect 44272 3340 44324 3392
rect 45468 3340 45520 3392
rect 46664 3340 46716 3392
rect 71136 3408 71188 3460
rect 76196 3340 76248 3392
rect 105728 3476 105780 3528
rect 106188 3476 106240 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 109316 3476 109368 3528
rect 110328 3476 110380 3528
rect 110512 3476 110564 3528
rect 111708 3476 111760 3528
rect 137284 3544 137336 3596
rect 267740 3544 267792 3596
rect 268936 3544 268988 3596
rect 307760 3544 307812 3596
rect 309048 3544 309100 3596
rect 328368 3544 328420 3596
rect 331588 3544 331640 3596
rect 336648 3544 336700 3596
rect 340972 3544 341024 3596
rect 357256 3544 357308 3596
rect 365812 3544 365864 3596
rect 366916 3544 366968 3596
rect 376484 3544 376536 3596
rect 376576 3544 376628 3596
rect 387156 3544 387208 3596
rect 387616 3544 387668 3596
rect 401324 3544 401376 3596
rect 402796 3544 402848 3596
rect 418988 3544 419040 3596
rect 419448 3544 419500 3596
rect 437940 3544 437992 3596
rect 442816 3544 442868 3596
rect 465172 3544 465224 3596
rect 473268 3544 473320 3596
rect 500592 3544 500644 3596
rect 500776 3544 500828 3596
rect 531320 3544 531372 3596
rect 538128 3544 538180 3596
rect 575112 3544 575164 3596
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 125876 3476 125928 3528
rect 126888 3476 126940 3528
rect 128176 3476 128228 3528
rect 130384 3476 130436 3528
rect 130568 3476 130620 3528
rect 131028 3476 131080 3528
rect 131764 3476 131816 3528
rect 132408 3476 132460 3528
rect 132960 3476 133012 3528
rect 133788 3476 133840 3528
rect 134156 3476 134208 3528
rect 135168 3476 135220 3528
rect 135260 3476 135312 3528
rect 136548 3476 136600 3528
rect 138848 3476 138900 3528
rect 139308 3476 139360 3528
rect 140044 3476 140096 3528
rect 140688 3476 140740 3528
rect 141240 3476 141292 3528
rect 142068 3476 142120 3528
rect 142436 3476 142488 3528
rect 143448 3476 143500 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 149520 3476 149572 3528
rect 150348 3476 150400 3528
rect 150624 3476 150676 3528
rect 151728 3476 151780 3528
rect 151820 3476 151872 3528
rect 153108 3476 153160 3528
rect 155408 3476 155460 3528
rect 155868 3476 155920 3528
rect 156604 3476 156656 3528
rect 157248 3476 157300 3528
rect 157800 3476 157852 3528
rect 158628 3476 158680 3528
rect 158904 3476 158956 3528
rect 160008 3476 160060 3528
rect 160100 3476 160152 3528
rect 161388 3476 161440 3528
rect 163688 3476 163740 3528
rect 164148 3476 164200 3528
rect 166080 3476 166132 3528
rect 166908 3476 166960 3528
rect 167184 3476 167236 3528
rect 168288 3476 168340 3528
rect 168380 3476 168432 3528
rect 169484 3476 169536 3528
rect 171968 3476 172020 3528
rect 172428 3476 172480 3528
rect 173164 3476 173216 3528
rect 173808 3476 173860 3528
rect 174268 3476 174320 3528
rect 175188 3476 175240 3528
rect 175464 3476 175516 3528
rect 176568 3476 176620 3528
rect 176660 3476 176712 3528
rect 177764 3476 177816 3528
rect 180248 3476 180300 3528
rect 180708 3476 180760 3528
rect 181444 3476 181496 3528
rect 182088 3476 182140 3528
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 184940 3476 184992 3528
rect 186228 3476 186280 3528
rect 188528 3476 188580 3528
rect 188988 3476 189040 3528
rect 190828 3476 190880 3528
rect 191748 3476 191800 3528
rect 192024 3476 192076 3528
rect 193128 3476 193180 3528
rect 193220 3476 193272 3528
rect 194324 3476 194376 3528
rect 197912 3476 197964 3528
rect 198648 3476 198700 3528
rect 199108 3476 199160 3528
rect 200028 3476 200080 3528
rect 201500 3476 201552 3528
rect 202788 3476 202840 3528
rect 205088 3476 205140 3528
rect 205548 3476 205600 3528
rect 206192 3476 206244 3528
rect 206928 3476 206980 3528
rect 207388 3476 207440 3528
rect 208308 3476 208360 3528
rect 209780 3476 209832 3528
rect 211068 3476 211120 3528
rect 213368 3476 213420 3528
rect 213828 3476 213880 3528
rect 214472 3476 214524 3528
rect 215208 3476 215260 3528
rect 215668 3476 215720 3528
rect 216588 3476 216640 3528
rect 216864 3476 216916 3528
rect 217968 3476 218020 3528
rect 218060 3476 218112 3528
rect 219164 3476 219216 3528
rect 222752 3476 222804 3528
rect 223488 3476 223540 3528
rect 223948 3476 224000 3528
rect 224868 3476 224920 3528
rect 226340 3476 226392 3528
rect 227628 3476 227680 3528
rect 229836 3476 229888 3528
rect 230388 3476 230440 3528
rect 231032 3476 231084 3528
rect 231768 3476 231820 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 234620 3476 234672 3528
rect 235908 3476 235960 3528
rect 238116 3476 238168 3528
rect 238668 3476 238720 3528
rect 239312 3476 239364 3528
rect 240048 3476 240100 3528
rect 240508 3476 240560 3528
rect 241428 3476 241480 3528
rect 242900 3476 242952 3528
rect 244004 3476 244056 3528
rect 247592 3476 247644 3528
rect 248328 3476 248380 3528
rect 249984 3476 250036 3528
rect 251088 3476 251140 3528
rect 251180 3476 251232 3528
rect 252468 3476 252520 3528
rect 254676 3476 254728 3528
rect 255228 3476 255280 3528
rect 255872 3476 255924 3528
rect 256608 3476 256660 3528
rect 257068 3476 257120 3528
rect 257988 3476 258040 3528
rect 258264 3476 258316 3528
rect 259368 3476 259420 3528
rect 259460 3476 259512 3528
rect 260748 3476 260800 3528
rect 262956 3476 263008 3528
rect 263508 3476 263560 3528
rect 264152 3476 264204 3528
rect 264888 3476 264940 3528
rect 266544 3476 266596 3528
rect 267648 3476 267700 3528
rect 272432 3476 272484 3528
rect 273168 3476 273220 3528
rect 273628 3476 273680 3528
rect 274548 3476 274600 3528
rect 274824 3476 274876 3528
rect 275928 3476 275980 3528
rect 280712 3476 280764 3528
rect 281448 3476 281500 3528
rect 281908 3476 281960 3528
rect 282828 3476 282880 3528
rect 287796 3476 287848 3528
rect 288348 3476 288400 3528
rect 288992 3476 289044 3528
rect 289728 3476 289780 3528
rect 290188 3476 290240 3528
rect 291292 3476 291344 3528
rect 291384 3476 291436 3528
rect 292488 3476 292540 3528
rect 293684 3476 293736 3528
rect 294236 3476 294288 3528
rect 296076 3476 296128 3528
rect 296628 3476 296680 3528
rect 300952 3476 301004 3528
rect 301964 3476 302016 3528
rect 302240 3476 302292 3528
rect 303160 3476 303212 3528
rect 309140 3476 309192 3528
rect 310244 3476 310296 3528
rect 310428 3476 310480 3528
rect 311440 3476 311492 3528
rect 311808 3476 311860 3528
rect 312636 3476 312688 3528
rect 314568 3476 314620 3528
rect 315028 3476 315080 3528
rect 317328 3476 317380 3528
rect 318524 3476 318576 3528
rect 318708 3476 318760 3528
rect 319720 3476 319772 3528
rect 329748 3476 329800 3528
rect 332692 3476 332744 3528
rect 336004 3476 336056 3528
rect 337476 3476 337528 3528
rect 342076 3476 342128 3528
rect 348056 3476 348108 3528
rect 350448 3476 350500 3528
rect 357532 3476 357584 3528
rect 360016 3476 360068 3528
rect 369400 3476 369452 3528
rect 372436 3476 372488 3528
rect 383568 3476 383620 3528
rect 384948 3476 385000 3528
rect 397736 3476 397788 3528
rect 400036 3476 400088 3528
rect 415492 3476 415544 3528
rect 422116 3476 422168 3528
rect 441528 3476 441580 3528
rect 445576 3476 445628 3528
rect 468668 3476 468720 3528
rect 470508 3476 470560 3528
rect 497096 3476 497148 3528
rect 498108 3476 498160 3528
rect 529020 3476 529072 3528
rect 531136 3476 531188 3528
rect 568028 3476 568080 3528
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 83280 3340 83332 3392
rect 84108 3340 84160 3392
rect 85672 3408 85724 3460
rect 88984 3408 89036 3460
rect 90364 3408 90416 3460
rect 91008 3408 91060 3460
rect 91560 3408 91612 3460
rect 92388 3408 92440 3460
rect 97448 3408 97500 3460
rect 97908 3408 97960 3460
rect 98644 3408 98696 3460
rect 99288 3408 99340 3460
rect 99840 3408 99892 3460
rect 100668 3408 100720 3460
rect 101036 3408 101088 3460
rect 102048 3408 102100 3460
rect 89168 3340 89220 3392
rect 91744 3340 91796 3392
rect 93952 3340 94004 3392
rect 122932 3408 122984 3460
rect 161296 3408 161348 3460
rect 180064 3408 180116 3460
rect 189724 3408 189776 3460
rect 190368 3408 190420 3460
rect 265348 3408 265400 3460
rect 267004 3408 267056 3460
rect 325608 3408 325660 3460
rect 329196 3408 329248 3460
rect 331128 3408 331180 3460
rect 335084 3408 335136 3460
rect 335268 3408 335320 3460
rect 339868 3408 339920 3460
rect 353116 3408 353168 3460
rect 361120 3408 361172 3460
rect 364156 3408 364208 3460
rect 374092 3408 374144 3460
rect 378048 3408 378100 3460
rect 389456 3408 389508 3460
rect 391848 3408 391900 3460
rect 406016 3408 406068 3460
rect 406936 3408 406988 3460
rect 423772 3408 423824 3460
rect 426348 3408 426400 3460
rect 446220 3408 446272 3460
rect 449716 3408 449768 3460
rect 473452 3408 473504 3460
rect 477408 3408 477460 3460
rect 504180 3408 504232 3460
rect 506388 3408 506440 3460
rect 538404 3408 538456 3460
rect 540336 3408 540388 3460
rect 543188 3408 543240 3460
rect 544476 3408 544528 3460
rect 546684 3408 546736 3460
rect 577412 3408 577464 3460
rect 114008 3340 114060 3392
rect 114468 3340 114520 3392
rect 115204 3340 115256 3392
rect 115848 3340 115900 3392
rect 116400 3340 116452 3392
rect 117228 3340 117280 3392
rect 117596 3340 117648 3392
rect 118608 3340 118660 3392
rect 118792 3340 118844 3392
rect 119804 3340 119856 3392
rect 122288 3340 122340 3392
rect 122748 3340 122800 3392
rect 329656 3340 329708 3392
rect 333888 3340 333940 3392
rect 339408 3340 339460 3392
rect 344560 3340 344612 3392
rect 347688 3340 347740 3392
rect 354036 3340 354088 3392
rect 371148 3340 371200 3392
rect 381176 3340 381228 3392
rect 387708 3340 387760 3392
rect 400128 3340 400180 3392
rect 400220 3340 400272 3392
rect 414296 3340 414348 3392
rect 415308 3340 415360 3392
rect 432052 3340 432104 3392
rect 437388 3340 437440 3392
rect 457996 3340 458048 3392
rect 458088 3340 458140 3392
rect 482836 3340 482888 3392
rect 482928 3340 482980 3392
rect 511264 3340 511316 3392
rect 511908 3340 511960 3392
rect 545488 3340 545540 3392
rect 547236 3340 547288 3392
rect 550272 3340 550324 3392
rect 578608 3340 578660 3392
rect 93124 3272 93176 3324
rect 196808 3272 196860 3324
rect 197268 3272 197320 3324
rect 221556 3272 221608 3324
rect 222108 3272 222160 3324
rect 271236 3272 271288 3324
rect 271788 3272 271840 3324
rect 276020 3272 276072 3324
rect 277308 3272 277360 3324
rect 279516 3272 279568 3324
rect 280068 3272 280120 3324
rect 305000 3272 305052 3324
rect 305552 3272 305604 3324
rect 325516 3272 325568 3324
rect 328000 3272 328052 3324
rect 338028 3272 338080 3324
rect 343364 3272 343416 3324
rect 375196 3272 375248 3324
rect 385960 3272 386012 3324
rect 389088 3272 389140 3324
rect 402520 3272 402572 3324
rect 402888 3272 402940 3324
rect 417884 3272 417936 3324
rect 418068 3272 418120 3324
rect 435548 3272 435600 3324
rect 440148 3272 440200 3324
rect 461584 3272 461636 3324
rect 462228 3272 462280 3324
rect 486424 3272 486476 3324
rect 488448 3272 488500 3324
rect 517152 3272 517204 3324
rect 520188 3272 520240 3324
rect 553768 3272 553820 3324
rect 28908 3204 28960 3256
rect 32312 3204 32364 3256
rect 183744 3204 183796 3256
rect 184848 3204 184900 3256
rect 200304 3204 200356 3256
rect 201408 3204 201460 3256
rect 225144 3204 225196 3256
rect 226248 3204 226300 3256
rect 322848 3204 322900 3256
rect 325608 3204 325660 3256
rect 338764 3204 338816 3256
rect 342168 3204 342220 3256
rect 390468 3204 390520 3256
rect 403624 3204 403676 3256
rect 412548 3204 412600 3256
rect 429660 3204 429712 3256
rect 430488 3204 430540 3256
rect 449808 3204 449860 3256
rect 453856 3204 453908 3256
rect 476948 3204 477000 3256
rect 478788 3204 478840 3256
rect 506480 3204 506532 3256
rect 512644 3204 512696 3256
rect 521844 3204 521896 3256
rect 522948 3204 523000 3256
rect 78588 3136 78640 3188
rect 81992 3136 82044 3188
rect 241704 3136 241756 3188
rect 242808 3136 242860 3188
rect 321376 3136 321428 3188
rect 324412 3136 324464 3188
rect 326988 3136 327040 3188
rect 330392 3136 330444 3188
rect 332508 3136 332560 3188
rect 336280 3136 336332 3188
rect 407028 3136 407080 3188
rect 422576 3136 422628 3188
rect 424968 3136 425020 3188
rect 443828 3136 443880 3188
rect 451188 3136 451240 3188
rect 474556 3136 474608 3188
rect 476028 3136 476080 3188
rect 502984 3136 503036 3188
rect 507768 3136 507820 3188
rect 539600 3136 539652 3188
rect 548524 3136 548576 3188
rect 102232 3068 102284 3120
rect 103428 3068 103480 3120
rect 126980 3068 127032 3120
rect 129464 3068 129516 3120
rect 246396 3068 246448 3120
rect 246948 3068 247000 3120
rect 349068 3068 349120 3120
rect 356336 3068 356388 3120
rect 394608 3068 394660 3120
rect 408408 3068 408460 3120
rect 423588 3068 423640 3120
rect 442632 3068 442684 3120
rect 449716 3068 449768 3120
rect 472256 3068 472308 3120
rect 480168 3068 480220 3120
rect 507676 3068 507728 3120
rect 516048 3068 516100 3120
rect 549076 3068 549128 3120
rect 557356 3136 557408 3188
rect 581000 3136 581052 3188
rect 25320 3000 25372 3052
rect 26148 3000 26200 3052
rect 143540 3000 143592 3052
rect 144644 3000 144696 3052
rect 164884 3000 164936 3052
rect 165528 3000 165580 3052
rect 208584 3000 208636 3052
rect 209688 3000 209740 3052
rect 248788 3000 248840 3052
rect 249708 3000 249760 3052
rect 283104 3000 283156 3052
rect 284944 3000 284996 3052
rect 318616 3000 318668 3052
rect 320916 3000 320968 3052
rect 340788 3000 340840 3052
rect 345756 3000 345808 3052
rect 346308 3000 346360 3052
rect 352840 3000 352892 3052
rect 355968 3000 356020 3052
rect 363512 3000 363564 3052
rect 416596 3000 416648 3052
rect 434444 3000 434496 3052
rect 444288 3000 444340 3052
rect 466276 3000 466328 3052
rect 466368 3000 466420 3052
rect 492312 3000 492364 3052
rect 509148 3000 509200 3052
rect 541992 3000 542044 3052
rect 284300 2932 284352 2984
rect 285864 2932 285916 2984
rect 314476 2932 314528 2984
rect 316224 2932 316276 2984
rect 321468 2932 321520 2984
rect 323308 2932 323360 2984
rect 409788 2932 409840 2984
rect 426164 2932 426216 2984
rect 434628 2932 434680 2984
rect 454500 2932 454552 2984
rect 460848 2932 460900 2984
rect 485228 2932 485280 2984
rect 503628 2932 503680 2984
rect 534908 2932 534960 2984
rect 539508 2932 539560 2984
rect 548616 3000 548668 3052
rect 582196 3000 582248 3052
rect 583392 3000 583444 3052
rect 545764 2932 545816 2984
rect 571524 2932 571576 2984
rect 48964 2864 49016 2916
rect 49608 2864 49660 2916
rect 84476 2864 84528 2916
rect 85488 2864 85540 2916
rect 292580 2864 292632 2916
rect 293960 2864 294012 2916
rect 324228 2864 324280 2916
rect 326804 2864 326856 2916
rect 408316 2864 408368 2916
rect 424968 2864 425020 2916
rect 452568 2864 452620 2916
rect 475752 2864 475804 2916
rect 497464 2864 497516 2916
rect 518348 2864 518400 2916
rect 522304 2864 522356 2916
rect 536104 2864 536156 2916
rect 540244 2864 540296 2916
rect 136456 2796 136508 2848
rect 139400 2796 139452 2848
rect 294880 2796 294932 2848
rect 295432 2796 295484 2848
rect 447048 2796 447100 2848
rect 469864 2796 469916 2848
rect 541624 2796 541676 2848
rect 564440 2864 564492 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299584 703582 299980 703610
rect 8128 700330 8156 703520
rect 24320 700466 24348 703520
rect 24308 700460 24360 700466
rect 24308 700402 24360 700408
rect 40512 700398 40540 703520
rect 72988 700602 73016 703520
rect 89180 700806 89208 703520
rect 89168 700800 89220 700806
rect 89168 700742 89220 700748
rect 93124 700800 93176 700806
rect 93124 700742 93176 700748
rect 72976 700596 73028 700602
rect 72976 700538 73028 700544
rect 65524 700460 65576 700466
rect 65524 700402 65576 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 61384 670744 61436 670750
rect 61384 670686 61436 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 557534 3464 566879
rect 3436 557506 3556 557534
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3528 549914 3556 557506
rect 61396 550050 61424 670686
rect 65536 550186 65564 700402
rect 68284 618316 68336 618322
rect 68284 618258 68336 618264
rect 65524 550180 65576 550186
rect 65524 550122 65576 550128
rect 61384 550044 61436 550050
rect 61384 549986 61436 549992
rect 68296 549982 68324 618258
rect 93136 550254 93164 700742
rect 105464 700670 105492 703520
rect 137848 700874 137876 703520
rect 154132 700942 154160 703520
rect 154120 700936 154172 700942
rect 154120 700878 154172 700884
rect 137836 700868 137888 700874
rect 137836 700810 137888 700816
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 170324 700466 170352 703520
rect 170312 700460 170364 700466
rect 170312 700402 170364 700408
rect 180064 700460 180116 700466
rect 180064 700402 180116 700408
rect 180076 550322 180104 700402
rect 202800 700262 202828 703520
rect 218992 700738 219020 703520
rect 218980 700732 219032 700738
rect 218980 700674 219032 700680
rect 235184 700466 235212 703520
rect 260748 700800 260800 700806
rect 260748 700742 260800 700748
rect 255964 700732 256016 700738
rect 255964 700674 256016 700680
rect 246948 700528 247000 700534
rect 246948 700470 247000 700476
rect 235172 700460 235224 700466
rect 235172 700402 235224 700408
rect 242164 700460 242216 700466
rect 242164 700402 242216 700408
rect 202788 700256 202840 700262
rect 202788 700198 202840 700204
rect 234528 696992 234580 696998
rect 234528 696934 234580 696940
rect 230388 670744 230440 670750
rect 230388 670686 230440 670692
rect 220728 643136 220780 643142
rect 220728 643078 220780 643084
rect 216588 616888 216640 616894
rect 216588 616830 216640 616836
rect 208308 590708 208360 590714
rect 208308 590650 208360 590656
rect 202788 563100 202840 563106
rect 202788 563042 202840 563048
rect 180064 550316 180116 550322
rect 180064 550258 180116 550264
rect 93124 550248 93176 550254
rect 93124 550190 93176 550196
rect 68284 549976 68336 549982
rect 68284 549918 68336 549924
rect 3516 549908 3568 549914
rect 3516 549850 3568 549856
rect 172060 549228 172112 549234
rect 172060 549170 172112 549176
rect 40868 549092 40920 549098
rect 40868 549034 40920 549040
rect 11796 548888 11848 548894
rect 11796 548830 11848 548836
rect 7562 548040 7618 548049
rect 7562 547975 7618 547984
rect 3514 547904 3570 547913
rect 3514 547839 3570 547848
rect 3422 545728 3478 545737
rect 3422 545663 3478 545672
rect 3332 528556 3384 528562
rect 3332 528498 3384 528504
rect 3344 527921 3372 528498
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3148 516112 3200 516118
rect 3148 516054 3200 516060
rect 3160 514865 3188 516054
rect 3146 514856 3202 514865
rect 3146 514791 3202 514800
rect 2964 502308 3016 502314
rect 2964 502250 3016 502256
rect 2976 501809 3004 502250
rect 2962 501800 3018 501809
rect 2962 501735 3018 501744
rect 3240 476060 3292 476066
rect 3240 476002 3292 476008
rect 3252 475697 3280 476002
rect 3238 475688 3294 475697
rect 3238 475623 3294 475632
rect 3056 463684 3108 463690
rect 3056 463626 3108 463632
rect 3068 462641 3096 463626
rect 3054 462632 3110 462641
rect 3054 462567 3110 462576
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3332 293956 3384 293962
rect 3332 293898 3384 293904
rect 3344 293185 3372 293898
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 2780 267300 2832 267306
rect 2780 267242 2832 267248
rect 2792 267209 2820 267242
rect 2778 267200 2834 267209
rect 2778 267135 2834 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3332 215008 3384 215014
rect 3330 214976 3332 214985
rect 3384 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 137964 3384 137970
rect 3332 137906 3384 137912
rect 3344 136785 3372 137906
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3240 97980 3292 97986
rect 3240 97922 3292 97928
rect 3252 97617 3280 97922
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3332 85536 3384 85542
rect 3332 85478 3384 85484
rect 3344 84697 3372 85478
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 2780 71664 2832 71670
rect 2778 71632 2780 71641
rect 2832 71632 2834 71641
rect 2778 71567 2834 71576
rect 3436 19417 3464 545663
rect 3528 58585 3556 547839
rect 4896 546984 4948 546990
rect 4896 546926 4948 546932
rect 4804 546508 4856 546514
rect 4804 546450 4856 546456
rect 3608 150408 3660 150414
rect 3608 150350 3660 150356
rect 3620 149841 3648 150350
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 4816 71670 4844 546450
rect 4908 267306 4936 546926
rect 4896 267300 4948 267306
rect 4896 267242 4948 267248
rect 4804 71664 4856 71670
rect 4804 71606 4856 71612
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 7576 45558 7604 547975
rect 7656 546916 7708 546922
rect 7656 546858 7708 546864
rect 7668 215014 7696 546858
rect 11704 546712 11756 546718
rect 11704 546654 11756 546660
rect 10324 545896 10376 545902
rect 10324 545838 10376 545844
rect 10336 463690 10364 545838
rect 10324 463684 10376 463690
rect 10324 463626 10376 463632
rect 7656 215008 7708 215014
rect 7656 214950 7708 214956
rect 11716 164218 11744 546654
rect 11808 516118 11836 548830
rect 40684 548616 40736 548622
rect 40684 548558 40736 548564
rect 17316 548548 17368 548554
rect 17316 548490 17368 548496
rect 15936 548208 15988 548214
rect 15936 548150 15988 548156
rect 14462 546544 14518 546553
rect 14462 546479 14518 546488
rect 11796 516112 11848 516118
rect 11796 516054 11848 516060
rect 11704 164212 11756 164218
rect 11704 164154 11756 164160
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 7564 45552 7616 45558
rect 3568 45520 3570 45529
rect 7564 45494 7616 45500
rect 3514 45455 3570 45464
rect 9588 39772 9640 39778
rect 9588 39714 9640 39720
rect 6828 39432 6880 39438
rect 6828 39374 6880 39380
rect 4068 39364 4120 39370
rect 4068 39306 4120 39312
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1688 480 1716 3538
rect 2884 480 2912 4082
rect 4080 480 4108 39306
rect 4804 38276 4856 38282
rect 4804 38218 4856 38224
rect 4816 3534 4844 38218
rect 6840 6914 6868 39374
rect 7564 38208 7616 38214
rect 7564 38150 7616 38156
rect 6472 6886 6868 6914
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6472 480 6500 6886
rect 7576 4146 7604 38150
rect 8208 37936 8260 37942
rect 8208 37878 8260 37884
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 8220 3534 8248 37878
rect 9600 3534 9628 39714
rect 10968 39704 11020 39710
rect 10968 39646 11020 39652
rect 10980 3534 11008 39646
rect 13728 39568 13780 39574
rect 13728 39510 13780 39516
rect 12348 39500 12400 39506
rect 12348 39442 12400 39448
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 7668 480 7696 3470
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 12268 1850 12296 3538
rect 12360 3534 12388 39442
rect 13740 6914 13768 39510
rect 14476 33114 14504 546479
rect 14556 545828 14608 545834
rect 14556 545770 14608 545776
rect 14568 411262 14596 545770
rect 15842 545184 15898 545193
rect 15842 545119 15898 545128
rect 14556 411256 14608 411262
rect 14556 411198 14608 411204
rect 14464 33108 14516 33114
rect 14464 33050 14516 33056
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 13556 6886 13768 6914
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12268 1822 12388 1850
rect 12360 480 12388 1822
rect 13556 480 13584 6886
rect 14568 3670 14596 32370
rect 15856 6866 15884 545119
rect 15948 189038 15976 548150
rect 17224 548072 17276 548078
rect 17224 548014 17276 548020
rect 15936 189032 15988 189038
rect 15936 188974 15988 188980
rect 17236 137970 17264 548014
rect 17328 358766 17356 548490
rect 22744 548480 22796 548486
rect 22744 548422 22796 548428
rect 18602 548176 18658 548185
rect 18602 548111 18658 548120
rect 17316 358760 17368 358766
rect 17316 358702 17368 358708
rect 17224 137964 17276 137970
rect 17224 137906 17276 137912
rect 18616 85542 18644 548111
rect 21364 546644 21416 546650
rect 21364 546586 21416 546592
rect 21376 111790 21404 546586
rect 22756 241466 22784 548422
rect 25596 548412 25648 548418
rect 25596 548354 25648 548360
rect 25504 547936 25556 547942
rect 25504 547878 25556 547884
rect 22744 241460 22796 241466
rect 22744 241402 22796 241408
rect 21364 111784 21416 111790
rect 21364 111726 21416 111732
rect 25516 97986 25544 547878
rect 25608 255270 25636 548354
rect 29644 548344 29696 548350
rect 29644 548286 29696 548292
rect 25596 255264 25648 255270
rect 25596 255206 25648 255212
rect 29656 202842 29684 548286
rect 32404 548140 32456 548146
rect 32404 548082 32456 548088
rect 29644 202836 29696 202842
rect 29644 202778 29696 202784
rect 32416 150414 32444 548082
rect 35256 547732 35308 547738
rect 35256 547674 35308 547680
rect 35164 547596 35216 547602
rect 35164 547538 35216 547544
rect 33784 547392 33836 547398
rect 33784 547334 33836 547340
rect 33796 320142 33824 547334
rect 33876 546304 33928 546310
rect 33876 546246 33928 546252
rect 33888 528562 33916 546246
rect 33876 528556 33928 528562
rect 33876 528498 33928 528504
rect 35176 398818 35204 547538
rect 35268 476066 35296 547674
rect 36636 547664 36688 547670
rect 36636 547606 36688 547612
rect 36544 545964 36596 545970
rect 36544 545906 36596 545912
rect 35256 476060 35308 476066
rect 35256 476002 35308 476008
rect 35164 398812 35216 398818
rect 35164 398754 35216 398760
rect 36556 346390 36584 545906
rect 36648 423638 36676 547606
rect 39396 547528 39448 547534
rect 39396 547470 39448 547476
rect 39304 547460 39356 547466
rect 39304 547402 39356 547408
rect 36636 423632 36688 423638
rect 36636 423574 36688 423580
rect 36544 346384 36596 346390
rect 36544 346326 36596 346332
rect 33784 320136 33836 320142
rect 33784 320078 33836 320084
rect 39316 293962 39344 547402
rect 39408 372570 39436 547470
rect 39396 372564 39448 372570
rect 39396 372506 39448 372512
rect 40696 306338 40724 548558
rect 40776 546168 40828 546174
rect 40776 546110 40828 546116
rect 40788 449886 40816 546110
rect 40880 502314 40908 549034
rect 132408 548956 132460 548962
rect 132408 548898 132460 548904
rect 101680 548276 101732 548282
rect 101680 548218 101732 548224
rect 75276 548004 75328 548010
rect 75276 547946 75328 547952
rect 53194 546816 53250 546825
rect 53194 546751 53250 546760
rect 70860 546780 70912 546786
rect 48778 546680 48834 546689
rect 48778 546615 48834 546624
rect 48792 545986 48820 546615
rect 53208 545986 53236 546751
rect 70860 546722 70912 546728
rect 62028 546576 62080 546582
rect 62028 546518 62080 546524
rect 62040 545986 62068 546518
rect 70872 545986 70900 546722
rect 75288 545986 75316 547946
rect 97264 547120 97316 547126
rect 97264 547062 97316 547068
rect 83924 547052 83976 547058
rect 83924 546994 83976 547000
rect 83936 545986 83964 546994
rect 88248 546848 88300 546854
rect 88248 546790 88300 546796
rect 88260 545986 88288 546790
rect 97276 545986 97304 547062
rect 101692 545986 101720 548218
rect 123668 547256 123720 547262
rect 123668 547198 123720 547204
rect 110328 547188 110380 547194
rect 110328 547130 110380 547136
rect 110340 545986 110368 547130
rect 123680 545986 123708 547198
rect 132420 545986 132448 548898
rect 167736 548820 167788 548826
rect 167736 548762 167788 548768
rect 150072 548752 150124 548758
rect 150072 548694 150124 548700
rect 136916 547324 136968 547330
rect 136916 547266 136968 547272
rect 136928 545986 136956 547266
rect 145656 546032 145708 546038
rect 48484 545958 48820 545986
rect 52900 545958 53236 545986
rect 61732 545958 62068 545986
rect 70564 545958 70900 545986
rect 74980 545958 75316 545986
rect 83720 545958 83964 545986
rect 88136 545958 88288 545986
rect 96968 545958 97304 545986
rect 101384 545958 101720 545986
rect 110124 545958 110368 545986
rect 123372 545958 123708 545986
rect 132204 545958 132448 545986
rect 136620 545958 136956 545986
rect 145360 545980 145656 545986
rect 150084 545986 150112 548694
rect 154304 548684 154356 548690
rect 154304 548626 154356 548632
rect 154316 545986 154344 548626
rect 163320 546100 163372 546106
rect 163320 546042 163372 546048
rect 163332 545986 163360 546042
rect 167748 545986 167776 548762
rect 172072 545986 172100 549170
rect 198556 549160 198608 549166
rect 198556 549102 198608 549108
rect 180708 549024 180760 549030
rect 180708 548966 180760 548972
rect 176154 546236 176206 546242
rect 176154 546178 176206 546184
rect 145360 545974 145708 545980
rect 145360 545958 145696 545974
rect 149776 545958 150112 545986
rect 154192 545958 154344 545986
rect 163024 545958 163360 545986
rect 167440 545958 167776 545986
rect 171764 545958 172100 545986
rect 176166 545972 176194 546178
rect 180720 545986 180748 548966
rect 180800 548956 180852 548962
rect 180800 548898 180852 548904
rect 185308 548956 185360 548962
rect 185308 548898 185360 548904
rect 180812 546446 180840 548898
rect 180800 546440 180852 546446
rect 180800 546382 180852 546388
rect 185320 545986 185348 548898
rect 189724 547800 189776 547806
rect 189724 547742 189776 547748
rect 189736 545986 189764 547742
rect 194140 546372 194192 546378
rect 194140 546314 194192 546320
rect 194152 545986 194180 546314
rect 198568 545986 198596 549102
rect 202800 545986 202828 563042
rect 208320 547874 208348 590650
rect 212448 576904 212500 576910
rect 212448 576846 212500 576852
rect 212460 547874 212488 576846
rect 216600 547874 216628 616830
rect 220740 547874 220768 643078
rect 224868 630692 224920 630698
rect 224868 630634 224920 630640
rect 207400 547846 208348 547874
rect 211816 547846 212488 547874
rect 216232 547846 216628 547874
rect 220648 547846 220768 547874
rect 207400 545986 207428 547846
rect 211816 545986 211844 547846
rect 216232 545986 216260 547846
rect 220648 545986 220676 547846
rect 224880 545986 224908 630634
rect 230400 547874 230428 670686
rect 234540 547874 234568 696934
rect 238668 683256 238720 683262
rect 238668 683198 238720 683204
rect 238680 547874 238708 683198
rect 242176 550526 242204 700402
rect 242164 550520 242216 550526
rect 242164 550462 242216 550468
rect 242532 550112 242584 550118
rect 242532 550054 242584 550060
rect 229480 547846 230428 547874
rect 233804 547846 234568 547874
rect 238220 547846 238708 547874
rect 229480 545986 229508 547846
rect 233804 545986 233832 547846
rect 238220 545986 238248 547846
rect 242544 545986 242572 550054
rect 246960 545986 246988 700470
rect 251088 700460 251140 700466
rect 251088 700402 251140 700408
rect 251100 546258 251128 700402
rect 255780 550452 255832 550458
rect 255780 550394 255832 550400
rect 180596 545958 180748 545986
rect 185012 545958 185348 545986
rect 189428 545958 189764 545986
rect 193844 545958 194180 545986
rect 198260 545958 198596 545986
rect 202584 545958 202828 545986
rect 207000 545958 207428 545986
rect 211416 545958 211844 545986
rect 215832 545958 216260 545986
rect 220248 545958 220676 545986
rect 224664 545958 224908 545986
rect 229080 545958 229508 545986
rect 233404 545958 233832 545986
rect 237820 545958 238248 545986
rect 242236 545958 242572 545986
rect 246652 545958 246988 545986
rect 251054 546230 251128 546258
rect 251054 545972 251082 546230
rect 255792 545986 255820 550394
rect 255976 549846 256004 700674
rect 255964 549840 256016 549846
rect 255964 549782 256016 549788
rect 260760 547874 260788 700742
rect 264888 700732 264940 700738
rect 264888 700674 264940 700680
rect 264900 547874 264928 700674
rect 267660 700058 267688 703520
rect 273168 701004 273220 701010
rect 273168 700946 273220 700952
rect 268384 700936 268436 700942
rect 268384 700878 268436 700884
rect 267648 700052 267700 700058
rect 267648 699994 267700 700000
rect 268396 550594 268424 700878
rect 268384 550588 268436 550594
rect 268384 550530 268436 550536
rect 268936 550384 268988 550390
rect 268936 550326 268988 550332
rect 260300 547846 260788 547874
rect 264624 547846 264928 547874
rect 260300 545986 260328 547846
rect 264624 545986 264652 547846
rect 268948 545986 268976 550326
rect 273180 545986 273208 700946
rect 278688 700936 278740 700942
rect 278688 700878 278740 700884
rect 278700 547874 278728 700878
rect 283852 699990 283880 703520
rect 291108 700188 291160 700194
rect 291108 700130 291160 700136
rect 286968 700120 287020 700126
rect 286968 700062 287020 700068
rect 283840 699984 283892 699990
rect 283840 699926 283892 699932
rect 282276 551336 282328 551342
rect 282276 551278 282328 551284
rect 277872 547846 278728 547874
rect 277872 545986 277900 547846
rect 282288 545986 282316 551278
rect 286980 547874 287008 700062
rect 286704 547846 287008 547874
rect 286704 545986 286732 547846
rect 291120 545986 291148 700130
rect 299480 700052 299532 700058
rect 299480 699994 299532 700000
rect 295248 549772 295300 549778
rect 295248 549714 295300 549720
rect 295260 545986 295288 549714
rect 299492 546258 299520 699994
rect 299584 549778 299612 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 325700 700868 325752 700874
rect 325700 700810 325752 700816
rect 331864 700868 331916 700874
rect 331864 700810 331916 700816
rect 311900 700256 311952 700262
rect 311900 700198 311952 700204
rect 324964 700256 325016 700262
rect 324964 700198 325016 700204
rect 303620 699984 303672 699990
rect 303620 699926 303672 699932
rect 299572 549772 299624 549778
rect 299572 549714 299624 549720
rect 255484 545958 255820 545986
rect 259900 545958 260328 545986
rect 264224 545958 264652 545986
rect 268640 545958 268976 545986
rect 273056 545958 273208 545986
rect 277472 545958 277900 545986
rect 281888 545958 282316 545986
rect 286304 545958 286732 545986
rect 290720 545958 291148 545986
rect 295136 545958 295288 545986
rect 299446 546230 299520 546258
rect 299446 545972 299474 546230
rect 303632 545986 303660 699926
rect 311912 557534 311940 700198
rect 311912 557506 312308 557534
rect 307944 550520 307996 550526
rect 307944 550462 307996 550468
rect 307956 545986 307984 550462
rect 312280 545986 312308 557506
rect 324976 551342 325004 700198
rect 324964 551336 325016 551342
rect 324964 551278 325016 551284
rect 321560 550316 321612 550322
rect 321560 550258 321612 550264
rect 316776 549840 316828 549846
rect 316776 549782 316828 549788
rect 316788 545986 316816 549782
rect 321572 546258 321600 550258
rect 321526 546230 321600 546258
rect 303632 545958 303876 545986
rect 307956 545958 308292 545986
rect 312280 545958 312708 545986
rect 316788 545958 317124 545986
rect 321526 545972 321554 546230
rect 325712 545986 325740 700810
rect 329932 550588 329984 550594
rect 329932 550530 329984 550536
rect 329944 545986 329972 550530
rect 331876 550458 331904 700810
rect 332520 700126 332548 703520
rect 333980 700664 334032 700670
rect 333980 700606 334032 700612
rect 332508 700120 332560 700126
rect 332508 700062 332560 700068
rect 333992 557534 334020 700606
rect 338120 700596 338172 700602
rect 338120 700538 338172 700544
rect 338132 557534 338160 700538
rect 347780 700392 347832 700398
rect 347780 700334 347832 700340
rect 333992 557506 334296 557534
rect 338132 557506 338712 557534
rect 331864 550452 331916 550458
rect 331864 550394 331916 550400
rect 334268 545986 334296 557506
rect 338684 545986 338712 557506
rect 343180 550248 343232 550254
rect 343180 550190 343232 550196
rect 343192 545986 343220 550190
rect 347792 545986 347820 700334
rect 348804 700194 348832 703520
rect 351920 700324 351972 700330
rect 351920 700266 351972 700272
rect 348792 700188 348844 700194
rect 348792 700130 348844 700136
rect 351932 545986 351960 700266
rect 364996 700262 365024 703520
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 413664 700942 413692 703520
rect 413652 700936 413704 700942
rect 413652 700878 413704 700884
rect 429856 700330 429884 703520
rect 462332 700806 462360 703520
rect 462320 700800 462372 700806
rect 462320 700742 462372 700748
rect 478524 700738 478552 703520
rect 494808 700874 494836 703520
rect 494796 700868 494848 700874
rect 494796 700810 494848 700816
rect 478512 700732 478564 700738
rect 478512 700674 478564 700680
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 700330 559696 703520
rect 400864 700324 400916 700330
rect 400864 700266 400916 700272
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 538864 700324 538916 700330
rect 538864 700266 538916 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 364984 700256 365036 700262
rect 364984 700198 365036 700204
rect 360200 683188 360252 683194
rect 360200 683130 360252 683136
rect 360212 557534 360240 683130
rect 364340 656940 364392 656946
rect 364340 656882 364392 656888
rect 364352 557534 364380 656882
rect 374000 632120 374052 632126
rect 374000 632062 374052 632068
rect 360212 557506 360700 557534
rect 364352 557506 365116 557534
rect 356428 550180 356480 550186
rect 356428 550122 356480 550128
rect 356440 545986 356468 550122
rect 360672 545986 360700 557506
rect 365088 545986 365116 557506
rect 370044 550044 370096 550050
rect 370044 549986 370096 549992
rect 325712 545958 325956 545986
rect 329944 545958 330280 545986
rect 334268 545958 334696 545986
rect 338684 545958 339112 545986
rect 343192 545958 343528 545986
rect 347792 545958 347944 545986
rect 351932 545958 352360 545986
rect 356440 545958 356776 545986
rect 360672 545958 361100 545986
rect 365088 545958 365516 545986
rect 158720 545760 158772 545766
rect 140944 545698 141280 545714
rect 158608 545708 158720 545714
rect 370056 545714 370084 549986
rect 374012 545986 374040 632062
rect 378140 605872 378192 605878
rect 378140 605814 378192 605820
rect 378152 557534 378180 605814
rect 386420 579692 386472 579698
rect 386420 579634 386472 579640
rect 386432 557534 386460 579634
rect 378152 557506 378364 557534
rect 386432 557506 387196 557534
rect 378336 545986 378364 557506
rect 382832 549976 382884 549982
rect 382832 549918 382884 549924
rect 382844 545986 382872 549918
rect 387168 545986 387196 557506
rect 391940 553444 391992 553450
rect 391940 553386 391992 553392
rect 391952 546258 391980 553386
rect 400876 550390 400904 700266
rect 400864 550384 400916 550390
rect 400864 550326 400916 550332
rect 538876 550118 538904 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 538864 550112 538916 550118
rect 538864 550054 538916 550060
rect 396172 549908 396224 549914
rect 396172 549850 396224 549856
rect 391906 546230 391980 546258
rect 374012 545958 374348 545986
rect 378336 545958 378764 545986
rect 382844 545958 383180 545986
rect 387168 545958 387596 545986
rect 391906 545972 391934 546230
rect 396184 545986 396212 549850
rect 431316 549228 431368 549234
rect 431316 549170 431368 549176
rect 404820 549092 404872 549098
rect 404820 549034 404872 549040
rect 400404 546304 400456 546310
rect 400404 546246 400456 546252
rect 400416 545986 400444 546246
rect 404832 545986 404860 549034
rect 409236 548888 409288 548894
rect 409236 548830 409288 548836
rect 409248 545986 409276 548830
rect 414112 547732 414164 547738
rect 414112 547674 414164 547680
rect 396184 545958 396336 545986
rect 400416 545958 400752 545986
rect 404832 545958 405168 545986
rect 409248 545958 409584 545986
rect 414124 545850 414152 547674
rect 426808 547664 426860 547670
rect 426808 547606 426860 547612
rect 418160 546168 418212 546174
rect 418160 546110 418212 546116
rect 418172 545986 418200 546110
rect 426820 545986 426848 547606
rect 431328 547602 431356 549170
rect 554044 549160 554096 549166
rect 554044 549102 554096 549108
rect 462504 548616 462556 548622
rect 462504 548558 462556 548564
rect 448888 548548 448940 548554
rect 448888 548490 448940 548496
rect 431224 547596 431276 547602
rect 431224 547538 431276 547544
rect 431316 547596 431368 547602
rect 431316 547538 431368 547544
rect 431236 545986 431264 547538
rect 440240 547528 440292 547534
rect 440240 547470 440292 547476
rect 440252 545986 440280 547470
rect 448900 545986 448928 548490
rect 457628 547460 457680 547466
rect 457628 547402 457680 547408
rect 453212 547392 453264 547398
rect 453212 547334 453264 547340
rect 453224 545986 453252 547334
rect 457640 545986 457668 547402
rect 418172 545958 418416 545986
rect 426820 545958 427156 545986
rect 431236 545958 431572 545986
rect 440252 545958 440404 545986
rect 444484 545970 444820 545986
rect 444472 545964 444820 545970
rect 444524 545958 444820 545964
rect 448900 545958 449236 545986
rect 453224 545958 453560 545986
rect 457640 545958 457976 545986
rect 444472 545906 444524 545912
rect 414000 545822 414152 545850
rect 422484 545896 422536 545902
rect 422536 545844 422740 545850
rect 422484 545838 422740 545844
rect 422496 545822 422740 545838
rect 435652 545834 435988 545850
rect 435640 545828 435988 545834
rect 435692 545822 435988 545828
rect 435640 545770 435692 545776
rect 462516 545714 462544 548558
rect 470876 548480 470928 548486
rect 470876 548422 470928 548428
rect 471520 548480 471572 548486
rect 471520 548422 471572 548428
rect 541348 548480 541400 548486
rect 541348 548422 541400 548428
rect 466460 546984 466512 546990
rect 466460 546926 466512 546932
rect 466472 545986 466500 546926
rect 470888 545986 470916 548422
rect 466472 545958 466808 545986
rect 470888 545958 471224 545986
rect 471532 545737 471560 548422
rect 475292 548412 475344 548418
rect 475292 548354 475344 548360
rect 475304 545986 475332 548354
rect 488540 548344 488592 548350
rect 488540 548286 488592 548292
rect 484400 548208 484452 548214
rect 484400 548150 484452 548156
rect 479708 546916 479760 546922
rect 479708 546858 479760 546864
rect 479720 545986 479748 546858
rect 484412 546258 484440 548150
rect 484366 546230 484440 546258
rect 475304 545958 475640 545986
rect 479720 545958 480056 545986
rect 484366 545972 484394 546230
rect 488552 545986 488580 548286
rect 510618 548176 510674 548185
rect 501696 548140 501748 548146
rect 510618 548111 510674 548120
rect 501696 548082 501748 548088
rect 497280 548072 497332 548078
rect 497280 548014 497332 548020
rect 492864 546712 492916 546718
rect 492864 546654 492916 546660
rect 492876 545986 492904 546654
rect 497292 545986 497320 548014
rect 501708 545986 501736 548082
rect 506572 546644 506624 546650
rect 506572 546586 506624 546592
rect 488552 545958 488796 545986
rect 492876 545958 493212 545986
rect 497292 545958 497628 545986
rect 501708 545958 502044 545986
rect 506584 545850 506612 546586
rect 510632 545986 510660 548111
rect 523682 548040 523738 548049
rect 523682 547975 523738 547984
rect 514852 547936 514904 547942
rect 514852 547878 514904 547884
rect 514864 545986 514892 547878
rect 519268 546508 519320 546514
rect 519268 546450 519320 546456
rect 519280 545986 519308 546450
rect 523696 545986 523724 547975
rect 528098 547904 528154 547913
rect 528098 547839 528154 547848
rect 528112 545986 528140 547839
rect 532698 546544 532754 546553
rect 532698 546479 532754 546488
rect 532712 545986 532740 546479
rect 541360 545986 541388 548422
rect 548616 547800 548668 547806
rect 548616 547742 548668 547748
rect 544384 547052 544436 547058
rect 544384 546994 544436 547000
rect 510632 545958 510876 545986
rect 514864 545958 515200 545986
rect 519280 545958 519616 545986
rect 523696 545958 524032 545986
rect 528112 545958 528448 545986
rect 532712 545958 532864 545986
rect 541360 545958 541696 545986
rect 506460 545822 506612 545850
rect 158608 545702 158772 545708
rect 140944 545692 141292 545698
rect 140944 545686 141240 545692
rect 158608 545686 158760 545702
rect 369932 545686 370084 545714
rect 462392 545686 462544 545714
rect 471518 545728 471574 545737
rect 471518 545663 471574 545672
rect 141240 545634 141292 545640
rect 128084 545624 128136 545630
rect 114540 545562 114876 545578
rect 127788 545572 128084 545578
rect 127788 545566 128136 545572
rect 114540 545556 114888 545562
rect 114540 545550 114836 545556
rect 127788 545550 128124 545566
rect 114836 545498 114888 545504
rect 119252 545488 119304 545494
rect 44454 545456 44510 545465
rect 44160 545414 44454 545442
rect 57316 545426 57652 545442
rect 66148 545426 66300 545442
rect 79304 545426 79640 545442
rect 92552 545426 92888 545442
rect 105800 545426 106136 545442
rect 118956 545436 119252 545442
rect 118956 545430 119304 545436
rect 536930 545456 536986 545465
rect 57316 545420 57664 545426
rect 57316 545414 57612 545420
rect 44454 545391 44510 545400
rect 66148 545420 66312 545426
rect 66148 545414 66260 545420
rect 57612 545362 57664 545368
rect 79304 545420 79652 545426
rect 79304 545414 79600 545420
rect 66260 545362 66312 545368
rect 92552 545420 92900 545426
rect 92552 545414 92848 545420
rect 79600 545362 79652 545368
rect 105800 545420 106148 545426
rect 105800 545414 106096 545420
rect 92848 545362 92900 545368
rect 118956 545414 119292 545430
rect 536986 545414 537280 545442
rect 536930 545391 536986 545400
rect 106096 545362 106148 545368
rect 40868 502308 40920 502314
rect 40868 502250 40920 502256
rect 40776 449880 40828 449886
rect 40776 449822 40828 449828
rect 40684 306332 40736 306338
rect 40684 306274 40736 306280
rect 39304 293956 39356 293962
rect 39304 293898 39356 293904
rect 32404 150408 32456 150414
rect 32404 150350 32456 150356
rect 544396 126954 544424 546994
rect 548524 546780 548576 546786
rect 548524 546722 548576 546728
rect 544476 546372 544528 546378
rect 544476 546314 544528 546320
rect 544488 538218 544516 546314
rect 545856 546236 545908 546242
rect 545856 546178 545908 546184
rect 545764 545284 545816 545290
rect 545764 545226 545816 545232
rect 544476 538212 544528 538218
rect 544476 538154 544528 538160
rect 544384 126948 544436 126954
rect 544384 126890 544436 126896
rect 25504 97980 25556 97986
rect 25504 97922 25556 97928
rect 18604 85536 18656 85542
rect 18604 85478 18656 85484
rect 545776 46918 545804 545226
rect 545868 458182 545896 546178
rect 547236 546032 547288 546038
rect 547236 545974 547288 545980
rect 547142 545320 547198 545329
rect 547142 545255 547198 545264
rect 545856 458176 545908 458182
rect 545856 458118 545908 458124
rect 545764 46912 545816 46918
rect 545764 46854 545816 46860
rect 42168 42078 42504 42106
rect 20628 40044 20680 40050
rect 20628 39986 20680 39992
rect 19248 39840 19300 39846
rect 19248 39782 19300 39788
rect 16488 39636 16540 39642
rect 16488 39578 16540 39584
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14752 480 14780 3878
rect 16500 3602 16528 39578
rect 17868 38072 17920 38078
rect 17868 38014 17920 38020
rect 17880 3602 17908 38014
rect 19260 3602 19288 39782
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 15948 480 15976 3538
rect 17052 480 17080 3538
rect 18248 480 18276 3538
rect 19444 480 19472 3538
rect 20548 1986 20576 3946
rect 20640 3602 20668 39986
rect 26148 39976 26200 39982
rect 26148 39918 26200 39924
rect 23388 39908 23440 39914
rect 23388 39850 23440 39856
rect 22008 38004 22060 38010
rect 22008 37946 22060 37952
rect 22020 6914 22048 37946
rect 23400 6914 23428 39850
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20548 1958 20668 1986
rect 20640 480 20668 1958
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24228 480 24256 3538
rect 26160 3058 26188 39918
rect 31668 39296 31720 39302
rect 31668 39238 31720 39244
rect 28908 39228 28960 39234
rect 28908 39170 28960 39176
rect 26516 3732 26568 3738
rect 26516 3674 26568 3680
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 25332 480 25360 2994
rect 26528 480 26556 3674
rect 28920 3398 28948 39170
rect 30288 38140 30340 38146
rect 30288 38082 30340 38088
rect 30300 6914 30328 38082
rect 31680 6914 31708 39238
rect 35808 39160 35860 39166
rect 35808 39102 35860 39108
rect 32404 38888 32456 38894
rect 32404 38830 32456 38836
rect 32416 6914 32444 38830
rect 34428 38344 34480 38350
rect 34428 38286 34480 38292
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 32324 6886 32444 6914
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27724 480 27752 3334
rect 28908 3256 28960 3262
rect 28908 3198 28960 3204
rect 28920 480 28948 3198
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 32324 3262 32352 6886
rect 32404 3868 32456 3874
rect 32404 3810 32456 3816
rect 32312 3256 32364 3262
rect 32312 3198 32364 3204
rect 32416 480 32444 3810
rect 34440 3398 34468 38286
rect 35820 3398 35848 39102
rect 39304 39092 39356 39098
rect 39304 39034 39356 39040
rect 37188 36576 37240 36582
rect 37188 36518 37240 36524
rect 35992 3800 36044 3806
rect 35992 3742 36044 3748
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 33612 480 33640 3334
rect 34808 480 34836 3334
rect 36004 480 36032 3742
rect 37200 480 37228 36518
rect 39316 3398 39344 39034
rect 42064 38752 42116 38758
rect 42064 38694 42116 38700
rect 41328 38412 41380 38418
rect 41328 38354 41380 38360
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 38396 480 38424 3334
rect 39592 480 39620 3606
rect 41340 3398 41368 38354
rect 41880 4072 41932 4078
rect 41880 4014 41932 4020
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 40696 480 40724 3334
rect 41892 480 41920 4014
rect 42076 3942 42104 38694
rect 42168 38282 42196 42078
rect 43502 41834 43530 42092
rect 44514 41834 44542 42092
rect 42812 41806 43530 41834
rect 44468 41806 44542 41834
rect 45526 41834 45554 42092
rect 46538 41834 46566 42092
rect 47550 41834 47578 42092
rect 48562 41834 48590 42092
rect 49574 41834 49602 42092
rect 50586 41834 50614 42092
rect 51598 41834 51626 42092
rect 52610 41834 52638 42092
rect 53622 41834 53650 42092
rect 54634 41834 54662 42092
rect 55646 41834 55674 42092
rect 56658 41834 56686 42092
rect 57762 41834 57790 42092
rect 58774 41834 58802 42092
rect 59786 41834 59814 42092
rect 60798 41834 60826 42092
rect 61810 41834 61838 42092
rect 62822 41834 62850 42092
rect 63834 41834 63862 42092
rect 45526 41806 45600 41834
rect 42156 38276 42208 38282
rect 42156 38218 42208 38224
rect 42812 32434 42840 41806
rect 44088 39024 44140 39030
rect 44088 38966 44140 38972
rect 42800 32428 42852 32434
rect 42800 32370 42852 32376
rect 42064 3936 42116 3942
rect 42064 3878 42116 3884
rect 44100 3398 44128 38966
rect 44468 38214 44496 41806
rect 45572 39370 45600 41806
rect 45756 41806 46566 41834
rect 47504 41806 47578 41834
rect 48516 41806 48590 41834
rect 49528 41806 49602 41834
rect 50540 41806 50614 41834
rect 51552 41806 51626 41834
rect 52564 41806 52638 41834
rect 53576 41806 53650 41834
rect 54588 41806 54662 41834
rect 55600 41806 55674 41834
rect 56612 41806 56686 41834
rect 57716 41806 57790 41834
rect 58728 41806 58802 41834
rect 59740 41806 59814 41834
rect 60752 41806 60826 41834
rect 61764 41806 61838 41834
rect 62776 41806 62850 41834
rect 63788 41806 63862 41834
rect 64846 41834 64874 42092
rect 65858 41834 65886 42092
rect 66870 41834 66898 42092
rect 67882 41834 67910 42092
rect 68894 41834 68922 42092
rect 69906 41834 69934 42092
rect 70918 41834 70946 42092
rect 71930 41834 71958 42092
rect 73034 41834 73062 42092
rect 74046 41834 74074 42092
rect 75058 41834 75086 42092
rect 76070 41834 76098 42092
rect 77082 41834 77110 42092
rect 78094 41834 78122 42092
rect 79106 41834 79134 42092
rect 80118 41834 80146 42092
rect 81130 41834 81158 42092
rect 82142 41834 82170 42092
rect 83154 41834 83182 42092
rect 64846 41806 64920 41834
rect 45560 39364 45612 39370
rect 45560 39306 45612 39312
rect 45468 38956 45520 38962
rect 45468 38898 45520 38904
rect 44456 38208 44508 38214
rect 44456 38150 44508 38156
rect 45376 3936 45428 3942
rect 45376 3878 45428 3884
rect 43076 3392 43128 3398
rect 43076 3334 43128 3340
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 43088 480 43116 3334
rect 44284 480 44312 3334
rect 45388 1986 45416 3878
rect 45480 3398 45508 38898
rect 45756 3466 45784 41806
rect 47504 39438 47532 41806
rect 47492 39432 47544 39438
rect 47492 39374 47544 39380
rect 46204 38752 46256 38758
rect 46204 38694 46256 38700
rect 46216 4010 46244 38694
rect 48228 38208 48280 38214
rect 48228 38150 48280 38156
rect 48240 6914 48268 38150
rect 48516 37942 48544 41806
rect 49528 39778 49556 41806
rect 49516 39772 49568 39778
rect 49516 39714 49568 39720
rect 50540 39710 50568 41806
rect 50528 39704 50580 39710
rect 50528 39646 50580 39652
rect 51552 39506 51580 41806
rect 51540 39500 51592 39506
rect 51540 39442 51592 39448
rect 49608 39364 49660 39370
rect 49608 39306 49660 39312
rect 48504 37936 48556 37942
rect 48504 37878 48556 37884
rect 47872 6886 48268 6914
rect 46204 4004 46256 4010
rect 46204 3946 46256 3952
rect 45744 3460 45796 3466
rect 45744 3402 45796 3408
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 46664 3392 46716 3398
rect 46664 3334 46716 3340
rect 45388 1958 45508 1986
rect 45480 480 45508 1958
rect 46676 480 46704 3334
rect 47872 480 47900 6886
rect 49620 2922 49648 39306
rect 50344 38820 50396 38826
rect 50344 38762 50396 38768
rect 50160 4140 50212 4146
rect 50160 4082 50212 4088
rect 48964 2916 49016 2922
rect 48964 2858 49016 2864
rect 49608 2916 49660 2922
rect 49608 2858 49660 2864
rect 48976 480 49004 2858
rect 50172 480 50200 4082
rect 50356 4078 50384 38762
rect 52368 37936 52420 37942
rect 52368 37878 52420 37884
rect 51724 30320 51776 30326
rect 51724 30262 51776 30268
rect 50344 4072 50396 4078
rect 50344 4014 50396 4020
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 51368 480 51396 3470
rect 51736 3466 51764 30262
rect 52380 3534 52408 37878
rect 52564 30326 52592 41806
rect 53576 39574 53604 41806
rect 53564 39568 53616 39574
rect 53564 39510 53616 39516
rect 53748 39568 53800 39574
rect 53748 39510 53800 39516
rect 52552 30320 52604 30326
rect 52552 30262 52604 30268
rect 53760 3942 53788 39510
rect 54588 38690 54616 41806
rect 55600 39642 55628 41806
rect 55588 39636 55640 39642
rect 55588 39578 55640 39584
rect 56508 39500 56560 39506
rect 56508 39442 56560 39448
rect 54576 38684 54628 38690
rect 54576 38626 54628 38632
rect 55128 38276 55180 38282
rect 55128 38218 55180 38224
rect 55140 6914 55168 38218
rect 54956 6886 55168 6914
rect 52552 3936 52604 3942
rect 52552 3878 52604 3884
rect 53748 3936 53800 3942
rect 53748 3878 53800 3884
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 51724 3460 51776 3466
rect 51724 3402 51776 3408
rect 52564 480 52592 3878
rect 53748 3528 53800 3534
rect 53748 3470 53800 3476
rect 53760 480 53788 3470
rect 54956 480 54984 6886
rect 56520 3466 56548 39442
rect 56612 38078 56640 41806
rect 57716 39846 57744 41806
rect 58728 40050 58756 41806
rect 58716 40044 58768 40050
rect 58716 39986 58768 39992
rect 57704 39840 57756 39846
rect 57704 39782 57756 39788
rect 57888 39432 57940 39438
rect 57888 39374 57940 39380
rect 57244 38684 57296 38690
rect 57244 38626 57296 38632
rect 56600 38072 56652 38078
rect 56600 38014 56652 38020
rect 57256 6914 57284 38626
rect 57164 6886 57284 6914
rect 57164 4010 57192 6886
rect 57152 4004 57204 4010
rect 57152 3946 57204 3952
rect 57900 3466 57928 39374
rect 59740 38758 59768 41806
rect 60648 39840 60700 39846
rect 60648 39782 60700 39788
rect 59728 38752 59780 38758
rect 59728 38694 59780 38700
rect 59268 38072 59320 38078
rect 59268 38014 59320 38020
rect 59280 3466 59308 38014
rect 60660 3466 60688 39782
rect 60752 38010 60780 41806
rect 61764 39914 61792 41806
rect 61752 39908 61804 39914
rect 61752 39850 61804 39856
rect 62776 38758 62804 41806
rect 63788 39982 63816 41806
rect 63776 39976 63828 39982
rect 63776 39918 63828 39924
rect 63408 39772 63460 39778
rect 63408 39714 63460 39720
rect 61384 38752 61436 38758
rect 61384 38694 61436 38700
rect 62764 38752 62816 38758
rect 62764 38694 62816 38700
rect 60740 38004 60792 38010
rect 60740 37946 60792 37952
rect 60832 4072 60884 4078
rect 60832 4014 60884 4020
rect 56048 3460 56100 3466
rect 56048 3402 56100 3408
rect 56508 3460 56560 3466
rect 56508 3402 56560 3408
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 57888 3460 57940 3466
rect 57888 3402 57940 3408
rect 58440 3460 58492 3466
rect 58440 3402 58492 3408
rect 59268 3460 59320 3466
rect 59268 3402 59320 3408
rect 59636 3460 59688 3466
rect 59636 3402 59688 3408
rect 60648 3460 60700 3466
rect 60648 3402 60700 3408
rect 56060 480 56088 3402
rect 57256 480 57284 3402
rect 58452 480 58480 3402
rect 59648 480 59676 3402
rect 60844 480 60872 4014
rect 61396 3602 61424 38694
rect 63420 6914 63448 39714
rect 64144 39636 64196 39642
rect 64144 39578 64196 39584
rect 63236 6886 63448 6914
rect 62120 4684 62172 4690
rect 62120 4626 62172 4632
rect 62132 3738 62160 4626
rect 62120 3732 62172 3738
rect 62120 3674 62172 3680
rect 61384 3596 61436 3602
rect 61384 3538 61436 3544
rect 62028 3460 62080 3466
rect 62028 3402 62080 3408
rect 62040 480 62068 3402
rect 63236 480 63264 6886
rect 64156 3874 64184 39578
rect 64892 4690 64920 41806
rect 65812 41806 65886 41834
rect 66824 41806 66898 41834
rect 67836 41806 67910 41834
rect 68848 41806 68922 41834
rect 69860 41806 69934 41834
rect 70872 41806 70946 41834
rect 71884 41806 71958 41834
rect 72988 41806 73062 41834
rect 74000 41806 74074 41834
rect 75012 41806 75086 41834
rect 75932 41806 76098 41834
rect 77036 41806 77110 41834
rect 78048 41806 78122 41834
rect 79060 41806 79134 41834
rect 80072 41806 80146 41834
rect 81084 41806 81158 41834
rect 82096 41806 82170 41834
rect 83108 41806 83182 41834
rect 84166 41834 84194 42092
rect 85178 41834 85206 42092
rect 86190 41834 86218 42092
rect 87202 41834 87230 42092
rect 84166 41806 84240 41834
rect 65812 39234 65840 41806
rect 65800 39228 65852 39234
rect 65800 39170 65852 39176
rect 66824 38894 66852 41806
rect 67548 39704 67600 39710
rect 67548 39646 67600 39652
rect 66812 38888 66864 38894
rect 66812 38830 66864 38836
rect 66168 38004 66220 38010
rect 66168 37946 66220 37952
rect 64880 4684 64932 4690
rect 64880 4626 64932 4632
rect 64144 3868 64196 3874
rect 64144 3810 64196 3816
rect 64328 3732 64380 3738
rect 64328 3674 64380 3680
rect 64340 480 64368 3674
rect 66180 3534 66208 37946
rect 67560 3534 67588 39646
rect 67836 38146 67864 41806
rect 68848 39302 68876 41806
rect 68928 39908 68980 39914
rect 68928 39850 68980 39856
rect 68836 39296 68888 39302
rect 68836 39238 68888 39244
rect 68284 39228 68336 39234
rect 68284 39170 68336 39176
rect 67824 38140 67876 38146
rect 67824 38082 67876 38088
rect 68296 4010 68324 39170
rect 68284 4004 68336 4010
rect 68284 3946 68336 3952
rect 68940 3534 68968 39850
rect 69860 39642 69888 41806
rect 69848 39636 69900 39642
rect 69848 39578 69900 39584
rect 70308 39636 70360 39642
rect 70308 39578 70360 39584
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 66720 3528 66772 3534
rect 66720 3470 66772 3476
rect 67548 3528 67600 3534
rect 67548 3470 67600 3476
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 65536 480 65564 3470
rect 66732 480 66760 3470
rect 67928 480 67956 3470
rect 69124 480 69152 3538
rect 70320 480 70348 39578
rect 70872 38350 70900 41806
rect 71780 39296 71832 39302
rect 71780 39238 71832 39244
rect 71044 38888 71096 38894
rect 71044 38830 71096 38836
rect 70860 38344 70912 38350
rect 70860 38286 70912 38292
rect 71056 3806 71084 38830
rect 71136 38684 71188 38690
rect 71136 38626 71188 38632
rect 71044 3800 71096 3806
rect 71044 3742 71096 3748
rect 71148 3466 71176 38626
rect 71792 36582 71820 39238
rect 71884 39166 71912 41806
rect 71872 39160 71924 39166
rect 71872 39102 71924 39108
rect 72424 39160 72476 39166
rect 72424 39102 72476 39108
rect 71780 36576 71832 36582
rect 71780 36518 71832 36524
rect 72436 4078 72464 39102
rect 72988 38894 73016 41806
rect 74000 39302 74028 41806
rect 74448 39976 74500 39982
rect 74448 39918 74500 39924
rect 73988 39296 74040 39302
rect 73988 39238 74040 39244
rect 73068 39160 73120 39166
rect 73068 39102 73120 39108
rect 73080 38894 73108 39102
rect 72976 38888 73028 38894
rect 72976 38830 73028 38836
rect 73068 38888 73120 38894
rect 73068 38830 73120 38836
rect 72608 4820 72660 4826
rect 72608 4762 72660 4768
rect 72424 4072 72476 4078
rect 72424 4014 72476 4020
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 71136 3460 71188 3466
rect 71136 3402 71188 3408
rect 71516 480 71544 3810
rect 72620 480 72648 4762
rect 74460 3534 74488 39918
rect 75012 39098 75040 41806
rect 75828 40044 75880 40050
rect 75828 39986 75880 39992
rect 75184 39296 75236 39302
rect 75184 39238 75236 39244
rect 75000 39092 75052 39098
rect 75000 39034 75052 39040
rect 75196 3942 75224 39238
rect 75184 3936 75236 3942
rect 75184 3878 75236 3884
rect 75840 3534 75868 39986
rect 75932 3670 75960 41806
rect 77036 38418 77064 41806
rect 78048 38826 78076 41806
rect 78588 39160 78640 39166
rect 78588 39102 78640 39108
rect 78036 38820 78088 38826
rect 78036 38762 78088 38768
rect 77024 38412 77076 38418
rect 77024 38354 77076 38360
rect 75920 3664 75972 3670
rect 75920 3606 75972 3612
rect 78600 3534 78628 39102
rect 79060 39030 79088 41806
rect 79048 39024 79100 39030
rect 79048 38966 79100 38972
rect 80072 38962 80100 41806
rect 80060 38956 80112 38962
rect 80060 38898 80112 38904
rect 80704 38820 80756 38826
rect 80704 38762 80756 38768
rect 79968 38140 80020 38146
rect 79968 38082 80020 38088
rect 79980 6914 80008 38082
rect 79704 6886 80008 6914
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 74448 3528 74500 3534
rect 74448 3470 74500 3476
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 77392 3528 77444 3534
rect 77392 3470 77444 3476
rect 78588 3528 78640 3534
rect 78588 3470 78640 3476
rect 73816 480 73844 3470
rect 75012 480 75040 3470
rect 76196 3392 76248 3398
rect 76196 3334 76248 3340
rect 76208 480 76236 3334
rect 77404 480 77432 3470
rect 78588 3188 78640 3194
rect 78588 3130 78640 3136
rect 78600 480 78628 3130
rect 79704 480 79732 6886
rect 80716 3874 80744 38762
rect 81084 38758 81112 41806
rect 82096 39302 82124 41806
rect 82084 39296 82136 39302
rect 82084 39238 82136 39244
rect 81348 39228 81400 39234
rect 81348 39170 81400 39176
rect 81072 38752 81124 38758
rect 81072 38694 81124 38700
rect 80704 3868 80756 3874
rect 80704 3810 80756 3816
rect 81360 3398 81388 39170
rect 82084 39092 82136 39098
rect 82084 39034 82136 39040
rect 82096 6914 82124 39034
rect 83108 38214 83136 41806
rect 84212 39370 84240 41806
rect 85132 41806 85206 41834
rect 86144 41806 86218 41834
rect 87156 41806 87230 41834
rect 88306 41834 88334 42092
rect 89318 41834 89346 42092
rect 90330 41834 90358 42092
rect 91342 41834 91370 42092
rect 92354 41834 92382 42092
rect 93366 41834 93394 42092
rect 94378 41834 94406 42092
rect 95390 41834 95418 42092
rect 96402 41834 96430 42092
rect 97414 41834 97442 42092
rect 98426 41834 98454 42092
rect 99438 41834 99466 42092
rect 100450 41834 100478 42092
rect 101462 41834 101490 42092
rect 102474 41834 102502 42092
rect 103578 41834 103606 42092
rect 104590 41834 104618 42092
rect 105602 41834 105630 42092
rect 106614 41834 106642 42092
rect 88306 41806 88380 41834
rect 84200 39364 84252 39370
rect 84200 39306 84252 39312
rect 84844 39160 84896 39166
rect 84844 39102 84896 39108
rect 83096 38208 83148 38214
rect 83096 38150 83148 38156
rect 84108 38208 84160 38214
rect 84108 38150 84160 38156
rect 82004 6886 82124 6914
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 80900 480 80928 3334
rect 82004 3194 82032 6886
rect 82084 4072 82136 4078
rect 82084 4014 82136 4020
rect 81992 3188 82044 3194
rect 81992 3130 82044 3136
rect 82096 480 82124 4014
rect 84120 3398 84148 38150
rect 84856 4078 84884 39102
rect 85132 39030 85160 41806
rect 85488 39364 85540 39370
rect 85488 39306 85540 39312
rect 85120 39024 85172 39030
rect 85120 38966 85172 38972
rect 84844 4072 84896 4078
rect 84844 4014 84896 4020
rect 83280 3392 83332 3398
rect 83280 3334 83332 3340
rect 84108 3392 84160 3398
rect 84108 3334 84160 3340
rect 83292 480 83320 3334
rect 85500 2922 85528 39306
rect 86144 37942 86172 41806
rect 87156 39574 87184 41806
rect 87144 39568 87196 39574
rect 87144 39510 87196 39516
rect 88248 39568 88300 39574
rect 88248 39510 88300 39516
rect 86132 37936 86184 37942
rect 86132 37878 86184 37884
rect 86868 37936 86920 37942
rect 86868 37878 86920 37884
rect 85672 3460 85724 3466
rect 85672 3402 85724 3408
rect 84476 2916 84528 2922
rect 84476 2858 84528 2864
rect 85488 2916 85540 2922
rect 85488 2858 85540 2864
rect 84488 480 84516 2858
rect 85684 480 85712 3402
rect 86880 480 86908 37878
rect 88260 6914 88288 39510
rect 88352 38690 88380 41806
rect 89272 41806 89346 41834
rect 90284 41806 90358 41834
rect 91296 41806 91370 41834
rect 92308 41806 92382 41834
rect 93320 41806 93394 41834
rect 94332 41806 94406 41834
rect 95344 41806 95418 41834
rect 96356 41806 96430 41834
rect 97368 41806 97442 41834
rect 98380 41806 98454 41834
rect 99392 41806 99466 41834
rect 100404 41806 100478 41834
rect 100772 41806 101490 41834
rect 102428 41806 102502 41834
rect 103532 41806 103606 41834
rect 103716 41806 104618 41834
rect 105556 41806 105630 41834
rect 106568 41806 106642 41834
rect 107626 41834 107654 42092
rect 108638 41834 108666 42092
rect 109650 41834 109678 42092
rect 110662 41834 110690 42092
rect 111674 41834 111702 42092
rect 112686 41834 112714 42092
rect 113698 41834 113726 42092
rect 114710 41834 114738 42092
rect 115722 41834 115750 42092
rect 116734 41834 116762 42092
rect 117746 41834 117774 42092
rect 118850 41834 118878 42092
rect 119862 41834 119890 42092
rect 120874 41834 120902 42092
rect 121886 41834 121914 42092
rect 107626 41806 107700 41834
rect 88984 38956 89036 38962
rect 88984 38898 89036 38904
rect 88340 38684 88392 38690
rect 88340 38626 88392 38632
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 88996 3466 89024 38898
rect 89076 38752 89128 38758
rect 89076 38694 89128 38700
rect 89088 3738 89116 38694
rect 89272 38282 89300 41806
rect 90284 39506 90312 41806
rect 90272 39500 90324 39506
rect 90272 39442 90324 39448
rect 91296 39438 91324 41806
rect 91284 39432 91336 39438
rect 91284 39374 91336 39380
rect 91744 39024 91796 39030
rect 91744 38966 91796 38972
rect 89260 38276 89312 38282
rect 89260 38218 89312 38224
rect 91008 38276 91060 38282
rect 91008 38218 91060 38224
rect 89076 3732 89128 3738
rect 89076 3674 89128 3680
rect 91020 3466 91048 38218
rect 88984 3460 89036 3466
rect 88984 3402 89036 3408
rect 90364 3460 90416 3466
rect 90364 3402 90416 3408
rect 91008 3460 91060 3466
rect 91008 3402 91060 3408
rect 91560 3460 91612 3466
rect 91560 3402 91612 3408
rect 89168 3392 89220 3398
rect 89168 3334 89220 3340
rect 89180 480 89208 3334
rect 90376 480 90404 3402
rect 91572 480 91600 3402
rect 91756 3398 91784 38966
rect 92308 38078 92336 41806
rect 93320 39846 93348 41806
rect 93308 39840 93360 39846
rect 93308 39782 93360 39788
rect 92388 39500 92440 39506
rect 92388 39442 92440 39448
rect 92296 38072 92348 38078
rect 92296 38014 92348 38020
rect 92400 3466 92428 39442
rect 94332 38894 94360 41806
rect 95148 39840 95200 39846
rect 95148 39782 95200 39788
rect 94320 38888 94372 38894
rect 94320 38830 94372 38836
rect 93124 37324 93176 37330
rect 93124 37266 93176 37272
rect 92756 4004 92808 4010
rect 92756 3946 92808 3952
rect 92388 3460 92440 3466
rect 92388 3402 92440 3408
rect 91744 3392 91796 3398
rect 91744 3334 91796 3340
rect 92768 480 92796 3946
rect 93136 3330 93164 37266
rect 93952 3392 94004 3398
rect 93952 3334 94004 3340
rect 93124 3324 93176 3330
rect 93124 3266 93176 3272
rect 93964 480 93992 3334
rect 95160 480 95188 39782
rect 95344 37330 95372 41806
rect 96356 39778 96384 41806
rect 96344 39772 96396 39778
rect 96344 39714 96396 39720
rect 95884 38888 95936 38894
rect 95884 38830 95936 38836
rect 95332 37324 95384 37330
rect 95332 37266 95384 37272
rect 95896 4010 95924 38830
rect 97368 38758 97396 41806
rect 97356 38752 97408 38758
rect 97356 38694 97408 38700
rect 98380 38010 98408 41806
rect 99392 39710 99420 41806
rect 100404 39914 100432 41806
rect 100392 39908 100444 39914
rect 100392 39850 100444 39856
rect 99380 39704 99432 39710
rect 99380 39646 99432 39652
rect 100668 39704 100720 39710
rect 100668 39646 100720 39652
rect 99288 39432 99340 39438
rect 99288 39374 99340 39380
rect 98368 38004 98420 38010
rect 98368 37946 98420 37952
rect 97908 36576 97960 36582
rect 97908 36518 97960 36524
rect 95884 4004 95936 4010
rect 95884 3946 95936 3952
rect 96252 3664 96304 3670
rect 96252 3606 96304 3612
rect 96264 480 96292 3606
rect 97920 3466 97948 36518
rect 99300 3466 99328 39374
rect 100680 3466 100708 39646
rect 100772 3602 100800 41806
rect 102428 39642 102456 41806
rect 103428 39908 103480 39914
rect 103428 39850 103480 39856
rect 102416 39636 102468 39642
rect 102416 39578 102468 39584
rect 103336 39636 103388 39642
rect 103336 39578 103388 39584
rect 102048 26920 102100 26926
rect 102048 26862 102100 26868
rect 100760 3596 100812 3602
rect 100760 3538 100812 3544
rect 102060 3466 102088 26862
rect 97448 3460 97500 3466
rect 97448 3402 97500 3408
rect 97908 3460 97960 3466
rect 97908 3402 97960 3408
rect 98644 3460 98696 3466
rect 98644 3402 98696 3408
rect 99288 3460 99340 3466
rect 99288 3402 99340 3408
rect 99840 3460 99892 3466
rect 99840 3402 99892 3408
rect 100668 3460 100720 3466
rect 100668 3402 100720 3408
rect 101036 3460 101088 3466
rect 101036 3402 101088 3408
rect 102048 3460 102100 3466
rect 102048 3402 102100 3408
rect 97460 480 97488 3402
rect 98656 480 98684 3402
rect 99852 480 99880 3402
rect 101048 480 101076 3402
rect 102232 3120 102284 3126
rect 102232 3062 102284 3068
rect 102244 480 102272 3062
rect 103348 480 103376 39578
rect 103440 3126 103468 39850
rect 103532 38826 103560 41806
rect 103520 38820 103572 38826
rect 103520 38762 103572 38768
rect 103716 4826 103744 41806
rect 105556 39982 105584 41806
rect 106568 40050 106596 41806
rect 106556 40044 106608 40050
rect 106556 39986 106608 39992
rect 105544 39976 105596 39982
rect 105544 39918 105596 39924
rect 107568 39976 107620 39982
rect 107568 39918 107620 39924
rect 106188 39772 106240 39778
rect 106188 39714 106240 39720
rect 104808 36644 104860 36650
rect 104808 36586 104860 36592
rect 104820 6914 104848 36586
rect 104544 6886 104848 6914
rect 103704 4820 103756 4826
rect 103704 4762 103756 4768
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 104544 480 104572 6886
rect 106200 3534 106228 39714
rect 106924 38752 106976 38758
rect 106924 38694 106976 38700
rect 106936 3670 106964 38694
rect 106924 3664 106976 3670
rect 106924 3606 106976 3612
rect 107580 3534 107608 39918
rect 107672 3602 107700 41806
rect 108592 41806 108666 41834
rect 109604 41806 109678 41834
rect 110616 41806 110690 41834
rect 111628 41806 111702 41834
rect 112640 41806 112714 41834
rect 113652 41806 113726 41834
rect 114664 41806 114738 41834
rect 115676 41806 115750 41834
rect 116688 41806 116762 41834
rect 117700 41806 117774 41834
rect 118804 41806 118878 41834
rect 119816 41806 119890 41834
rect 120828 41806 120902 41834
rect 121840 41806 121914 41834
rect 122898 41834 122926 42092
rect 123910 41834 123938 42092
rect 124922 41834 124950 42092
rect 125934 41834 125962 42092
rect 122898 41806 122972 41834
rect 108592 39234 108620 41806
rect 108580 39228 108632 39234
rect 108580 39170 108632 39176
rect 109604 39098 109632 41806
rect 110328 40044 110380 40050
rect 110328 39986 110380 39992
rect 109592 39092 109644 39098
rect 109592 39034 109644 39040
rect 108120 3664 108172 3670
rect 108120 3606 108172 3612
rect 107660 3596 107712 3602
rect 107660 3538 107712 3544
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 105740 480 105768 3470
rect 106936 480 106964 3470
rect 108132 480 108160 3606
rect 110340 3534 110368 39986
rect 110616 38146 110644 41806
rect 111628 39302 111656 41806
rect 111616 39296 111668 39302
rect 111616 39238 111668 39244
rect 112640 39166 112668 41806
rect 113088 39296 113140 39302
rect 113088 39238 113140 39244
rect 112628 39160 112680 39166
rect 112628 39102 112680 39108
rect 111708 39092 111760 39098
rect 111708 39034 111760 39040
rect 110604 38140 110656 38146
rect 110604 38082 110656 38088
rect 111616 3596 111668 3602
rect 111616 3538 111668 3544
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 110328 3528 110380 3534
rect 110328 3470 110380 3476
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 109328 480 109356 3470
rect 110524 480 110552 3470
rect 111628 480 111656 3538
rect 111720 3534 111748 39034
rect 113100 6914 113128 39238
rect 113652 38214 113680 41806
rect 114664 39370 114692 41806
rect 114652 39364 114704 39370
rect 114652 39306 114704 39312
rect 114468 39228 114520 39234
rect 114468 39170 114520 39176
rect 113640 38208 113692 38214
rect 113640 38150 113692 38156
rect 112824 6886 113128 6914
rect 111708 3528 111760 3534
rect 111708 3470 111760 3476
rect 112824 480 112852 6886
rect 114480 3398 114508 39170
rect 115676 38962 115704 41806
rect 115848 39160 115900 39166
rect 115848 39102 115900 39108
rect 115664 38956 115716 38962
rect 115664 38898 115716 38904
rect 115860 3398 115888 39102
rect 116688 37942 116716 41806
rect 117700 39574 117728 41806
rect 117688 39568 117740 39574
rect 117688 39510 117740 39516
rect 117228 39364 117280 39370
rect 117228 39306 117280 39312
rect 116676 37936 116728 37942
rect 116676 37878 116728 37884
rect 117240 3398 117268 39306
rect 118804 39030 118832 41806
rect 118792 39024 118844 39030
rect 118792 38966 118844 38972
rect 118608 38956 118660 38962
rect 118608 38898 118660 38904
rect 118620 3398 118648 38898
rect 119816 38282 119844 41806
rect 119988 39568 120040 39574
rect 119988 39510 120040 39516
rect 119896 39024 119948 39030
rect 119896 38966 119948 38972
rect 119804 38276 119856 38282
rect 119804 38218 119856 38224
rect 119908 16574 119936 38966
rect 119816 16546 119936 16574
rect 119816 3398 119844 16546
rect 120000 6914 120028 39510
rect 120828 39506 120856 41806
rect 120816 39500 120868 39506
rect 120816 39442 120868 39448
rect 121368 39500 121420 39506
rect 121368 39442 121420 39448
rect 121380 6914 121408 39442
rect 121840 38894 121868 41806
rect 121828 38888 121880 38894
rect 121828 38830 121880 38836
rect 122748 38820 122800 38826
rect 122748 38762 122800 38768
rect 119908 6886 120028 6914
rect 121104 6886 121408 6914
rect 114008 3392 114060 3398
rect 114008 3334 114060 3340
rect 114468 3392 114520 3398
rect 114468 3334 114520 3340
rect 115204 3392 115256 3398
rect 115204 3334 115256 3340
rect 115848 3392 115900 3398
rect 115848 3334 115900 3340
rect 116400 3392 116452 3398
rect 116400 3334 116452 3340
rect 117228 3392 117280 3398
rect 117228 3334 117280 3340
rect 117596 3392 117648 3398
rect 117596 3334 117648 3340
rect 118608 3392 118660 3398
rect 118608 3334 118660 3340
rect 118792 3392 118844 3398
rect 118792 3334 118844 3340
rect 119804 3392 119856 3398
rect 119804 3334 119856 3340
rect 114020 480 114048 3334
rect 115216 480 115244 3334
rect 116412 480 116440 3334
rect 117608 480 117636 3334
rect 118804 480 118832 3334
rect 119908 480 119936 6886
rect 121104 480 121132 6886
rect 122760 3398 122788 38762
rect 122944 3466 122972 41806
rect 123864 41806 123938 41834
rect 124876 41806 124950 41834
rect 125888 41806 125962 41834
rect 126946 41834 126974 42092
rect 127958 41834 127986 42092
rect 128970 41834 128998 42092
rect 129982 41834 130010 42092
rect 130994 41834 131022 42092
rect 132006 41834 132034 42092
rect 133018 41834 133046 42092
rect 126946 41806 127020 41834
rect 123864 39846 123892 41806
rect 123852 39840 123904 39846
rect 123852 39782 123904 39788
rect 124128 39840 124180 39846
rect 124128 39782 124180 39788
rect 124140 3534 124168 39782
rect 124876 38758 124904 41806
rect 125508 38888 125560 38894
rect 125508 38830 125560 38836
rect 124864 38752 124916 38758
rect 124864 38694 124916 38700
rect 125520 3534 125548 38830
rect 125888 36582 125916 41806
rect 126992 39438 127020 41806
rect 127912 41806 127986 41834
rect 128372 41806 128998 41834
rect 129936 41806 130010 41834
rect 130948 41806 131022 41834
rect 131960 41806 132034 41834
rect 132972 41806 133046 41834
rect 133972 41880 134024 41886
rect 134122 41834 134150 42092
rect 135134 41886 135162 42092
rect 133972 41822 134024 41828
rect 127912 39710 127940 41806
rect 127900 39704 127952 39710
rect 127900 39646 127952 39652
rect 126980 39432 127032 39438
rect 126980 39374 127032 39380
rect 126888 37936 126940 37942
rect 126888 37878 126940 37884
rect 125876 36576 125928 36582
rect 125876 36518 125928 36524
rect 126900 3534 126928 37878
rect 128372 26926 128400 41806
rect 129936 39914 129964 41806
rect 129924 39908 129976 39914
rect 129924 39850 129976 39856
rect 130948 39642 130976 41806
rect 130936 39636 130988 39642
rect 130936 39578 130988 39584
rect 131960 38758 131988 41806
rect 132972 39778 133000 41806
rect 132960 39772 133012 39778
rect 132960 39714 133012 39720
rect 132408 39432 132460 39438
rect 132408 39374 132460 39380
rect 129740 38752 129792 38758
rect 129740 38694 129792 38700
rect 131948 38752 132000 38758
rect 131948 38694 132000 38700
rect 129648 38004 129700 38010
rect 129648 37946 129700 37952
rect 128360 26920 128412 26926
rect 128360 26862 128412 26868
rect 129464 8968 129516 8974
rect 129464 8910 129516 8916
rect 128360 4548 128412 4554
rect 128360 4490 128412 4496
rect 128372 3670 128400 4490
rect 128360 3664 128412 3670
rect 128360 3606 128412 3612
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 128176 3528 128228 3534
rect 128176 3470 128228 3476
rect 122932 3460 122984 3466
rect 122932 3402 122984 3408
rect 122288 3392 122340 3398
rect 122288 3334 122340 3340
rect 122748 3392 122800 3398
rect 122748 3334 122800 3340
rect 122300 480 122328 3334
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 126980 3120 127032 3126
rect 126980 3062 127032 3068
rect 126992 480 127020 3062
rect 128188 480 128216 3470
rect 129476 3126 129504 8910
rect 129660 6914 129688 37946
rect 129752 36650 129780 38694
rect 130384 38140 130436 38146
rect 130384 38082 130436 38088
rect 129740 36644 129792 36650
rect 129740 36586 129792 36592
rect 129568 6886 129688 6914
rect 129464 3120 129516 3126
rect 129464 3062 129516 3068
rect 129568 2938 129596 6886
rect 130396 3534 130424 38082
rect 131028 36576 131080 36582
rect 131028 36518 131080 36524
rect 131040 3534 131068 36518
rect 132420 3534 132448 39374
rect 133788 38072 133840 38078
rect 133788 38014 133840 38020
rect 133800 3534 133828 38014
rect 133984 4554 134012 41822
rect 134076 41806 134150 41834
rect 135122 41880 135174 41886
rect 136146 41834 136174 42092
rect 137158 41834 137186 42092
rect 138170 41834 138198 42092
rect 139182 41834 139210 42092
rect 140194 41834 140222 42092
rect 141206 41834 141234 42092
rect 142218 41834 142246 42092
rect 143230 41834 143258 42092
rect 144242 41834 144270 42092
rect 145254 41834 145282 42092
rect 135122 41822 135174 41828
rect 136100 41806 136174 41834
rect 137112 41806 137186 41834
rect 138124 41806 138198 41834
rect 139136 41806 139210 41834
rect 140148 41806 140222 41834
rect 141160 41806 141234 41834
rect 142172 41806 142246 41834
rect 143184 41806 143258 41834
rect 144196 41806 144270 41834
rect 145208 41806 145282 41834
rect 146266 41834 146294 42092
rect 147278 41834 147306 42092
rect 148290 41834 148318 42092
rect 149394 41834 149422 42092
rect 146266 41806 146340 41834
rect 134076 39982 134104 41806
rect 136100 40050 136128 41806
rect 136088 40044 136140 40050
rect 136088 39986 136140 39992
rect 136548 40044 136600 40050
rect 136548 39986 136600 39992
rect 134064 39976 134116 39982
rect 134064 39918 134116 39924
rect 135168 39704 135220 39710
rect 135168 39646 135220 39652
rect 133972 4548 134024 4554
rect 133972 4490 134024 4496
rect 135180 3534 135208 39646
rect 136560 3534 136588 39986
rect 137112 39098 137140 41806
rect 137928 39636 137980 39642
rect 137928 39578 137980 39584
rect 137100 39092 137152 39098
rect 137100 39034 137152 39040
rect 137284 39092 137336 39098
rect 137284 39034 137336 39040
rect 137296 3602 137324 39034
rect 137940 6914 137968 39578
rect 138124 39098 138152 41806
rect 139136 39302 139164 41806
rect 139308 39772 139360 39778
rect 139308 39714 139360 39720
rect 139124 39296 139176 39302
rect 139124 39238 139176 39244
rect 138112 39092 138164 39098
rect 138112 39034 138164 39040
rect 137664 6886 137968 6914
rect 137284 3596 137336 3602
rect 137284 3538 137336 3544
rect 130384 3528 130436 3534
rect 130384 3470 130436 3476
rect 130568 3528 130620 3534
rect 130568 3470 130620 3476
rect 131028 3528 131080 3534
rect 131028 3470 131080 3476
rect 131764 3528 131816 3534
rect 131764 3470 131816 3476
rect 132408 3528 132460 3534
rect 132408 3470 132460 3476
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 134156 3528 134208 3534
rect 134156 3470 134208 3476
rect 135168 3528 135220 3534
rect 135168 3470 135220 3476
rect 135260 3528 135312 3534
rect 135260 3470 135312 3476
rect 136548 3528 136600 3534
rect 136548 3470 136600 3476
rect 129384 2910 129596 2938
rect 129384 480 129412 2910
rect 130580 480 130608 3470
rect 131776 480 131804 3470
rect 132972 480 133000 3470
rect 134168 480 134196 3470
rect 135272 480 135300 3470
rect 136456 2848 136508 2854
rect 136456 2790 136508 2796
rect 136468 480 136496 2790
rect 137664 480 137692 6886
rect 139320 3534 139348 39714
rect 140148 39234 140176 41806
rect 140136 39228 140188 39234
rect 140136 39170 140188 39176
rect 140688 39228 140740 39234
rect 140688 39170 140740 39176
rect 139400 4820 139452 4826
rect 139400 4762 139452 4768
rect 138848 3528 138900 3534
rect 138848 3470 138900 3476
rect 139308 3528 139360 3534
rect 139308 3470 139360 3476
rect 138860 480 138888 3470
rect 139412 2854 139440 4762
rect 140700 3534 140728 39170
rect 141160 39166 141188 41806
rect 142068 39908 142120 39914
rect 142068 39850 142120 39856
rect 141148 39160 141200 39166
rect 141148 39102 141200 39108
rect 142080 3534 142108 39850
rect 142172 39370 142200 41806
rect 142160 39364 142212 39370
rect 142160 39306 142212 39312
rect 143184 38962 143212 41806
rect 143448 39296 143500 39302
rect 143448 39238 143500 39244
rect 143172 38956 143224 38962
rect 143172 38898 143224 38904
rect 143460 3534 143488 39238
rect 144196 39030 144224 41806
rect 144828 39976 144880 39982
rect 144828 39918 144880 39924
rect 144736 39364 144788 39370
rect 144736 39306 144788 39312
rect 144184 39024 144236 39030
rect 144184 38966 144236 38972
rect 144748 16574 144776 39306
rect 144656 16546 144776 16574
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 140688 3528 140740 3534
rect 140688 3470 140740 3476
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 142068 3528 142120 3534
rect 142068 3470 142120 3476
rect 142436 3528 142488 3534
rect 142436 3470 142488 3476
rect 143448 3528 143500 3534
rect 143448 3470 143500 3476
rect 139400 2848 139452 2854
rect 139400 2790 139452 2796
rect 140056 480 140084 3470
rect 141252 480 141280 3470
rect 142448 480 142476 3470
rect 144656 3058 144684 16546
rect 144840 6914 144868 39918
rect 145208 39574 145236 41806
rect 145196 39568 145248 39574
rect 145196 39510 145248 39516
rect 146312 39506 146340 41806
rect 147232 41806 147306 41834
rect 148244 41806 148318 41834
rect 149348 41806 149422 41834
rect 150406 41834 150434 42092
rect 151418 41834 151446 42092
rect 152430 41834 152458 42092
rect 153442 41834 153470 42092
rect 154454 41834 154482 42092
rect 155466 41834 155494 42092
rect 156478 41834 156506 42092
rect 157490 41834 157518 42092
rect 158502 41834 158530 42092
rect 159514 41834 159542 42092
rect 160526 41834 160554 42092
rect 161538 41834 161566 42092
rect 162550 41834 162578 42092
rect 163562 41834 163590 42092
rect 164666 41834 164694 42092
rect 165678 41834 165706 42092
rect 166690 41834 166718 42092
rect 167702 41834 167730 42092
rect 168714 41834 168742 42092
rect 150406 41806 150480 41834
rect 146944 39568 146996 39574
rect 146944 39510 146996 39516
rect 146300 39500 146352 39506
rect 146300 39442 146352 39448
rect 146208 38752 146260 38758
rect 146208 38694 146260 38700
rect 146220 6914 146248 38694
rect 146956 36582 146984 39510
rect 147232 38826 147260 41806
rect 148244 39846 148272 41806
rect 148232 39840 148284 39846
rect 148232 39782 148284 39788
rect 148968 39500 149020 39506
rect 148968 39442 149020 39448
rect 147588 39160 147640 39166
rect 147588 39102 147640 39108
rect 147220 38820 147272 38826
rect 147220 38762 147272 38768
rect 146944 36576 146996 36582
rect 146944 36518 146996 36524
rect 144748 6886 144868 6914
rect 145944 6886 146248 6914
rect 143540 3052 143592 3058
rect 143540 2994 143592 3000
rect 144644 3052 144696 3058
rect 144644 2994 144696 3000
rect 143552 480 143580 2994
rect 144748 480 144776 6886
rect 145944 480 145972 6886
rect 147600 3534 147628 39102
rect 148980 3534 149008 39442
rect 149348 38894 149376 41806
rect 150348 39024 150400 39030
rect 150348 38966 150400 38972
rect 149336 38888 149388 38894
rect 149336 38830 149388 38836
rect 150360 3534 150388 38966
rect 150452 37942 150480 41806
rect 150636 41806 151446 41834
rect 152384 41806 152458 41834
rect 153396 41806 153470 41834
rect 154408 41806 154482 41834
rect 155420 41806 155494 41834
rect 156432 41806 156506 41834
rect 157444 41806 157518 41834
rect 158456 41806 158530 41834
rect 158732 41806 159542 41834
rect 160480 41806 160554 41834
rect 161492 41806 161566 41834
rect 162504 41806 162578 41834
rect 163516 41806 163590 41834
rect 164620 41806 164694 41834
rect 165632 41806 165706 41834
rect 166644 41806 166718 41834
rect 167656 41806 167730 41834
rect 168668 41806 168742 41834
rect 169726 41834 169754 42092
rect 170738 41834 170766 42092
rect 171750 41834 171778 42092
rect 172762 41834 172790 42092
rect 173774 41834 173802 42092
rect 174786 41834 174814 42092
rect 175798 41834 175826 42092
rect 176810 41834 176838 42092
rect 177822 41834 177850 42092
rect 178834 41834 178862 42092
rect 179938 41834 179966 42092
rect 180950 41834 180978 42092
rect 181962 41834 181990 42092
rect 182974 41834 183002 42092
rect 183986 41834 184014 42092
rect 184998 41834 185026 42092
rect 186010 41834 186038 42092
rect 187022 41834 187050 42092
rect 188034 41834 188062 42092
rect 169726 41806 169800 41834
rect 150440 37936 150492 37942
rect 150440 37878 150492 37884
rect 150636 8974 150664 41806
rect 151728 38888 151780 38894
rect 151728 38830 151780 38836
rect 150624 8968 150676 8974
rect 150624 8910 150676 8916
rect 151740 3534 151768 38830
rect 152384 38146 152412 41806
rect 153016 39840 153068 39846
rect 153016 39782 153068 39788
rect 152372 38140 152424 38146
rect 152372 38082 152424 38088
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 150348 3528 150400 3534
rect 150348 3470 150400 3476
rect 150624 3528 150676 3534
rect 150624 3470 150676 3476
rect 151728 3528 151780 3534
rect 151728 3470 151780 3476
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 147140 480 147168 3470
rect 148336 480 148364 3470
rect 149532 480 149560 3470
rect 150636 480 150664 3470
rect 151832 480 151860 3470
rect 153028 480 153056 39782
rect 153108 39092 153160 39098
rect 153108 39034 153160 39040
rect 153120 3534 153148 39034
rect 153396 38010 153424 41806
rect 154408 39574 154436 41806
rect 154396 39568 154448 39574
rect 154396 39510 154448 39516
rect 155420 39438 155448 41806
rect 155408 39432 155460 39438
rect 155408 39374 155460 39380
rect 155868 39432 155920 39438
rect 155868 39374 155920 39380
rect 154488 38956 154540 38962
rect 154488 38898 154540 38904
rect 153384 38004 153436 38010
rect 153384 37946 153436 37952
rect 154500 6914 154528 38898
rect 154224 6886 154528 6914
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 154224 480 154252 6886
rect 155880 3534 155908 39374
rect 156432 38078 156460 41806
rect 157444 39710 157472 41806
rect 158456 40050 158484 41806
rect 158444 40044 158496 40050
rect 158444 39986 158496 39992
rect 158628 40044 158680 40050
rect 158628 39986 158680 39992
rect 157432 39704 157484 39710
rect 157432 39646 157484 39652
rect 157248 38820 157300 38826
rect 157248 38762 157300 38768
rect 156420 38072 156472 38078
rect 156420 38014 156472 38020
rect 157260 3534 157288 38762
rect 158640 3534 158668 39986
rect 158732 4826 158760 41806
rect 160008 39704 160060 39710
rect 160008 39646 160060 39652
rect 158720 4820 158772 4826
rect 158720 4762 158772 4768
rect 160020 3534 160048 39646
rect 160480 39642 160508 41806
rect 161492 39778 161520 41806
rect 161480 39772 161532 39778
rect 161480 39714 161532 39720
rect 160468 39636 160520 39642
rect 160468 39578 160520 39584
rect 162504 39234 162532 41806
rect 163516 39914 163544 41806
rect 163504 39908 163556 39914
rect 163504 39850 163556 39856
rect 162768 39772 162820 39778
rect 162768 39714 162820 39720
rect 162492 39228 162544 39234
rect 162492 39170 162544 39176
rect 161388 38752 161440 38758
rect 161388 38694 161440 38700
rect 161400 3534 161428 38694
rect 162780 6914 162808 39714
rect 164148 39636 164200 39642
rect 164148 39578 164200 39584
rect 162504 6886 162808 6914
rect 155408 3528 155460 3534
rect 155408 3470 155460 3476
rect 155868 3528 155920 3534
rect 155868 3470 155920 3476
rect 156604 3528 156656 3534
rect 156604 3470 156656 3476
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 157800 3528 157852 3534
rect 157800 3470 157852 3476
rect 158628 3528 158680 3534
rect 158628 3470 158680 3476
rect 158904 3528 158956 3534
rect 158904 3470 158956 3476
rect 160008 3528 160060 3534
rect 160008 3470 160060 3476
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 161388 3528 161440 3534
rect 161388 3470 161440 3476
rect 155420 480 155448 3470
rect 156616 480 156644 3470
rect 157812 480 157840 3470
rect 158916 480 158944 3470
rect 160112 480 160140 3470
rect 161296 3460 161348 3466
rect 161296 3402 161348 3408
rect 161308 480 161336 3402
rect 162504 480 162532 6886
rect 164160 3534 164188 39578
rect 164620 39302 164648 41806
rect 165528 39908 165580 39914
rect 165528 39850 165580 39856
rect 164608 39296 164660 39302
rect 164608 39238 164660 39244
rect 163688 3528 163740 3534
rect 163688 3470 163740 3476
rect 164148 3528 164200 3534
rect 164148 3470 164200 3476
rect 163700 480 163728 3470
rect 165540 3058 165568 39850
rect 165632 39370 165660 41806
rect 166644 39982 166672 41806
rect 166632 39976 166684 39982
rect 166632 39918 166684 39924
rect 167656 39574 167684 41806
rect 167644 39568 167696 39574
rect 167644 39510 167696 39516
rect 165620 39364 165672 39370
rect 165620 39306 165672 39312
rect 166908 39364 166960 39370
rect 166908 39306 166960 39312
rect 166920 3534 166948 39306
rect 168288 39228 168340 39234
rect 168288 39170 168340 39176
rect 168300 3534 168328 39170
rect 168668 39166 168696 41806
rect 169576 39976 169628 39982
rect 169576 39918 169628 39924
rect 168656 39160 168708 39166
rect 168656 39102 168708 39108
rect 169588 16574 169616 39918
rect 169668 39568 169720 39574
rect 169668 39510 169720 39516
rect 169496 16546 169616 16574
rect 169496 3534 169524 16546
rect 169680 6914 169708 39510
rect 169772 39506 169800 41806
rect 170692 41806 170766 41834
rect 171704 41806 171778 41834
rect 172716 41806 172790 41834
rect 173728 41806 173802 41834
rect 174740 41806 174814 41834
rect 175752 41806 175826 41834
rect 176764 41806 176838 41834
rect 177776 41806 177850 41834
rect 178788 41806 178862 41834
rect 179892 41806 179966 41834
rect 180904 41806 180978 41834
rect 181916 41806 181990 41834
rect 182928 41806 183002 41834
rect 183940 41806 184014 41834
rect 184952 41806 185026 41834
rect 185964 41806 186038 41834
rect 186976 41806 187050 41834
rect 187988 41806 188062 41834
rect 189046 41834 189074 42092
rect 190058 41834 190086 42092
rect 191070 41834 191098 42092
rect 192082 41834 192110 42092
rect 193094 41834 193122 42092
rect 194106 41834 194134 42092
rect 195210 41834 195238 42092
rect 196222 41834 196250 42092
rect 197234 41834 197262 42092
rect 198246 41834 198274 42092
rect 199258 41834 199286 42092
rect 200270 41834 200298 42092
rect 201282 41834 201310 42092
rect 202294 41834 202322 42092
rect 203306 41834 203334 42092
rect 204318 41834 204346 42092
rect 205330 41834 205358 42092
rect 206342 41834 206370 42092
rect 207354 41834 207382 42092
rect 189046 41806 189120 41834
rect 169760 39500 169812 39506
rect 169760 39442 169812 39448
rect 170692 39030 170720 41806
rect 171048 39500 171100 39506
rect 171048 39442 171100 39448
rect 170680 39024 170732 39030
rect 170680 38966 170732 38972
rect 171060 6914 171088 39442
rect 171704 38894 171732 41806
rect 172428 39296 172480 39302
rect 172428 39238 172480 39244
rect 171692 38888 171744 38894
rect 171692 38830 171744 38836
rect 169588 6886 169708 6914
rect 170784 6886 171088 6914
rect 166080 3528 166132 3534
rect 166080 3470 166132 3476
rect 166908 3528 166960 3534
rect 166908 3470 166960 3476
rect 167184 3528 167236 3534
rect 167184 3470 167236 3476
rect 168288 3528 168340 3534
rect 168288 3470 168340 3476
rect 168380 3528 168432 3534
rect 168380 3470 168432 3476
rect 169484 3528 169536 3534
rect 169484 3470 169536 3476
rect 164884 3052 164936 3058
rect 164884 2994 164936 3000
rect 165528 3052 165580 3058
rect 165528 2994 165580 3000
rect 164896 480 164924 2994
rect 166092 480 166120 3470
rect 167196 480 167224 3470
rect 168392 480 168420 3470
rect 169588 480 169616 6886
rect 170784 480 170812 6886
rect 172440 3534 172468 39238
rect 172716 39098 172744 41806
rect 173728 39846 173756 41806
rect 173716 39840 173768 39846
rect 173716 39782 173768 39788
rect 173808 39840 173860 39846
rect 173808 39782 173860 39788
rect 172704 39092 172756 39098
rect 172704 39034 172756 39040
rect 173820 3534 173848 39782
rect 174740 38962 174768 41806
rect 175752 39438 175780 41806
rect 175740 39432 175792 39438
rect 175740 39374 175792 39380
rect 175188 39160 175240 39166
rect 175188 39102 175240 39108
rect 174728 38956 174780 38962
rect 174728 38898 174780 38904
rect 175200 3534 175228 39102
rect 176568 39024 176620 39030
rect 176568 38966 176620 38972
rect 176580 3534 176608 38966
rect 176764 38826 176792 41806
rect 177776 40050 177804 41806
rect 177764 40044 177816 40050
rect 177764 39986 177816 39992
rect 177948 40044 178000 40050
rect 177948 39986 178000 39992
rect 177856 39092 177908 39098
rect 177856 39034 177908 39040
rect 176752 38820 176804 38826
rect 176752 38762 176804 38768
rect 177868 16574 177896 39034
rect 177776 16546 177896 16574
rect 177776 3534 177804 16546
rect 177960 6914 177988 39986
rect 178788 39710 178816 41806
rect 178776 39704 178828 39710
rect 178776 39646 178828 39652
rect 179328 39432 179380 39438
rect 179328 39374 179380 39380
rect 179340 6914 179368 39374
rect 179892 38758 179920 41806
rect 180904 40050 180932 41806
rect 180064 40044 180116 40050
rect 180064 39986 180116 39992
rect 180892 40044 180944 40050
rect 180892 39986 180944 39992
rect 179880 38752 179932 38758
rect 179880 38694 179932 38700
rect 177868 6886 177988 6914
rect 179064 6886 179368 6914
rect 171968 3528 172020 3534
rect 171968 3470 172020 3476
rect 172428 3528 172480 3534
rect 172428 3470 172480 3476
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 175188 3528 175240 3534
rect 175188 3470 175240 3476
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 176568 3528 176620 3534
rect 176568 3470 176620 3476
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 177764 3528 177816 3534
rect 177764 3470 177816 3476
rect 171980 480 172008 3470
rect 173176 480 173204 3470
rect 174280 480 174308 3470
rect 175476 480 175504 3470
rect 176672 480 176700 3470
rect 177868 480 177896 6886
rect 179064 480 179092 6886
rect 180076 3466 180104 39986
rect 181916 39778 181944 41806
rect 181904 39772 181956 39778
rect 181904 39714 181956 39720
rect 180708 39704 180760 39710
rect 180708 39646 180760 39652
rect 180720 3534 180748 39646
rect 182928 39642 182956 41806
rect 183940 39914 183968 41806
rect 183928 39908 183980 39914
rect 183928 39850 183980 39856
rect 184848 39772 184900 39778
rect 184848 39714 184900 39720
rect 182916 39636 182968 39642
rect 182916 39578 182968 39584
rect 183468 39636 183520 39642
rect 183468 39578 183520 39584
rect 182088 38956 182140 38962
rect 182088 38898 182140 38904
rect 182100 3534 182128 38898
rect 183480 3534 183508 39578
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 181444 3528 181496 3534
rect 181444 3470 181496 3476
rect 182088 3528 182140 3534
rect 182088 3470 182140 3476
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 180064 3460 180116 3466
rect 180064 3402 180116 3408
rect 180260 480 180288 3470
rect 181456 480 181484 3470
rect 182560 480 182588 3470
rect 184860 3262 184888 39714
rect 184952 39370 184980 41806
rect 184940 39364 184992 39370
rect 184940 39306 184992 39312
rect 185964 39234 185992 41806
rect 186976 39982 187004 41806
rect 186964 39976 187016 39982
rect 186964 39918 187016 39924
rect 187608 39908 187660 39914
rect 187608 39850 187660 39856
rect 186136 39364 186188 39370
rect 186136 39306 186188 39312
rect 185952 39228 186004 39234
rect 185952 39170 186004 39176
rect 184940 3528 184992 3534
rect 184940 3470 184992 3476
rect 183744 3256 183796 3262
rect 183744 3198 183796 3204
rect 184848 3256 184900 3262
rect 184848 3198 184900 3204
rect 183756 480 183784 3198
rect 184952 480 184980 3470
rect 186148 480 186176 39306
rect 186228 38888 186280 38894
rect 186228 38830 186280 38836
rect 186240 3534 186268 38830
rect 187620 6914 187648 39850
rect 187988 39574 188016 41806
rect 187976 39568 188028 39574
rect 187976 39510 188028 39516
rect 188988 39568 189040 39574
rect 188988 39510 189040 39516
rect 187344 6886 187648 6914
rect 186228 3528 186280 3534
rect 186228 3470 186280 3476
rect 187344 480 187372 6886
rect 189000 3534 189028 39510
rect 189092 39506 189120 41806
rect 190012 41806 190086 41834
rect 191024 41806 191098 41834
rect 192036 41806 192110 41834
rect 193048 41806 193122 41834
rect 194060 41806 194134 41834
rect 195164 41806 195238 41834
rect 196176 41806 196250 41834
rect 197188 41806 197262 41834
rect 198200 41806 198274 41834
rect 199212 41806 199286 41834
rect 200224 41806 200298 41834
rect 201236 41806 201310 41834
rect 202248 41806 202322 41834
rect 203260 41806 203334 41834
rect 204272 41806 204346 41834
rect 205284 41806 205358 41834
rect 206296 41806 206370 41834
rect 207308 41806 207382 41834
rect 208366 41834 208394 42092
rect 209378 41834 209406 42092
rect 210482 41834 210510 42092
rect 211494 41834 211522 42092
rect 208366 41806 208440 41834
rect 189080 39500 189132 39506
rect 189080 39442 189132 39448
rect 190012 39302 190040 41806
rect 190368 39976 190420 39982
rect 190368 39918 190420 39924
rect 190000 39296 190052 39302
rect 190000 39238 190052 39244
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 188988 3528 189040 3534
rect 188988 3470 189040 3476
rect 188540 480 188568 3470
rect 190380 3466 190408 39918
rect 191024 39846 191052 41806
rect 191012 39840 191064 39846
rect 191012 39782 191064 39788
rect 191748 39228 191800 39234
rect 191748 39170 191800 39176
rect 191760 3534 191788 39170
rect 192036 39166 192064 41806
rect 192024 39160 192076 39166
rect 192024 39102 192076 39108
rect 193048 39030 193076 41806
rect 193128 39296 193180 39302
rect 193128 39238 193180 39244
rect 193036 39024 193088 39030
rect 193036 38966 193088 38972
rect 193140 3534 193168 39238
rect 194060 39098 194088 41806
rect 195164 40050 195192 41806
rect 195152 40044 195204 40050
rect 195152 39986 195204 39992
rect 195888 39840 195940 39846
rect 195888 39782 195940 39788
rect 194416 39500 194468 39506
rect 194416 39442 194468 39448
rect 194048 39092 194100 39098
rect 194048 39034 194100 39040
rect 194428 16574 194456 39442
rect 194508 39160 194560 39166
rect 194508 39102 194560 39108
rect 194336 16546 194456 16574
rect 194336 3534 194364 16546
rect 194520 6914 194548 39102
rect 195900 6914 195928 39782
rect 196176 39438 196204 41806
rect 197188 39710 197216 41806
rect 197176 39704 197228 39710
rect 197176 39646 197228 39652
rect 196164 39432 196216 39438
rect 196164 39374 196216 39380
rect 197268 39432 197320 39438
rect 197268 39374 197320 39380
rect 194428 6886 194548 6914
rect 195624 6886 195928 6914
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 191748 3528 191800 3534
rect 191748 3470 191800 3476
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 193128 3528 193180 3534
rect 193128 3470 193180 3476
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 194324 3528 194376 3534
rect 194324 3470 194376 3476
rect 189724 3460 189776 3466
rect 189724 3402 189776 3408
rect 190368 3460 190420 3466
rect 190368 3402 190420 3408
rect 189736 480 189764 3402
rect 190840 480 190868 3470
rect 192036 480 192064 3470
rect 193232 480 193260 3470
rect 194428 480 194456 6886
rect 195624 480 195652 6886
rect 197280 3330 197308 39374
rect 198200 38962 198228 41806
rect 198648 39704 198700 39710
rect 198648 39646 198700 39652
rect 198188 38956 198240 38962
rect 198188 38898 198240 38904
rect 198660 3534 198688 39646
rect 199212 39642 199240 41806
rect 200028 40044 200080 40050
rect 200028 39986 200080 39992
rect 199200 39636 199252 39642
rect 199200 39578 199252 39584
rect 200040 3534 200068 39986
rect 200224 39778 200252 41806
rect 200212 39772 200264 39778
rect 200212 39714 200264 39720
rect 201236 38894 201264 41806
rect 201408 39772 201460 39778
rect 201408 39714 201460 39720
rect 201224 38888 201276 38894
rect 201224 38830 201276 38836
rect 197912 3528 197964 3534
rect 197912 3470 197964 3476
rect 198648 3528 198700 3534
rect 198648 3470 198700 3476
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 200028 3528 200080 3534
rect 200028 3470 200080 3476
rect 196808 3324 196860 3330
rect 196808 3266 196860 3272
rect 197268 3324 197320 3330
rect 197268 3266 197320 3272
rect 196820 480 196848 3266
rect 197924 480 197952 3470
rect 199120 480 199148 3470
rect 201420 3262 201448 39714
rect 202248 39370 202276 41806
rect 203260 39914 203288 41806
rect 203248 39908 203300 39914
rect 203248 39850 203300 39856
rect 204168 39908 204220 39914
rect 204168 39850 204220 39856
rect 202696 39636 202748 39642
rect 202696 39578 202748 39584
rect 202236 39364 202288 39370
rect 202236 39306 202288 39312
rect 201500 3528 201552 3534
rect 201500 3470 201552 3476
rect 200304 3256 200356 3262
rect 200304 3198 200356 3204
rect 201408 3256 201460 3262
rect 201408 3198 201460 3204
rect 200316 480 200344 3198
rect 201512 480 201540 3470
rect 202708 480 202736 39578
rect 202788 39092 202840 39098
rect 202788 39034 202840 39040
rect 202800 3534 202828 39034
rect 204180 6914 204208 39850
rect 204272 39574 204300 41806
rect 205284 39982 205312 41806
rect 205272 39976 205324 39982
rect 205272 39918 205324 39924
rect 205548 39976 205600 39982
rect 205548 39918 205600 39924
rect 204260 39568 204312 39574
rect 204260 39510 204312 39516
rect 203904 6886 204208 6914
rect 202788 3528 202840 3534
rect 202788 3470 202840 3476
rect 203904 480 203932 6886
rect 205560 3534 205588 39918
rect 206296 39234 206324 41806
rect 206928 39568 206980 39574
rect 206928 39510 206980 39516
rect 206284 39228 206336 39234
rect 206284 39170 206336 39176
rect 206940 3534 206968 39510
rect 207308 39302 207336 41806
rect 208412 39506 208440 41806
rect 209332 41806 209406 41834
rect 210436 41806 210510 41834
rect 211448 41806 211522 41834
rect 212506 41834 212534 42092
rect 213518 41834 213546 42092
rect 214530 41834 214558 42092
rect 215542 41834 215570 42092
rect 216554 41834 216582 42092
rect 217566 41834 217594 42092
rect 218578 41834 218606 42092
rect 219590 41834 219618 42092
rect 220602 41834 220630 42092
rect 221614 41834 221642 42092
rect 222626 41834 222654 42092
rect 223638 41834 223666 42092
rect 224650 41834 224678 42092
rect 225754 41834 225782 42092
rect 226766 41834 226794 42092
rect 227778 41834 227806 42092
rect 228790 41834 228818 42092
rect 229802 41834 229830 42092
rect 230814 41834 230842 42092
rect 212506 41806 212580 41834
rect 208400 39500 208452 39506
rect 208400 39442 208452 39448
rect 207296 39296 207348 39302
rect 207296 39238 207348 39244
rect 208308 39296 208360 39302
rect 208308 39238 208360 39244
rect 208320 3534 208348 39238
rect 209332 39166 209360 41806
rect 210436 39846 210464 41806
rect 210424 39840 210476 39846
rect 210424 39782 210476 39788
rect 211068 39840 211120 39846
rect 211068 39782 211120 39788
rect 210976 39364 211028 39370
rect 210976 39306 211028 39312
rect 209688 39228 209740 39234
rect 209688 39170 209740 39176
rect 209320 39160 209372 39166
rect 209320 39102 209372 39108
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 206192 3528 206244 3534
rect 206192 3470 206244 3476
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 207388 3528 207440 3534
rect 207388 3470 207440 3476
rect 208308 3528 208360 3534
rect 208308 3470 208360 3476
rect 205100 480 205128 3470
rect 206204 480 206232 3470
rect 207400 480 207428 3470
rect 209700 3058 209728 39170
rect 209780 3528 209832 3534
rect 209780 3470 209832 3476
rect 208584 3052 208636 3058
rect 208584 2994 208636 3000
rect 209688 3052 209740 3058
rect 209688 2994 209740 3000
rect 208596 480 208624 2994
rect 209792 480 209820 3470
rect 210988 480 211016 39306
rect 211080 3534 211108 39782
rect 211448 39438 211476 41806
rect 212552 39710 212580 41806
rect 213472 41806 213546 41834
rect 214484 41806 214558 41834
rect 215496 41806 215570 41834
rect 216508 41806 216582 41834
rect 217520 41806 217594 41834
rect 218532 41806 218606 41834
rect 219544 41806 219618 41834
rect 220556 41806 220630 41834
rect 221568 41806 221642 41834
rect 222580 41806 222654 41834
rect 223592 41806 223666 41834
rect 224604 41806 224678 41834
rect 225708 41806 225782 41834
rect 226720 41806 226794 41834
rect 227732 41806 227806 41834
rect 228744 41806 228818 41834
rect 229756 41806 229830 41834
rect 230768 41806 230842 41834
rect 231826 41834 231854 42092
rect 232838 41834 232866 42092
rect 233850 41834 233878 42092
rect 234862 41834 234890 42092
rect 235874 41834 235902 42092
rect 236886 41834 236914 42092
rect 237898 41834 237926 42092
rect 238910 41834 238938 42092
rect 239922 41834 239950 42092
rect 241026 41834 241054 42092
rect 242038 41834 242066 42092
rect 243050 41834 243078 42092
rect 244062 41834 244090 42092
rect 245074 41834 245102 42092
rect 246086 41834 246114 42092
rect 247098 41834 247126 42092
rect 248110 41834 248138 42092
rect 249122 41834 249150 42092
rect 250134 41834 250162 42092
rect 231826 41806 231900 41834
rect 213472 40050 213500 41806
rect 213460 40044 213512 40050
rect 213460 39986 213512 39992
rect 214484 39778 214512 41806
rect 214472 39772 214524 39778
rect 214472 39714 214524 39720
rect 212540 39704 212592 39710
rect 212540 39646 212592 39652
rect 215208 39500 215260 39506
rect 215208 39442 215260 39448
rect 211436 39432 211488 39438
rect 211436 39374 211488 39380
rect 213828 39432 213880 39438
rect 213828 39374 213880 39380
rect 212448 39160 212500 39166
rect 212448 39102 212500 39108
rect 212460 6914 212488 39102
rect 212184 6886 212488 6914
rect 211068 3528 211120 3534
rect 211068 3470 211120 3476
rect 212184 480 212212 6886
rect 213840 3534 213868 39374
rect 215220 3534 215248 39442
rect 215496 39098 215524 41806
rect 216508 39642 216536 41806
rect 217520 39914 217548 41806
rect 218532 39982 218560 41806
rect 218520 39976 218572 39982
rect 218520 39918 218572 39924
rect 217508 39908 217560 39914
rect 217508 39850 217560 39856
rect 217968 39908 218020 39914
rect 217968 39850 218020 39856
rect 216496 39636 216548 39642
rect 216496 39578 216548 39584
rect 216588 39636 216640 39642
rect 216588 39578 216640 39584
rect 215484 39092 215536 39098
rect 215484 39034 215536 39040
rect 216600 3534 216628 39578
rect 217980 3534 218008 39850
rect 219256 39772 219308 39778
rect 219256 39714 219308 39720
rect 219268 16574 219296 39714
rect 219348 39704 219400 39710
rect 219348 39646 219400 39652
rect 219176 16546 219296 16574
rect 219176 3534 219204 16546
rect 219360 6914 219388 39646
rect 219544 39574 219572 41806
rect 219532 39568 219584 39574
rect 219532 39510 219584 39516
rect 220556 39302 220584 41806
rect 220728 39568 220780 39574
rect 220728 39510 220780 39516
rect 220544 39296 220596 39302
rect 220544 39238 220596 39244
rect 220740 6914 220768 39510
rect 221568 39234 221596 41806
rect 222108 39976 222160 39982
rect 222108 39918 222160 39924
rect 221556 39228 221608 39234
rect 221556 39170 221608 39176
rect 219268 6886 219388 6914
rect 220464 6886 220768 6914
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213828 3528 213880 3534
rect 213828 3470 213880 3476
rect 214472 3528 214524 3534
rect 214472 3470 214524 3476
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 216864 3528 216916 3534
rect 216864 3470 216916 3476
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 219164 3528 219216 3534
rect 219164 3470 219216 3476
rect 213380 480 213408 3470
rect 214484 480 214512 3470
rect 215680 480 215708 3470
rect 216876 480 216904 3470
rect 218072 480 218100 3470
rect 219268 480 219296 6886
rect 220464 480 220492 6886
rect 222120 3330 222148 39918
rect 222580 39846 222608 41806
rect 223488 40044 223540 40050
rect 223488 39986 223540 39992
rect 222568 39840 222620 39846
rect 222568 39782 222620 39788
rect 223500 3534 223528 39986
rect 223592 39370 223620 41806
rect 223580 39364 223632 39370
rect 223580 39306 223632 39312
rect 224604 39166 224632 41806
rect 224868 39840 224920 39846
rect 224868 39782 224920 39788
rect 224592 39160 224644 39166
rect 224592 39102 224644 39108
rect 224880 3534 224908 39782
rect 225708 39438 225736 41806
rect 226720 39506 226748 41806
rect 227732 39642 227760 41806
rect 228744 39914 228772 41806
rect 228732 39908 228784 39914
rect 228732 39850 228784 39856
rect 229756 39778 229784 41806
rect 229744 39772 229796 39778
rect 229744 39714 229796 39720
rect 230388 39772 230440 39778
rect 230388 39714 230440 39720
rect 227720 39636 227772 39642
rect 227720 39578 227772 39584
rect 226708 39500 226760 39506
rect 226708 39442 226760 39448
rect 225696 39432 225748 39438
rect 225696 39374 225748 39380
rect 229008 39432 229060 39438
rect 229008 39374 229060 39380
rect 227536 39364 227588 39370
rect 227536 39306 227588 39312
rect 226248 39228 226300 39234
rect 226248 39170 226300 39176
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 221556 3324 221608 3330
rect 221556 3266 221608 3272
rect 222108 3324 222160 3330
rect 222108 3266 222160 3272
rect 221568 480 221596 3266
rect 222764 480 222792 3470
rect 223960 480 223988 3470
rect 226260 3262 226288 39170
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 225144 3256 225196 3262
rect 225144 3198 225196 3204
rect 226248 3256 226300 3262
rect 226248 3198 226300 3204
rect 225156 480 225184 3198
rect 226352 480 226380 3470
rect 227548 480 227576 39306
rect 227628 39296 227680 39302
rect 227628 39238 227680 39244
rect 227640 3534 227668 39238
rect 229020 6914 229048 39374
rect 228744 6886 229048 6914
rect 227628 3528 227680 3534
rect 227628 3470 227680 3476
rect 228744 480 228772 6886
rect 230400 3534 230428 39714
rect 230768 39710 230796 41806
rect 230756 39704 230808 39710
rect 230756 39646 230808 39652
rect 231768 39636 231820 39642
rect 231768 39578 231820 39584
rect 231780 3534 231808 39578
rect 231872 39574 231900 41806
rect 232792 41806 232866 41834
rect 233804 41806 233878 41834
rect 234816 41806 234890 41834
rect 235736 41806 235902 41834
rect 236840 41806 236914 41834
rect 237852 41806 237926 41834
rect 238864 41806 238938 41834
rect 239876 41806 239950 41834
rect 240980 41806 241054 41834
rect 241992 41806 242066 41834
rect 243004 41806 243078 41834
rect 244016 41806 244090 41834
rect 245028 41806 245102 41834
rect 246040 41806 246114 41834
rect 247052 41806 247126 41834
rect 248064 41806 248138 41834
rect 249076 41806 249150 41834
rect 250088 41806 250162 41834
rect 251146 41834 251174 42092
rect 252158 41834 252186 42092
rect 253170 41834 253198 42092
rect 254182 41834 254210 42092
rect 255194 41834 255222 42092
rect 256298 41834 256326 42092
rect 257310 41834 257338 42092
rect 258322 41834 258350 42092
rect 259334 41834 259362 42092
rect 260346 41834 260374 42092
rect 261358 41834 261386 42092
rect 262370 41834 262398 42092
rect 263382 41834 263410 42092
rect 264394 41834 264422 42092
rect 265406 41834 265434 42092
rect 266418 41834 266446 42092
rect 267430 41834 267458 42092
rect 268442 41834 268470 42092
rect 269454 41834 269482 42092
rect 251146 41806 251220 41834
rect 232792 39982 232820 41806
rect 233804 40050 233832 41806
rect 233792 40044 233844 40050
rect 233792 39986 233844 39992
rect 232780 39976 232832 39982
rect 232780 39918 232832 39924
rect 234816 39846 234844 41806
rect 234804 39840 234856 39846
rect 234804 39782 234856 39788
rect 233148 39704 233200 39710
rect 233148 39646 233200 39652
rect 231860 39568 231912 39574
rect 231860 39510 231912 39516
rect 233160 3534 233188 39646
rect 234528 39568 234580 39574
rect 234528 39510 234580 39516
rect 234540 3534 234568 39510
rect 235736 39234 235764 41806
rect 235908 39908 235960 39914
rect 235908 39850 235960 39856
rect 235816 39500 235868 39506
rect 235816 39442 235868 39448
rect 235724 39228 235776 39234
rect 235724 39170 235776 39176
rect 229836 3528 229888 3534
rect 229836 3470 229888 3476
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 229848 480 229876 3470
rect 231044 480 231072 3470
rect 232240 480 232268 3470
rect 233436 480 233464 3470
rect 234632 480 234660 3470
rect 235828 480 235856 39442
rect 235920 3534 235948 39850
rect 236840 39302 236868 41806
rect 237288 39840 237340 39846
rect 237288 39782 237340 39788
rect 236828 39296 236880 39302
rect 236828 39238 236880 39244
rect 237300 6914 237328 39782
rect 237852 39370 237880 41806
rect 238864 39438 238892 41806
rect 239876 39778 239904 41806
rect 239864 39772 239916 39778
rect 239864 39714 239916 39720
rect 240980 39642 241008 41806
rect 241428 39772 241480 39778
rect 241428 39714 241480 39720
rect 240968 39636 241020 39642
rect 240968 39578 241020 39584
rect 238852 39432 238904 39438
rect 238852 39374 238904 39380
rect 237840 39364 237892 39370
rect 237840 39306 237892 39312
rect 238668 39364 238720 39370
rect 238668 39306 238720 39312
rect 237024 6886 237328 6914
rect 235908 3528 235960 3534
rect 235908 3470 235960 3476
rect 237024 480 237052 6886
rect 238680 3534 238708 39306
rect 240048 39024 240100 39030
rect 240048 38966 240100 38972
rect 240060 3534 240088 38966
rect 241440 3534 241468 39714
rect 241992 39710 242020 41806
rect 242808 40044 242860 40050
rect 242808 39986 242860 39992
rect 241980 39704 242032 39710
rect 241980 39646 242032 39652
rect 238116 3528 238168 3534
rect 238116 3470 238168 3476
rect 238668 3528 238720 3534
rect 238668 3470 238720 3476
rect 239312 3528 239364 3534
rect 239312 3470 239364 3476
rect 240048 3528 240100 3534
rect 240048 3470 240100 3476
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 238128 480 238156 3470
rect 239324 480 239352 3470
rect 240520 480 240548 3470
rect 242820 3194 242848 39986
rect 243004 39574 243032 41806
rect 244016 39914 244044 41806
rect 244004 39908 244056 39914
rect 244004 39850 244056 39856
rect 244188 39704 244240 39710
rect 244188 39646 244240 39652
rect 242992 39568 243044 39574
rect 242992 39510 243044 39516
rect 244096 39432 244148 39438
rect 244096 39374 244148 39380
rect 244108 16574 244136 39374
rect 244016 16546 244136 16574
rect 244016 3534 244044 16546
rect 244200 6914 244228 39646
rect 245028 39506 245056 41806
rect 246040 39846 246068 41806
rect 246028 39840 246080 39846
rect 246028 39782 246080 39788
rect 245568 39568 245620 39574
rect 245568 39510 245620 39516
rect 245016 39500 245068 39506
rect 245016 39442 245068 39448
rect 244108 6886 244228 6914
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 244004 3528 244056 3534
rect 244004 3470 244056 3476
rect 241704 3188 241756 3194
rect 241704 3130 241756 3136
rect 242808 3188 242860 3194
rect 242808 3130 242860 3136
rect 241716 480 241744 3130
rect 242912 480 242940 3470
rect 244108 480 244136 6886
rect 245212 598 245424 626
rect 245212 480 245240 598
rect 245396 490 245424 598
rect 245580 490 245608 39510
rect 246948 39500 247000 39506
rect 246948 39442 247000 39448
rect 246960 3126 246988 39442
rect 247052 39370 247080 41806
rect 247040 39364 247092 39370
rect 247040 39306 247092 39312
rect 248064 39030 248092 41806
rect 248328 39840 248380 39846
rect 248328 39782 248380 39788
rect 248052 39024 248104 39030
rect 248052 38966 248104 38972
rect 248340 3534 248368 39782
rect 249076 39778 249104 41806
rect 250088 40050 250116 41806
rect 250076 40044 250128 40050
rect 250076 39986 250128 39992
rect 249064 39772 249116 39778
rect 249064 39714 249116 39720
rect 251192 39438 251220 41806
rect 252112 41806 252186 41834
rect 253124 41806 253198 41834
rect 254136 41806 254210 41834
rect 255148 41806 255222 41834
rect 256252 41806 256326 41834
rect 257264 41806 257338 41834
rect 258276 41806 258350 41834
rect 259288 41806 259362 41834
rect 260300 41806 260374 41834
rect 261312 41806 261386 41834
rect 262324 41806 262398 41834
rect 263336 41806 263410 41834
rect 264348 41806 264422 41834
rect 265360 41806 265434 41834
rect 266372 41806 266446 41834
rect 267384 41806 267458 41834
rect 268396 41806 268470 41834
rect 269408 41806 269482 41834
rect 270466 41834 270494 42092
rect 271570 41834 271598 42092
rect 272582 41834 272610 42092
rect 273594 41834 273622 42092
rect 270466 41806 270540 41834
rect 252112 39710 252140 41806
rect 252100 39704 252152 39710
rect 252100 39646 252152 39652
rect 253124 39574 253152 41806
rect 253848 40044 253900 40050
rect 253848 39986 253900 39992
rect 253112 39568 253164 39574
rect 253112 39510 253164 39516
rect 251180 39432 251232 39438
rect 251180 39374 251232 39380
rect 252376 39092 252428 39098
rect 252376 39034 252428 39040
rect 251088 39024 251140 39030
rect 251088 38966 251140 38972
rect 249708 38888 249760 38894
rect 249708 38830 249760 38836
rect 247592 3528 247644 3534
rect 247592 3470 247644 3476
rect 248328 3528 248380 3534
rect 248328 3470 248380 3476
rect 246396 3120 246448 3126
rect 246396 3062 246448 3068
rect 246948 3120 247000 3126
rect 246948 3062 247000 3068
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245396 462 245608 490
rect 246408 480 246436 3062
rect 247604 480 247632 3470
rect 249720 3058 249748 38830
rect 251100 3534 251128 38966
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 248788 3052 248840 3058
rect 248788 2994 248840 3000
rect 249708 3052 249760 3058
rect 249708 2994 249760 3000
rect 248800 480 248828 2994
rect 249996 480 250024 3470
rect 251192 480 251220 3470
rect 252388 480 252416 39034
rect 252468 38956 252520 38962
rect 252468 38898 252520 38904
rect 252480 3534 252508 38898
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 253492 598 253704 626
rect 253492 480 253520 598
rect 253676 490 253704 598
rect 253860 490 253888 39986
rect 254136 39506 254164 41806
rect 255148 39846 255176 41806
rect 255136 39840 255188 39846
rect 255136 39782 255188 39788
rect 254124 39500 254176 39506
rect 254124 39442 254176 39448
rect 255228 39500 255280 39506
rect 255228 39442 255280 39448
rect 255240 3534 255268 39442
rect 256252 38894 256280 41806
rect 256608 39568 256660 39574
rect 256608 39510 256660 39516
rect 256240 38888 256292 38894
rect 256240 38830 256292 38836
rect 256620 3534 256648 39510
rect 257264 39030 257292 41806
rect 257988 39772 258040 39778
rect 257988 39714 258040 39720
rect 257252 39024 257304 39030
rect 257252 38966 257304 38972
rect 258000 3534 258028 39714
rect 258276 38962 258304 41806
rect 259288 39098 259316 41806
rect 260300 40050 260328 41806
rect 260288 40044 260340 40050
rect 260288 39986 260340 39992
rect 261312 39506 261340 41806
rect 262324 39574 262352 41806
rect 263336 39778 263364 41806
rect 263324 39772 263376 39778
rect 263324 39714 263376 39720
rect 262312 39568 262364 39574
rect 262312 39510 262364 39516
rect 261300 39500 261352 39506
rect 261300 39442 261352 39448
rect 264348 39098 264376 41806
rect 264888 39636 264940 39642
rect 264888 39578 264940 39584
rect 259276 39092 259328 39098
rect 259276 39034 259328 39040
rect 259368 39092 259420 39098
rect 259368 39034 259420 39040
rect 264336 39092 264388 39098
rect 264336 39034 264388 39040
rect 258264 38956 258316 38962
rect 258264 38898 258316 38904
rect 259380 3534 259408 39034
rect 260748 39024 260800 39030
rect 260748 38966 260800 38972
rect 260656 38820 260708 38826
rect 260656 38762 260708 38768
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 255228 3528 255280 3534
rect 255228 3470 255280 3476
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 256608 3528 256660 3534
rect 256608 3470 256660 3476
rect 257068 3528 257120 3534
rect 257068 3470 257120 3476
rect 257988 3528 258040 3534
rect 257988 3470 258040 3476
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 253676 462 253888 490
rect 254688 480 254716 3470
rect 255884 480 255912 3470
rect 257080 480 257108 3470
rect 258276 480 258304 3470
rect 259472 480 259500 3470
rect 260668 480 260696 38762
rect 260760 3534 260788 38966
rect 263508 38956 263560 38962
rect 263508 38898 263560 38904
rect 262128 38888 262180 38894
rect 262128 38830 262180 38836
rect 260748 3528 260800 3534
rect 260748 3470 260800 3476
rect 261772 598 261984 626
rect 261772 480 261800 598
rect 261956 490 261984 598
rect 262140 490 262168 38830
rect 263520 3534 263548 38898
rect 264900 3534 264928 39578
rect 265360 39030 265388 41806
rect 265348 39024 265400 39030
rect 265348 38966 265400 38972
rect 266372 38826 266400 41806
rect 267004 39500 267056 39506
rect 267004 39442 267056 39448
rect 266360 38820 266412 38826
rect 266360 38762 266412 38768
rect 262956 3528 263008 3534
rect 262956 3470 263008 3476
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 264888 3528 264940 3534
rect 264888 3470 264940 3476
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 261956 462 262168 490
rect 262968 480 262996 3470
rect 264164 480 264192 3470
rect 265348 3460 265400 3466
rect 265348 3402 265400 3408
rect 265360 480 265388 3402
rect 266556 480 266584 3470
rect 267016 3466 267044 39442
rect 267384 38894 267412 41806
rect 267648 39704 267700 39710
rect 267648 39646 267700 39652
rect 267372 38888 267424 38894
rect 267372 38830 267424 38836
rect 267660 3534 267688 39646
rect 268396 38962 268424 41806
rect 269408 39642 269436 41806
rect 269396 39636 269448 39642
rect 269396 39578 269448 39584
rect 270512 39506 270540 41806
rect 271524 41806 271598 41834
rect 272536 41806 272610 41834
rect 273548 41806 273622 41834
rect 274606 41834 274634 42092
rect 275618 41834 275646 42092
rect 276630 41834 276658 42092
rect 277642 41834 277670 42092
rect 278654 41834 278682 42092
rect 279666 41834 279694 42092
rect 280678 41834 280706 42092
rect 281690 41834 281718 42092
rect 282702 41834 282730 42092
rect 283714 41834 283742 42092
rect 284726 41834 284754 42092
rect 285738 41834 285766 42092
rect 286842 41834 286870 42092
rect 287854 41834 287882 42092
rect 288866 41834 288894 42092
rect 289878 41834 289906 42092
rect 290890 41834 290918 42092
rect 291902 41834 291930 42092
rect 292914 41834 292942 42092
rect 274606 41806 274680 41834
rect 271524 39710 271552 41806
rect 271512 39704 271564 39710
rect 271512 39646 271564 39652
rect 270500 39500 270552 39506
rect 270500 39442 270552 39448
rect 269028 39092 269080 39098
rect 269028 39034 269080 39040
rect 268384 38956 268436 38962
rect 268384 38898 268436 38904
rect 268936 38888 268988 38894
rect 268936 38830 268988 38836
rect 268948 3602 268976 38830
rect 267740 3596 267792 3602
rect 267740 3538 267792 3544
rect 268936 3596 268988 3602
rect 268936 3538 268988 3544
rect 267648 3528 267700 3534
rect 267648 3470 267700 3476
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 267752 480 267780 3538
rect 269040 3482 269068 39034
rect 271788 39024 271840 39030
rect 271788 38966 271840 38972
rect 270408 38956 270460 38962
rect 270408 38898 270460 38904
rect 268856 3454 269068 3482
rect 268856 480 268884 3454
rect 270052 598 270264 626
rect 270052 480 270080 598
rect 270236 490 270264 598
rect 270420 490 270448 38898
rect 271800 3330 271828 38966
rect 272536 38894 272564 41806
rect 273548 39098 273576 41806
rect 274548 39228 274600 39234
rect 274548 39170 274600 39176
rect 273536 39092 273588 39098
rect 273536 39034 273588 39040
rect 272524 38888 272576 38894
rect 272524 38830 272576 38836
rect 273168 38888 273220 38894
rect 273168 38830 273220 38836
rect 273180 3534 273208 38830
rect 274560 3534 274588 39170
rect 274652 38962 274680 41806
rect 275572 41806 275646 41834
rect 276584 41806 276658 41834
rect 277596 41806 277670 41834
rect 278608 41806 278682 41834
rect 279620 41806 279694 41834
rect 280632 41806 280706 41834
rect 281644 41806 281718 41834
rect 282656 41806 282730 41834
rect 283668 41806 283742 41834
rect 284680 41806 284754 41834
rect 285692 41806 285766 41834
rect 285876 41806 286870 41834
rect 287808 41806 287882 41834
rect 288820 41806 288894 41834
rect 289832 41806 289906 41834
rect 290844 41806 290918 41834
rect 291304 41806 291930 41834
rect 292592 41806 292942 41834
rect 293926 41834 293954 42092
rect 294938 41834 294966 42092
rect 295950 41834 295978 42092
rect 296962 41834 296990 42092
rect 297974 41834 298002 42092
rect 298986 41834 299014 42092
rect 299998 41834 300026 42092
rect 301102 41834 301130 42092
rect 302114 41834 302142 42092
rect 303126 41834 303154 42092
rect 304138 41834 304166 42092
rect 305150 41834 305178 42092
rect 293926 41806 294000 41834
rect 275572 39030 275600 41806
rect 275928 39976 275980 39982
rect 275928 39918 275980 39924
rect 275560 39024 275612 39030
rect 275560 38966 275612 38972
rect 274640 38956 274692 38962
rect 274640 38898 274692 38904
rect 275940 3534 275968 39918
rect 276584 38894 276612 41806
rect 277308 40044 277360 40050
rect 277308 39986 277360 39992
rect 277216 39364 277268 39370
rect 277216 39306 277268 39312
rect 276572 38888 276624 38894
rect 276572 38830 276624 38836
rect 277228 6914 277256 39306
rect 277136 6886 277256 6914
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 273168 3528 273220 3534
rect 273168 3470 273220 3476
rect 273628 3528 273680 3534
rect 273628 3470 273680 3476
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 274824 3528 274876 3534
rect 274824 3470 274876 3476
rect 275928 3528 275980 3534
rect 275928 3470 275980 3476
rect 271236 3324 271288 3330
rect 271236 3266 271288 3272
rect 271788 3324 271840 3330
rect 271788 3266 271840 3272
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270236 462 270448 490
rect 271248 480 271276 3266
rect 272444 480 272472 3470
rect 273640 480 273668 3470
rect 274836 480 274864 3470
rect 276020 3324 276072 3330
rect 276020 3266 276072 3272
rect 276032 480 276060 3266
rect 277136 480 277164 6886
rect 277320 3330 277348 39986
rect 277596 39234 277624 41806
rect 278608 39982 278636 41806
rect 279620 40050 279648 41806
rect 279608 40044 279660 40050
rect 279608 39986 279660 39992
rect 278596 39976 278648 39982
rect 278596 39918 278648 39924
rect 280632 39370 280660 41806
rect 280620 39364 280672 39370
rect 280620 39306 280672 39312
rect 277584 39228 277636 39234
rect 277584 39170 277636 39176
rect 281448 38956 281500 38962
rect 281448 38898 281500 38904
rect 280068 38752 280120 38758
rect 280068 38694 280120 38700
rect 278688 38684 278740 38690
rect 278688 38626 278740 38632
rect 277308 3324 277360 3330
rect 277308 3266 277360 3272
rect 278332 598 278544 626
rect 278332 480 278360 598
rect 278516 490 278544 598
rect 278700 490 278728 38626
rect 280080 3330 280108 38694
rect 281460 3534 281488 38898
rect 281644 38690 281672 41806
rect 282656 38758 282684 41806
rect 282828 39024 282880 39030
rect 282828 38966 282880 38972
rect 282644 38752 282696 38758
rect 282644 38694 282696 38700
rect 281632 38684 281684 38690
rect 281632 38626 281684 38632
rect 282840 3534 282868 38966
rect 283668 38962 283696 41806
rect 284680 39030 284708 41806
rect 285588 39976 285640 39982
rect 285588 39918 285640 39924
rect 284668 39024 284720 39030
rect 284668 38966 284720 38972
rect 284944 39024 284996 39030
rect 284944 38966 284996 38972
rect 283656 38956 283708 38962
rect 283656 38898 283708 38904
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 281908 3528 281960 3534
rect 281908 3470 281960 3476
rect 282828 3528 282880 3534
rect 282828 3470 282880 3476
rect 279516 3324 279568 3330
rect 279516 3266 279568 3272
rect 280068 3324 280120 3330
rect 280068 3266 280120 3272
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 278516 462 278728 490
rect 279528 480 279556 3266
rect 280724 480 280752 3470
rect 281920 480 281948 3470
rect 284956 3058 284984 38966
rect 285600 6914 285628 39918
rect 285692 39030 285720 41806
rect 285680 39024 285732 39030
rect 285680 38966 285732 38972
rect 285416 6886 285628 6914
rect 283104 3052 283156 3058
rect 283104 2994 283156 3000
rect 284944 3052 284996 3058
rect 284944 2994 284996 3000
rect 283116 480 283144 2994
rect 284300 2984 284352 2990
rect 284300 2926 284352 2932
rect 284312 480 284340 2926
rect 285416 480 285444 6886
rect 285876 2990 285904 41806
rect 286968 40044 287020 40050
rect 286968 39986 287020 39992
rect 285864 2984 285916 2990
rect 285864 2926 285916 2932
rect 286612 598 286824 626
rect 286612 480 286640 598
rect 286796 490 286824 598
rect 286980 490 287008 39986
rect 287808 39982 287836 41806
rect 288820 40050 288848 41806
rect 288808 40044 288860 40050
rect 288808 39986 288860 39992
rect 287796 39976 287848 39982
rect 287796 39918 287848 39924
rect 289728 39024 289780 39030
rect 289728 38966 289780 38972
rect 288348 38956 288400 38962
rect 288348 38898 288400 38904
rect 288360 3534 288388 38898
rect 289740 3534 289768 38966
rect 289832 38962 289860 41806
rect 290844 39030 290872 41806
rect 290832 39024 290884 39030
rect 290832 38966 290884 38972
rect 289820 38956 289872 38962
rect 289820 38898 289872 38904
rect 291304 3534 291332 41806
rect 292592 38978 292620 41806
rect 292500 38950 292620 38978
rect 292500 3534 292528 38950
rect 287796 3528 287848 3534
rect 287796 3470 287848 3476
rect 288348 3528 288400 3534
rect 288348 3470 288400 3476
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 291292 3528 291344 3534
rect 291292 3470 291344 3476
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 292488 3528 292540 3534
rect 292488 3470 292540 3476
rect 293684 3528 293736 3534
rect 293684 3470 293736 3476
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 286796 462 287008 490
rect 287808 480 287836 3470
rect 289004 480 289032 3470
rect 290200 480 290228 3470
rect 291396 480 291424 3470
rect 292580 2916 292632 2922
rect 292580 2858 292632 2864
rect 292592 480 292620 2858
rect 293696 480 293724 3470
rect 293972 2922 294000 41806
rect 294248 41806 294966 41834
rect 295444 41806 295978 41834
rect 296732 41806 296990 41834
rect 297928 41806 298002 41834
rect 298112 41806 299014 41834
rect 299492 41806 300026 41834
rect 300872 41806 301130 41834
rect 301240 41806 302142 41834
rect 302252 41806 303154 41834
rect 304092 41806 304166 41834
rect 305012 41806 305178 41834
rect 306162 41834 306190 42092
rect 307174 41834 307202 42092
rect 308186 41834 308214 42092
rect 309198 41834 309226 42092
rect 306162 41806 306328 41834
rect 307174 41806 307248 41834
rect 294248 3534 294276 41806
rect 294236 3528 294288 3534
rect 294236 3470 294288 3476
rect 293960 2916 294012 2922
rect 293960 2858 294012 2864
rect 295444 2854 295472 41806
rect 296732 39930 296760 41806
rect 296640 39902 296760 39930
rect 296640 3534 296668 39902
rect 297928 39030 297956 41806
rect 296720 39024 296772 39030
rect 296720 38966 296772 38972
rect 297916 39024 297968 39030
rect 297916 38966 297968 38972
rect 296732 16574 296760 38966
rect 296732 16546 297312 16574
rect 296076 3528 296128 3534
rect 296076 3470 296128 3476
rect 296628 3528 296680 3534
rect 296628 3470 296680 3476
rect 294880 2848 294932 2854
rect 294880 2790 294932 2796
rect 295432 2848 295484 2854
rect 295432 2790 295484 2796
rect 294892 480 294920 2790
rect 296088 480 296116 3470
rect 297284 480 297312 16546
rect 298112 490 298140 41806
rect 299492 16574 299520 41806
rect 300872 38978 300900 41806
rect 300780 38950 300900 38978
rect 299492 16546 299704 16574
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 16546
rect 300780 480 300808 38950
rect 301240 26234 301268 41806
rect 300964 26206 301268 26234
rect 300964 3534 300992 26206
rect 302252 3534 302280 41806
rect 304092 39030 304120 41806
rect 303620 39024 303672 39030
rect 303620 38966 303672 38972
rect 304080 39024 304132 39030
rect 304080 38966 304132 38972
rect 303632 16574 303660 38966
rect 303632 16546 303936 16574
rect 300952 3528 301004 3534
rect 300952 3470 301004 3476
rect 301964 3528 302016 3534
rect 301964 3470 302016 3476
rect 302240 3528 302292 3534
rect 302240 3470 302292 3476
rect 303160 3528 303212 3534
rect 303160 3470 303212 3476
rect 301976 480 302004 3470
rect 303172 480 303200 3470
rect 303908 490 303936 16546
rect 305012 3330 305040 41806
rect 305000 3324 305052 3330
rect 305000 3266 305052 3272
rect 305552 3324 305604 3330
rect 305552 3266 305604 3272
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3266
rect 306300 2802 306328 41806
rect 307220 39030 307248 41806
rect 307772 41806 308214 41834
rect 309152 41806 309226 41834
rect 310210 41834 310238 42092
rect 311222 41834 311250 42092
rect 312234 41834 312262 42092
rect 313246 41834 313274 42092
rect 314258 41834 314286 42092
rect 315270 41834 315298 42092
rect 316374 41834 316402 42092
rect 317386 41834 317414 42092
rect 318398 41834 318426 42092
rect 319410 41834 319438 42092
rect 320422 41834 320450 42092
rect 321434 41834 321462 42092
rect 310210 41806 310468 41834
rect 311222 41806 311296 41834
rect 312234 41806 312308 41834
rect 313246 41806 313320 41834
rect 314258 41806 314516 41834
rect 315270 41806 315344 41834
rect 316374 41806 316448 41834
rect 317386 41806 317460 41834
rect 318398 41806 318656 41834
rect 319410 41806 319484 41834
rect 320422 41806 320496 41834
rect 307208 39024 307260 39030
rect 307208 38966 307260 38972
rect 307668 39024 307720 39030
rect 307668 38966 307720 38972
rect 307680 3482 307708 38966
rect 307772 3602 307800 41806
rect 307760 3596 307812 3602
rect 307760 3538 307812 3544
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 307680 3454 307984 3482
rect 306300 2774 306420 2802
rect 306392 490 306420 2774
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 3454
rect 309060 480 309088 3538
rect 309152 3534 309180 41806
rect 310440 3534 310468 41806
rect 311268 39030 311296 41806
rect 311256 39024 311308 39030
rect 311256 38966 311308 38972
rect 311808 39024 311860 39030
rect 311808 38966 311860 38972
rect 311820 3534 311848 38966
rect 312280 38758 312308 41806
rect 313292 39030 313320 41806
rect 313280 39024 313332 39030
rect 313280 38966 313332 38972
rect 312268 38752 312320 38758
rect 312268 38694 312320 38700
rect 313464 38752 313516 38758
rect 313464 38694 313516 38700
rect 313476 16574 313504 38694
rect 313476 16546 313872 16574
rect 309140 3528 309192 3534
rect 309140 3470 309192 3476
rect 310244 3528 310296 3534
rect 310244 3470 310296 3476
rect 310428 3528 310480 3534
rect 310428 3470 310480 3476
rect 311440 3528 311492 3534
rect 311440 3470 311492 3476
rect 311808 3528 311860 3534
rect 311808 3470 311860 3476
rect 312636 3528 312688 3534
rect 312636 3470 312688 3476
rect 310256 480 310284 3470
rect 311452 480 311480 3470
rect 312648 480 312676 3470
rect 313844 480 313872 16546
rect 314488 2990 314516 41806
rect 315316 40050 315344 41806
rect 315304 40044 315356 40050
rect 315304 39986 315356 39992
rect 316132 40044 316184 40050
rect 316132 39986 316184 39992
rect 314568 39024 314620 39030
rect 314568 38966 314620 38972
rect 314580 3534 314608 38966
rect 316144 16574 316172 39986
rect 316420 39030 316448 41806
rect 317432 39030 317460 41806
rect 316408 39024 316460 39030
rect 316408 38966 316460 38972
rect 317328 39024 317380 39030
rect 317328 38966 317380 38972
rect 317420 39024 317472 39030
rect 317420 38966 317472 38972
rect 316144 16546 317276 16574
rect 314568 3528 314620 3534
rect 314568 3470 314620 3476
rect 315028 3528 315080 3534
rect 315028 3470 315080 3476
rect 314476 2984 314528 2990
rect 314476 2926 314528 2932
rect 315040 480 315068 3470
rect 317248 3346 317276 16546
rect 317340 3534 317368 38966
rect 317328 3528 317380 3534
rect 317328 3470 317380 3476
rect 318524 3528 318576 3534
rect 318524 3470 318576 3476
rect 317248 3318 317368 3346
rect 316224 2984 316276 2990
rect 316224 2926 316276 2932
rect 316236 480 316264 2926
rect 317340 480 317368 3318
rect 318536 480 318564 3470
rect 318628 3058 318656 41806
rect 318708 39024 318760 39030
rect 318708 38966 318760 38972
rect 318720 3534 318748 38966
rect 319456 38962 319484 41806
rect 320468 39030 320496 41806
rect 321388 41806 321462 41834
rect 322446 41834 322474 42092
rect 323458 41834 323486 42092
rect 324470 41834 324498 42092
rect 325482 41834 325510 42092
rect 326494 41834 326522 42092
rect 327506 41834 327534 42092
rect 328518 41834 328546 42092
rect 329530 41834 329558 42092
rect 330542 41834 330570 42092
rect 331646 41834 331674 42092
rect 332658 41834 332686 42092
rect 333670 41834 333698 42092
rect 334682 41834 334710 42092
rect 335694 41834 335722 42092
rect 336706 41834 336734 42092
rect 337718 41834 337746 42092
rect 338730 41834 338758 42092
rect 339742 41834 339770 42092
rect 340754 41834 340782 42092
rect 322446 41806 322888 41834
rect 323458 41806 323532 41834
rect 324470 41806 324544 41834
rect 325482 41806 325648 41834
rect 326494 41806 326568 41834
rect 327506 41806 327580 41834
rect 328518 41806 328592 41834
rect 329530 41806 329696 41834
rect 330542 41806 330616 41834
rect 331646 41806 331720 41834
rect 332658 41806 332732 41834
rect 333670 41806 333744 41834
rect 334682 41806 334756 41834
rect 335694 41806 335768 41834
rect 336706 41806 336780 41834
rect 337718 41806 338068 41834
rect 338730 41806 338804 41834
rect 339742 41806 339816 41834
rect 320456 39024 320508 39030
rect 320456 38966 320508 38972
rect 319444 38956 319496 38962
rect 319444 38898 319496 38904
rect 318708 3528 318760 3534
rect 318708 3470 318760 3476
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 318616 3052 318668 3058
rect 318616 2994 318668 3000
rect 319732 480 319760 3470
rect 321388 3194 321416 41806
rect 321468 39024 321520 39030
rect 321468 38966 321520 38972
rect 321376 3188 321428 3194
rect 321376 3130 321428 3136
rect 320916 3052 320968 3058
rect 320916 2994 320968 3000
rect 320928 480 320956 2994
rect 321480 2990 321508 38966
rect 321652 38956 321704 38962
rect 321652 38898 321704 38904
rect 321664 16574 321692 38898
rect 321664 16546 322152 16574
rect 321468 2984 321520 2990
rect 321468 2926 321520 2932
rect 322124 480 322152 16546
rect 322860 3262 322888 41806
rect 323504 39030 323532 41806
rect 324516 39030 324544 41806
rect 323492 39024 323544 39030
rect 323492 38966 323544 38972
rect 324228 39024 324280 39030
rect 324228 38966 324280 38972
rect 324504 39024 324556 39030
rect 324504 38966 324556 38972
rect 325516 39024 325568 39030
rect 325516 38966 325568 38972
rect 322848 3256 322900 3262
rect 322848 3198 322900 3204
rect 323308 2984 323360 2990
rect 323308 2926 323360 2932
rect 323320 480 323348 2926
rect 324240 2922 324268 38966
rect 325528 3330 325556 38966
rect 325620 3466 325648 41806
rect 326540 39030 326568 41806
rect 327552 39030 327580 41806
rect 328564 39030 328592 41806
rect 326528 39024 326580 39030
rect 326528 38966 326580 38972
rect 326988 39024 327040 39030
rect 326988 38966 327040 38972
rect 327540 39024 327592 39030
rect 327540 38966 327592 38972
rect 328368 39024 328420 39030
rect 328368 38966 328420 38972
rect 328552 39024 328604 39030
rect 328552 38966 328604 38972
rect 325608 3460 325660 3466
rect 325608 3402 325660 3408
rect 325516 3324 325568 3330
rect 325516 3266 325568 3272
rect 325608 3256 325660 3262
rect 325608 3198 325660 3204
rect 324412 3188 324464 3194
rect 324412 3130 324464 3136
rect 324228 2916 324280 2922
rect 324228 2858 324280 2864
rect 324424 480 324452 3130
rect 325620 480 325648 3198
rect 327000 3194 327028 38966
rect 328380 3602 328408 38966
rect 328368 3596 328420 3602
rect 328368 3538 328420 3544
rect 329196 3460 329248 3466
rect 329196 3402 329248 3408
rect 328000 3324 328052 3330
rect 328000 3266 328052 3272
rect 326988 3188 327040 3194
rect 326988 3130 327040 3136
rect 326804 2916 326856 2922
rect 326804 2858 326856 2864
rect 326816 480 326844 2858
rect 328012 480 328040 3266
rect 329208 480 329236 3402
rect 329668 3398 329696 41806
rect 330588 39030 330616 41806
rect 331692 39030 331720 41806
rect 332704 39506 332732 41806
rect 332692 39500 332744 39506
rect 332692 39442 332744 39448
rect 333716 39030 333744 41806
rect 334728 39030 334756 41806
rect 335740 39030 335768 41806
rect 336004 39500 336056 39506
rect 336004 39442 336056 39448
rect 329748 39024 329800 39030
rect 329748 38966 329800 38972
rect 330576 39024 330628 39030
rect 330576 38966 330628 38972
rect 331128 39024 331180 39030
rect 331128 38966 331180 38972
rect 331680 39024 331732 39030
rect 331680 38966 331732 38972
rect 332508 39024 332560 39030
rect 332508 38966 332560 38972
rect 333704 39024 333756 39030
rect 333704 38966 333756 38972
rect 334624 39024 334676 39030
rect 334624 38966 334676 38972
rect 334716 39024 334768 39030
rect 334716 38966 334768 38972
rect 335268 39024 335320 39030
rect 335268 38966 335320 38972
rect 335728 39024 335780 39030
rect 335728 38966 335780 38972
rect 329760 3534 329788 38966
rect 329748 3528 329800 3534
rect 329748 3470 329800 3476
rect 331140 3466 331168 38966
rect 331588 3596 331640 3602
rect 331588 3538 331640 3544
rect 331128 3460 331180 3466
rect 331128 3402 331180 3408
rect 329656 3392 329708 3398
rect 329656 3334 329708 3340
rect 330392 3188 330444 3194
rect 330392 3130 330444 3136
rect 330404 480 330432 3130
rect 331600 480 331628 3538
rect 332520 3194 332548 38966
rect 334636 3670 334664 38966
rect 334624 3664 334676 3670
rect 334624 3606 334676 3612
rect 332692 3528 332744 3534
rect 332692 3470 332744 3476
rect 332508 3188 332560 3194
rect 332508 3130 332560 3136
rect 332704 480 332732 3470
rect 335280 3466 335308 38966
rect 336016 3534 336044 39442
rect 336648 39024 336700 39030
rect 336648 38966 336700 38972
rect 336660 3602 336688 38966
rect 336752 38894 336780 41806
rect 336740 38888 336792 38894
rect 336740 38830 336792 38836
rect 336648 3596 336700 3602
rect 336648 3538 336700 3544
rect 336004 3528 336056 3534
rect 336004 3470 336056 3476
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 335084 3460 335136 3466
rect 335084 3402 335136 3408
rect 335268 3460 335320 3466
rect 335268 3402 335320 3408
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 335096 480 335124 3402
rect 336280 3188 336332 3194
rect 336280 3130 336332 3136
rect 336292 480 336320 3130
rect 337488 480 337516 3470
rect 338040 3330 338068 41806
rect 338776 39030 338804 41806
rect 339788 39030 339816 41806
rect 340708 41806 340782 41834
rect 341766 41834 341794 42092
rect 342778 41834 342806 42092
rect 343790 41834 343818 42092
rect 344802 41834 344830 42092
rect 345814 41834 345842 42092
rect 346918 41834 346946 42092
rect 347930 41834 347958 42092
rect 348942 41834 348970 42092
rect 349954 41834 349982 42092
rect 350966 41834 350994 42092
rect 351978 41834 352006 42092
rect 352990 41834 353018 42092
rect 354002 41834 354030 42092
rect 355014 41834 355042 42092
rect 356026 41834 356054 42092
rect 357038 41834 357066 42092
rect 358050 41834 358078 42092
rect 359062 41834 359090 42092
rect 360074 41834 360102 42092
rect 341766 41806 342208 41834
rect 342778 41806 342852 41834
rect 343790 41806 343864 41834
rect 344802 41806 344968 41834
rect 345814 41806 345888 41834
rect 346918 41806 346992 41834
rect 347930 41806 348004 41834
rect 348942 41806 349108 41834
rect 349954 41806 350028 41834
rect 350966 41806 351040 41834
rect 351978 41806 352052 41834
rect 352990 41806 353156 41834
rect 354002 41806 354076 41834
rect 355014 41806 355088 41834
rect 356026 41806 356100 41834
rect 357038 41806 357296 41834
rect 358050 41806 358124 41834
rect 359062 41806 359136 41834
rect 338764 39024 338816 39030
rect 338764 38966 338816 38972
rect 339408 39024 339460 39030
rect 339408 38966 339460 38972
rect 339776 39024 339828 39030
rect 339776 38966 339828 38972
rect 338764 38888 338816 38894
rect 338764 38830 338816 38836
rect 338672 3664 338724 3670
rect 338672 3606 338724 3612
rect 338028 3324 338080 3330
rect 338028 3266 338080 3272
rect 338684 480 338712 3606
rect 338776 3262 338804 38830
rect 339420 3398 339448 38966
rect 340708 4078 340736 41806
rect 340788 39024 340840 39030
rect 340788 38966 340840 38972
rect 340696 4072 340748 4078
rect 340696 4014 340748 4020
rect 339868 3460 339920 3466
rect 339868 3402 339920 3408
rect 339408 3392 339460 3398
rect 339408 3334 339460 3340
rect 338764 3256 338816 3262
rect 338764 3198 338816 3204
rect 339880 480 339908 3402
rect 340800 3058 340828 38966
rect 342180 6914 342208 41806
rect 342824 39030 342852 41806
rect 343836 39370 343864 41806
rect 343824 39364 343876 39370
rect 343824 39306 343876 39312
rect 342812 39024 342864 39030
rect 342812 38966 342864 38972
rect 343548 39024 343600 39030
rect 343548 38966 343600 38972
rect 342088 6886 342208 6914
rect 340972 3596 341024 3602
rect 340972 3538 341024 3544
rect 340788 3052 340840 3058
rect 340788 2994 340840 3000
rect 340984 480 341012 3538
rect 342088 3534 342116 6886
rect 343560 3942 343588 38966
rect 343548 3936 343600 3942
rect 343548 3878 343600 3884
rect 344940 3874 344968 41806
rect 345860 39030 345888 41806
rect 346964 39030 346992 41806
rect 347976 39030 348004 41806
rect 345848 39024 345900 39030
rect 345848 38966 345900 38972
rect 346308 39024 346360 39030
rect 346308 38966 346360 38972
rect 346952 39024 347004 39030
rect 346952 38966 347004 38972
rect 347688 39024 347740 39030
rect 347688 38966 347740 38972
rect 347964 39024 348016 39030
rect 347964 38966 348016 38972
rect 348976 39024 349028 39030
rect 348976 38966 349028 38972
rect 344928 3868 344980 3874
rect 344928 3810 344980 3816
rect 342076 3528 342128 3534
rect 342076 3470 342128 3476
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 343364 3324 343416 3330
rect 343364 3266 343416 3272
rect 342168 3256 342220 3262
rect 342168 3198 342220 3204
rect 342180 480 342208 3198
rect 343376 480 343404 3266
rect 344572 480 344600 3334
rect 346320 3058 346348 38966
rect 346952 4072 347004 4078
rect 346952 4014 347004 4020
rect 345756 3052 345808 3058
rect 345756 2994 345808 3000
rect 346308 3052 346360 3058
rect 346308 2994 346360 3000
rect 345768 480 345796 2994
rect 346964 480 346992 4014
rect 347700 3398 347728 38966
rect 348988 4146 349016 38966
rect 348976 4140 349028 4146
rect 348976 4082 349028 4088
rect 348056 3528 348108 3534
rect 348056 3470 348108 3476
rect 347688 3392 347740 3398
rect 347688 3334 347740 3340
rect 348068 480 348096 3470
rect 349080 3126 349108 41806
rect 349252 39364 349304 39370
rect 349252 39306 349304 39312
rect 349264 16574 349292 39306
rect 350000 39030 350028 41806
rect 351012 39030 351040 41806
rect 352024 39030 352052 41806
rect 349988 39024 350040 39030
rect 349988 38966 350040 38972
rect 350448 39024 350500 39030
rect 350448 38966 350500 38972
rect 351000 39024 351052 39030
rect 351000 38966 351052 38972
rect 351828 39024 351880 39030
rect 351828 38966 351880 38972
rect 352012 39024 352064 39030
rect 352012 38966 352064 38972
rect 349264 16546 350396 16574
rect 349252 3936 349304 3942
rect 349252 3878 349304 3884
rect 349068 3120 349120 3126
rect 349068 3062 349120 3068
rect 349264 480 349292 3878
rect 350368 3346 350396 16546
rect 350460 3534 350488 38966
rect 351840 3874 351868 38966
rect 351644 3868 351696 3874
rect 351644 3810 351696 3816
rect 351828 3868 351880 3874
rect 351828 3810 351880 3816
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 350368 3318 350488 3346
rect 350460 480 350488 3318
rect 351656 480 351684 3810
rect 353128 3466 353156 41806
rect 354048 39030 354076 41806
rect 355060 39030 355088 41806
rect 356072 39030 356100 41806
rect 353208 39024 353260 39030
rect 353208 38966 353260 38972
rect 354036 39024 354088 39030
rect 354036 38966 354088 38972
rect 354588 39024 354640 39030
rect 354588 38966 354640 38972
rect 355048 39024 355100 39030
rect 355048 38966 355100 38972
rect 355968 39024 356020 39030
rect 355968 38966 356020 38972
rect 356060 39024 356112 39030
rect 356060 38966 356112 38972
rect 353220 3806 353248 38966
rect 353208 3800 353260 3806
rect 353208 3742 353260 3748
rect 354600 3738 354628 38966
rect 355232 4140 355284 4146
rect 355232 4082 355284 4088
rect 354588 3732 354640 3738
rect 354588 3674 354640 3680
rect 353116 3460 353168 3466
rect 353116 3402 353168 3408
rect 354036 3392 354088 3398
rect 354036 3334 354088 3340
rect 352840 3052 352892 3058
rect 352840 2994 352892 3000
rect 352852 480 352880 2994
rect 354048 480 354076 3334
rect 355244 480 355272 4082
rect 355980 3058 356008 38966
rect 357268 3602 357296 41806
rect 358096 39030 358124 41806
rect 359108 39030 359136 41806
rect 360028 41806 360102 41834
rect 361086 41834 361114 42092
rect 362190 41834 362218 42092
rect 363202 41834 363230 42092
rect 364214 41834 364242 42092
rect 361086 41806 361528 41834
rect 362190 41806 362264 41834
rect 363202 41806 363276 41834
rect 357348 39024 357400 39030
rect 357348 38966 357400 38972
rect 358084 39024 358136 39030
rect 358084 38966 358136 38972
rect 358728 39024 358780 39030
rect 358728 38966 358780 38972
rect 359096 39024 359148 39030
rect 359096 38966 359148 38972
rect 357360 3942 357388 38966
rect 358740 4146 358768 38966
rect 358728 4140 358780 4146
rect 358728 4082 358780 4088
rect 357348 3936 357400 3942
rect 357348 3878 357400 3884
rect 358728 3868 358780 3874
rect 358728 3810 358780 3816
rect 357256 3596 357308 3602
rect 357256 3538 357308 3544
rect 357532 3528 357584 3534
rect 357532 3470 357584 3476
rect 356336 3120 356388 3126
rect 356336 3062 356388 3068
rect 355968 3052 356020 3058
rect 355968 2994 356020 3000
rect 356348 480 356376 3062
rect 357544 480 357572 3470
rect 358740 480 358768 3810
rect 359924 3800 359976 3806
rect 359924 3742 359976 3748
rect 359936 480 359964 3742
rect 360028 3534 360056 41806
rect 360108 39024 360160 39030
rect 360108 38966 360160 38972
rect 360120 3806 360148 38966
rect 361500 4078 361528 41806
rect 362236 38826 362264 41806
rect 363248 39030 363276 41806
rect 364168 41806 364242 41834
rect 365226 41834 365254 42092
rect 366238 41834 366266 42092
rect 367250 41834 367278 42092
rect 368262 41834 368290 42092
rect 369274 41834 369302 42092
rect 370286 41834 370314 42092
rect 371298 41834 371326 42092
rect 372310 41834 372338 42092
rect 373322 41834 373350 42092
rect 374334 41834 374362 42092
rect 375346 41834 375374 42092
rect 376358 41834 376386 42092
rect 377462 41834 377490 42092
rect 378474 41834 378502 42092
rect 379486 41834 379514 42092
rect 380498 41834 380526 42092
rect 381510 41834 381538 42092
rect 382522 41834 382550 42092
rect 383534 41834 383562 42092
rect 384546 41834 384574 42092
rect 385558 41834 385586 42092
rect 386570 41834 386598 42092
rect 387582 41834 387610 42092
rect 388594 41834 388622 42092
rect 389606 41834 389634 42092
rect 390618 41834 390646 42092
rect 391630 41834 391658 42092
rect 392734 41834 392762 42092
rect 393746 41834 393774 42092
rect 394758 41834 394786 42092
rect 395770 41834 395798 42092
rect 396782 41834 396810 42092
rect 397794 41834 397822 42092
rect 398806 41834 398834 42092
rect 399818 41834 399846 42092
rect 400830 41834 400858 42092
rect 401842 41834 401870 42092
rect 402854 41834 402882 42092
rect 365226 41806 365668 41834
rect 366238 41806 366312 41834
rect 367250 41806 367324 41834
rect 368262 41806 368428 41834
rect 369274 41806 369348 41834
rect 370286 41806 370360 41834
rect 371298 41806 371372 41834
rect 372310 41806 372476 41834
rect 373322 41806 373396 41834
rect 374334 41806 374408 41834
rect 375346 41806 375420 41834
rect 376358 41806 376708 41834
rect 377462 41806 377536 41834
rect 378474 41806 378548 41834
rect 379486 41806 379560 41834
rect 380498 41806 380848 41834
rect 381510 41806 381584 41834
rect 382522 41806 382596 41834
rect 383534 41806 383608 41834
rect 384546 41806 384988 41834
rect 385558 41806 385632 41834
rect 386570 41806 386644 41834
rect 387582 41806 387656 41834
rect 388594 41806 388668 41834
rect 389606 41806 389680 41834
rect 390618 41806 390692 41834
rect 391630 41806 391888 41834
rect 392734 41806 392808 41834
rect 393746 41806 393820 41834
rect 394758 41806 394832 41834
rect 395770 41806 396028 41834
rect 396782 41806 396856 41834
rect 397794 41806 397868 41834
rect 398806 41806 398880 41834
rect 399818 41806 400076 41834
rect 400830 41806 400904 41834
rect 401842 41806 401916 41834
rect 363236 39024 363288 39030
rect 363236 38966 363288 38972
rect 362224 38820 362276 38826
rect 362224 38762 362276 38768
rect 362868 38820 362920 38826
rect 362868 38762 362920 38768
rect 361488 4072 361540 4078
rect 361488 4014 361540 4020
rect 362880 3874 362908 38762
rect 362868 3868 362920 3874
rect 362868 3810 362920 3816
rect 360108 3800 360160 3806
rect 360108 3742 360160 3748
rect 362316 3732 362368 3738
rect 362316 3674 362368 3680
rect 360016 3528 360068 3534
rect 360016 3470 360068 3476
rect 361120 3460 361172 3466
rect 361120 3402 361172 3408
rect 361132 480 361160 3402
rect 362328 480 362356 3674
rect 364168 3466 364196 41806
rect 364248 39024 364300 39030
rect 364248 38966 364300 38972
rect 364260 3670 364288 38966
rect 364616 3936 364668 3942
rect 364616 3878 364668 3884
rect 364248 3664 364300 3670
rect 364248 3606 364300 3612
rect 364156 3460 364208 3466
rect 364156 3402 364208 3408
rect 363512 3052 363564 3058
rect 363512 2994 363564 3000
rect 363524 480 363552 2994
rect 364628 480 364656 3878
rect 365640 3738 365668 41806
rect 366284 39030 366312 41806
rect 367296 39030 367324 41806
rect 366272 39024 366324 39030
rect 366272 38966 366324 38972
rect 367008 39024 367060 39030
rect 367008 38966 367060 38972
rect 367284 39024 367336 39030
rect 367284 38966 367336 38972
rect 368296 39024 368348 39030
rect 368296 38966 368348 38972
rect 367020 6914 367048 38966
rect 366928 6886 367048 6914
rect 365628 3732 365680 3738
rect 365628 3674 365680 3680
rect 366928 3602 366956 6886
rect 367008 4140 367060 4146
rect 367008 4082 367060 4088
rect 365812 3596 365864 3602
rect 365812 3538 365864 3544
rect 366916 3596 366968 3602
rect 366916 3538 366968 3544
rect 365824 480 365852 3538
rect 367020 480 367048 4082
rect 368308 4010 368336 38966
rect 368296 4004 368348 4010
rect 368296 3946 368348 3952
rect 368400 3806 368428 41806
rect 369320 39030 369348 41806
rect 370332 39030 370360 41806
rect 371344 39030 371372 41806
rect 369308 39024 369360 39030
rect 369308 38966 369360 38972
rect 369768 39024 369820 39030
rect 369768 38966 369820 38972
rect 370320 39024 370372 39030
rect 370320 38966 370372 38972
rect 371148 39024 371200 39030
rect 371148 38966 371200 38972
rect 371332 39024 371384 39030
rect 371332 38966 371384 38972
rect 369780 3942 369808 38966
rect 370596 4072 370648 4078
rect 370596 4014 370648 4020
rect 369768 3936 369820 3942
rect 369768 3878 369820 3884
rect 368204 3800 368256 3806
rect 368204 3742 368256 3748
rect 368388 3800 368440 3806
rect 368388 3742 368440 3748
rect 368216 480 368244 3742
rect 369400 3528 369452 3534
rect 369400 3470 369452 3476
rect 369412 480 369440 3470
rect 370608 480 370636 4014
rect 371160 3398 371188 38966
rect 371700 3868 371752 3874
rect 371700 3810 371752 3816
rect 371148 3392 371200 3398
rect 371148 3334 371200 3340
rect 371712 480 371740 3810
rect 372448 3534 372476 41806
rect 373368 39030 373396 41806
rect 374380 39030 374408 41806
rect 372528 39024 372580 39030
rect 372528 38966 372580 38972
rect 373356 39024 373408 39030
rect 373356 38966 373408 38972
rect 373908 39024 373960 39030
rect 373908 38966 373960 38972
rect 374368 39024 374420 39030
rect 374368 38966 374420 38972
rect 375288 39024 375340 39030
rect 375288 38966 375340 38972
rect 372540 3874 372568 38966
rect 372528 3868 372580 3874
rect 372528 3810 372580 3816
rect 373920 3670 373948 38966
rect 375300 6914 375328 38966
rect 375392 38826 375420 41806
rect 375380 38820 375432 38826
rect 375380 38762 375432 38768
rect 376576 38820 376628 38826
rect 376576 38762 376628 38768
rect 375208 6886 375328 6914
rect 372896 3664 372948 3670
rect 372896 3606 372948 3612
rect 373908 3664 373960 3670
rect 373908 3606 373960 3612
rect 372436 3528 372488 3534
rect 372436 3470 372488 3476
rect 372908 480 372936 3606
rect 374092 3460 374144 3466
rect 374092 3402 374144 3408
rect 374104 480 374132 3402
rect 375208 3330 375236 6886
rect 375288 3732 375340 3738
rect 375288 3674 375340 3680
rect 375196 3324 375248 3330
rect 375196 3266 375248 3272
rect 375300 480 375328 3674
rect 376588 3602 376616 38762
rect 376680 3738 376708 41806
rect 377508 39030 377536 41806
rect 378520 39030 378548 41806
rect 379532 39030 379560 41806
rect 377496 39024 377548 39030
rect 377496 38966 377548 38972
rect 378048 39024 378100 39030
rect 378048 38966 378100 38972
rect 378508 39024 378560 39030
rect 378508 38966 378560 38972
rect 379428 39024 379480 39030
rect 379428 38966 379480 38972
rect 379520 39024 379572 39030
rect 379520 38966 379572 38972
rect 380716 39024 380768 39030
rect 380716 38966 380768 38972
rect 377680 4004 377732 4010
rect 377680 3946 377732 3952
rect 376668 3732 376720 3738
rect 376668 3674 376720 3680
rect 376484 3596 376536 3602
rect 376484 3538 376536 3544
rect 376576 3596 376628 3602
rect 376576 3538 376628 3544
rect 376496 480 376524 3538
rect 377692 480 377720 3946
rect 378060 3466 378088 38966
rect 379440 4010 379468 38966
rect 380728 4146 380756 38966
rect 380716 4140 380768 4146
rect 380716 4082 380768 4088
rect 380820 4078 380848 41806
rect 381556 38826 381584 41806
rect 382568 39030 382596 41806
rect 382556 39024 382608 39030
rect 382556 38966 382608 38972
rect 383476 39024 383528 39030
rect 383476 38966 383528 38972
rect 381544 38820 381596 38826
rect 381544 38762 381596 38768
rect 382188 38820 382240 38826
rect 382188 38762 382240 38768
rect 380808 4072 380860 4078
rect 380808 4014 380860 4020
rect 379428 4004 379480 4010
rect 379428 3946 379480 3952
rect 382200 3942 382228 38762
rect 379980 3936 380032 3942
rect 379980 3878 380032 3884
rect 382188 3936 382240 3942
rect 382188 3878 382240 3884
rect 378876 3800 378928 3806
rect 378876 3742 378928 3748
rect 378048 3460 378100 3466
rect 378048 3402 378100 3408
rect 378888 480 378916 3742
rect 379992 480 380020 3878
rect 382372 3868 382424 3874
rect 382372 3810 382424 3816
rect 381176 3392 381228 3398
rect 381176 3334 381228 3340
rect 381188 480 381216 3334
rect 382384 480 382412 3810
rect 383488 3806 383516 38966
rect 383580 3874 383608 41806
rect 383568 3868 383620 3874
rect 383568 3810 383620 3816
rect 383476 3800 383528 3806
rect 383476 3742 383528 3748
rect 384764 3664 384816 3670
rect 384764 3606 384816 3612
rect 383568 3528 383620 3534
rect 383568 3470 383620 3476
rect 383580 480 383608 3470
rect 384776 480 384804 3606
rect 384960 3534 384988 41806
rect 385604 39030 385632 41806
rect 386616 39030 386644 41806
rect 385592 39024 385644 39030
rect 385592 38966 385644 38972
rect 386328 39024 386380 39030
rect 386328 38966 386380 38972
rect 386604 39024 386656 39030
rect 386604 38966 386656 38972
rect 386340 3670 386368 38966
rect 386328 3664 386380 3670
rect 386328 3606 386380 3612
rect 387628 3602 387656 41806
rect 388640 39030 388668 41806
rect 389652 39030 389680 41806
rect 390664 39030 390692 41806
rect 387708 39024 387760 39030
rect 387708 38966 387760 38972
rect 388628 39024 388680 39030
rect 388628 38966 388680 38972
rect 389088 39024 389140 39030
rect 389088 38966 389140 38972
rect 389640 39024 389692 39030
rect 389640 38966 389692 38972
rect 390468 39024 390520 39030
rect 390468 38966 390520 38972
rect 390652 39024 390704 39030
rect 390652 38966 390704 38972
rect 391756 39024 391808 39030
rect 391756 38966 391808 38972
rect 387156 3596 387208 3602
rect 387156 3538 387208 3544
rect 387616 3596 387668 3602
rect 387616 3538 387668 3544
rect 384948 3528 385000 3534
rect 384948 3470 385000 3476
rect 385960 3324 386012 3330
rect 385960 3266 386012 3272
rect 385972 480 386000 3266
rect 387168 480 387196 3538
rect 387720 3398 387748 38966
rect 388260 3732 388312 3738
rect 388260 3674 388312 3680
rect 387708 3392 387760 3398
rect 387708 3334 387760 3340
rect 388272 480 388300 3674
rect 389100 3330 389128 38966
rect 389456 3460 389508 3466
rect 389456 3402 389508 3408
rect 389088 3324 389140 3330
rect 389088 3266 389140 3272
rect 389468 480 389496 3402
rect 390480 3262 390508 38966
rect 391664 4140 391716 4146
rect 391664 4082 391716 4088
rect 390652 4004 390704 4010
rect 390652 3946 390704 3952
rect 390468 3256 390520 3262
rect 390468 3198 390520 3204
rect 390664 480 390692 3946
rect 391676 2122 391704 4082
rect 391768 4010 391796 38966
rect 391756 4004 391808 4010
rect 391756 3946 391808 3952
rect 391860 3466 391888 41806
rect 392780 39030 392808 41806
rect 393792 39030 393820 41806
rect 392768 39024 392820 39030
rect 392768 38966 392820 38972
rect 393228 39024 393280 39030
rect 393228 38966 393280 38972
rect 393780 39024 393832 39030
rect 393780 38966 393832 38972
rect 394608 39024 394660 39030
rect 394608 38966 394660 38972
rect 393044 4072 393096 4078
rect 393044 4014 393096 4020
rect 391848 3460 391900 3466
rect 391848 3402 391900 3408
rect 391676 2094 391888 2122
rect 391860 480 391888 2094
rect 393056 480 393084 4014
rect 393240 3738 393268 38966
rect 394240 3936 394292 3942
rect 394240 3878 394292 3884
rect 393228 3732 393280 3738
rect 393228 3674 393280 3680
rect 394252 480 394280 3878
rect 394620 3126 394648 38966
rect 394804 38962 394832 41806
rect 394792 38956 394844 38962
rect 394792 38898 394844 38904
rect 395896 38956 395948 38962
rect 395896 38898 395948 38904
rect 395908 4078 395936 38898
rect 395896 4072 395948 4078
rect 395896 4014 395948 4020
rect 396000 3806 396028 41806
rect 396828 39030 396856 41806
rect 397840 39030 397868 41806
rect 398852 39030 398880 41806
rect 396816 39024 396868 39030
rect 396816 38966 396868 38972
rect 397368 39024 397420 39030
rect 397368 38966 397420 38972
rect 397828 39024 397880 39030
rect 397828 38966 397880 38972
rect 398748 39024 398800 39030
rect 398748 38966 398800 38972
rect 398840 39024 398892 39030
rect 398840 38966 398892 38972
rect 397380 3942 397408 38966
rect 398760 4146 398788 38966
rect 398748 4140 398800 4146
rect 398748 4082 398800 4088
rect 397368 3936 397420 3942
rect 397368 3878 397420 3884
rect 396540 3868 396592 3874
rect 396540 3810 396592 3816
rect 395344 3800 395396 3806
rect 395344 3742 395396 3748
rect 395988 3800 396040 3806
rect 395988 3742 396040 3748
rect 394608 3120 394660 3126
rect 394608 3062 394660 3068
rect 395356 480 395384 3742
rect 396552 480 396580 3810
rect 398932 3664 398984 3670
rect 398932 3606 398984 3612
rect 397736 3528 397788 3534
rect 397736 3470 397788 3476
rect 397748 480 397776 3470
rect 398944 480 398972 3606
rect 400048 3534 400076 41806
rect 400128 39024 400180 39030
rect 400128 38966 400180 38972
rect 400036 3528 400088 3534
rect 400036 3470 400088 3476
rect 400140 3482 400168 38966
rect 400876 38826 400904 41806
rect 401888 39030 401916 41806
rect 402808 41806 402882 41834
rect 403866 41834 403894 42092
rect 404878 41834 404906 42092
rect 405890 41834 405918 42092
rect 406902 41834 406930 42092
rect 408006 41834 408034 42092
rect 409018 41834 409046 42092
rect 410030 41834 410058 42092
rect 411042 41834 411070 42092
rect 412054 41834 412082 42092
rect 413066 41834 413094 42092
rect 414078 41834 414106 42092
rect 415090 41834 415118 42092
rect 416102 41834 416130 42092
rect 417114 41834 417142 42092
rect 418126 41834 418154 42092
rect 419138 41834 419166 42092
rect 420150 41834 420178 42092
rect 421162 41834 421190 42092
rect 422174 41834 422202 42092
rect 403866 41806 404308 41834
rect 404878 41806 404952 41834
rect 405890 41806 405964 41834
rect 406902 41806 406976 41834
rect 408006 41806 408448 41834
rect 409018 41806 409092 41834
rect 410030 41806 410104 41834
rect 411042 41806 411208 41834
rect 412054 41806 412128 41834
rect 413066 41806 413140 41834
rect 414078 41806 414152 41834
rect 415090 41806 415256 41834
rect 416102 41806 416176 41834
rect 417114 41806 417188 41834
rect 418126 41806 418200 41834
rect 419138 41806 419488 41834
rect 420150 41806 420224 41834
rect 421162 41806 421236 41834
rect 401876 39024 401928 39030
rect 401876 38966 401928 38972
rect 400864 38820 400916 38826
rect 400864 38762 400916 38768
rect 401508 38820 401560 38826
rect 401508 38762 401560 38768
rect 401520 3874 401548 38762
rect 401508 3868 401560 3874
rect 401508 3810 401560 3816
rect 402808 3602 402836 41806
rect 402888 39024 402940 39030
rect 402888 38966 402940 38972
rect 401324 3596 401376 3602
rect 401324 3538 401376 3544
rect 402796 3596 402848 3602
rect 402796 3538 402848 3544
rect 400140 3454 400260 3482
rect 400232 3398 400260 3454
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400220 3392 400272 3398
rect 400220 3334 400272 3340
rect 400140 480 400168 3334
rect 401336 480 401364 3538
rect 402900 3330 402928 38966
rect 404280 3670 404308 41806
rect 404924 39030 404952 41806
rect 405936 39030 405964 41806
rect 404912 39024 404964 39030
rect 404912 38966 404964 38972
rect 405648 39024 405700 39030
rect 405648 38966 405700 38972
rect 405924 39024 405976 39030
rect 405924 38966 405976 38972
rect 405660 4010 405688 38966
rect 404820 4004 404872 4010
rect 404820 3946 404872 3952
rect 405648 4004 405700 4010
rect 405648 3946 405700 3952
rect 404268 3664 404320 3670
rect 404268 3606 404320 3612
rect 402520 3324 402572 3330
rect 402520 3266 402572 3272
rect 402888 3324 402940 3330
rect 402888 3266 402940 3272
rect 402532 480 402560 3266
rect 403624 3256 403676 3262
rect 403624 3198 403676 3204
rect 403636 480 403664 3198
rect 404832 480 404860 3946
rect 406948 3466 406976 41806
rect 407028 39024 407080 39030
rect 407028 38966 407080 38972
rect 406016 3460 406068 3466
rect 406016 3402 406068 3408
rect 406936 3460 406988 3466
rect 406936 3402 406988 3408
rect 406028 480 406056 3402
rect 407040 3194 407068 38966
rect 408420 6914 408448 41806
rect 409064 39030 409092 41806
rect 410076 39030 410104 41806
rect 409052 39024 409104 39030
rect 409052 38966 409104 38972
rect 409788 39024 409840 39030
rect 409788 38966 409840 38972
rect 410064 39024 410116 39030
rect 410064 38966 410116 38972
rect 411076 39024 411128 39030
rect 411076 38966 411128 38972
rect 408328 6886 408448 6914
rect 407212 3732 407264 3738
rect 407212 3674 407264 3680
rect 407028 3188 407080 3194
rect 407028 3130 407080 3136
rect 407224 480 407252 3674
rect 408328 2922 408356 6886
rect 409604 4072 409656 4078
rect 409604 4014 409656 4020
rect 408408 3120 408460 3126
rect 408408 3062 408460 3068
rect 408316 2916 408368 2922
rect 408316 2858 408368 2864
rect 408420 480 408448 3062
rect 409616 480 409644 4014
rect 409800 2990 409828 38966
rect 410800 3800 410852 3806
rect 410800 3742 410852 3748
rect 409788 2984 409840 2990
rect 409788 2926 409840 2932
rect 410812 480 410840 3742
rect 411088 3738 411116 38966
rect 411180 4078 411208 41806
rect 412100 39030 412128 41806
rect 413112 39030 413140 41806
rect 414124 39030 414152 41806
rect 412088 39024 412140 39030
rect 412088 38966 412140 38972
rect 412548 39024 412600 39030
rect 412548 38966 412600 38972
rect 413100 39024 413152 39030
rect 413100 38966 413152 38972
rect 413928 39024 413980 39030
rect 413928 38966 413980 38972
rect 414112 39024 414164 39030
rect 414112 38966 414164 38972
rect 411168 4072 411220 4078
rect 411168 4014 411220 4020
rect 411904 3936 411956 3942
rect 411904 3878 411956 3884
rect 411076 3732 411128 3738
rect 411076 3674 411128 3680
rect 411916 480 411944 3878
rect 412560 3262 412588 38966
rect 413940 4146 413968 38966
rect 413100 4140 413152 4146
rect 413100 4082 413152 4088
rect 413928 4140 413980 4146
rect 413928 4082 413980 4088
rect 412548 3256 412600 3262
rect 412548 3198 412600 3204
rect 413112 480 413140 4082
rect 415228 3806 415256 41806
rect 416148 39030 416176 41806
rect 417160 39030 417188 41806
rect 418172 39030 418200 41806
rect 415308 39024 415360 39030
rect 415308 38966 415360 38972
rect 416136 39024 416188 39030
rect 416136 38966 416188 38972
rect 416688 39024 416740 39030
rect 416688 38966 416740 38972
rect 417148 39024 417200 39030
rect 417148 38966 417200 38972
rect 418068 39024 418120 39030
rect 418068 38966 418120 38972
rect 418160 39024 418212 39030
rect 418160 38966 418212 38972
rect 419356 39024 419408 39030
rect 419356 38966 419408 38972
rect 415216 3800 415268 3806
rect 415216 3742 415268 3748
rect 415320 3398 415348 38966
rect 416700 6914 416728 38966
rect 416608 6886 416728 6914
rect 415492 3528 415544 3534
rect 415492 3470 415544 3476
rect 414296 3392 414348 3398
rect 414296 3334 414348 3340
rect 415308 3392 415360 3398
rect 415308 3334 415360 3340
rect 414308 480 414336 3334
rect 415504 480 415532 3470
rect 416608 3058 416636 6886
rect 416688 3868 416740 3874
rect 416688 3810 416740 3816
rect 416596 3052 416648 3058
rect 416596 2994 416648 3000
rect 416700 480 416728 3810
rect 418080 3330 418108 38966
rect 419368 3942 419396 38966
rect 419356 3936 419408 3942
rect 419356 3878 419408 3884
rect 419460 3602 419488 41806
rect 420196 38826 420224 41806
rect 421208 39030 421236 41806
rect 422128 41806 422202 41834
rect 423278 41834 423306 42092
rect 424290 41834 424318 42092
rect 425302 41834 425330 42092
rect 426314 41834 426342 42092
rect 427326 41834 427354 42092
rect 428338 41834 428366 42092
rect 429350 41834 429378 42092
rect 430362 41834 430390 42092
rect 431374 41834 431402 42092
rect 432386 41834 432414 42092
rect 433398 41834 433426 42092
rect 434410 41834 434438 42092
rect 435422 41834 435450 42092
rect 436434 41834 436462 42092
rect 437446 41834 437474 42092
rect 438550 41834 438578 42092
rect 439562 41834 439590 42092
rect 440574 41834 440602 42092
rect 441586 41834 441614 42092
rect 442598 41834 442626 42092
rect 443610 41834 443638 42092
rect 444622 41834 444650 42092
rect 445634 41834 445662 42092
rect 423278 41806 423628 41834
rect 424290 41806 424364 41834
rect 425302 41806 425376 41834
rect 426314 41806 426388 41834
rect 427326 41806 427768 41834
rect 428338 41806 428412 41834
rect 429350 41806 429424 41834
rect 430362 41806 430436 41834
rect 431374 41806 431448 41834
rect 432386 41806 432460 41834
rect 433398 41806 433472 41834
rect 434410 41806 434484 41834
rect 435422 41806 435496 41834
rect 436434 41806 436508 41834
rect 437446 41806 437520 41834
rect 438550 41806 438808 41834
rect 439562 41806 439636 41834
rect 440574 41806 440648 41834
rect 441586 41806 441660 41834
rect 442598 41806 442856 41834
rect 443610 41806 443684 41834
rect 444622 41806 444696 41834
rect 421196 39024 421248 39030
rect 421196 38966 421248 38972
rect 420184 38820 420236 38826
rect 420184 38762 420236 38768
rect 420828 38820 420880 38826
rect 420828 38762 420880 38768
rect 420840 3874 420868 38762
rect 421380 4004 421432 4010
rect 421380 3946 421432 3952
rect 420828 3868 420880 3874
rect 420828 3810 420880 3816
rect 420184 3664 420236 3670
rect 420184 3606 420236 3612
rect 418988 3596 419040 3602
rect 418988 3538 419040 3544
rect 419448 3596 419500 3602
rect 419448 3538 419500 3544
rect 417884 3324 417936 3330
rect 417884 3266 417936 3272
rect 418068 3324 418120 3330
rect 418068 3266 418120 3272
rect 417896 480 417924 3266
rect 419000 480 419028 3538
rect 420196 480 420224 3606
rect 421392 480 421420 3946
rect 422128 3534 422156 41806
rect 422208 39024 422260 39030
rect 422208 38966 422260 38972
rect 422220 4010 422248 38966
rect 422208 4004 422260 4010
rect 422208 3946 422260 3952
rect 422116 3528 422168 3534
rect 422116 3470 422168 3476
rect 422576 3188 422628 3194
rect 422576 3130 422628 3136
rect 422588 480 422616 3130
rect 423600 3126 423628 41806
rect 424336 39030 424364 41806
rect 425348 39030 425376 41806
rect 424324 39024 424376 39030
rect 424324 38966 424376 38972
rect 424968 39024 425020 39030
rect 424968 38966 425020 38972
rect 425336 39024 425388 39030
rect 425336 38966 425388 38972
rect 426256 39024 426308 39030
rect 426256 38966 426308 38972
rect 423772 3460 423824 3466
rect 423772 3402 423824 3408
rect 423588 3120 423640 3126
rect 423588 3062 423640 3068
rect 423784 480 423812 3402
rect 424980 3194 425008 38966
rect 426268 3670 426296 38966
rect 426256 3664 426308 3670
rect 426256 3606 426308 3612
rect 426360 3466 426388 41806
rect 427740 3738 427768 41806
rect 428384 39030 428412 41806
rect 429396 39030 429424 41806
rect 428372 39024 428424 39030
rect 428372 38966 428424 38972
rect 429108 39024 429160 39030
rect 429108 38966 429160 38972
rect 429384 39024 429436 39030
rect 429384 38966 429436 38972
rect 429120 4894 429148 38966
rect 429108 4888 429160 4894
rect 429108 4830 429160 4836
rect 430408 4078 430436 41806
rect 431420 39030 431448 41806
rect 432432 39030 432460 41806
rect 433444 39030 433472 41806
rect 434456 39438 434484 41806
rect 434444 39432 434496 39438
rect 434444 39374 434496 39380
rect 435468 39030 435496 41806
rect 436480 39030 436508 41806
rect 437492 39370 437520 41806
rect 437480 39364 437532 39370
rect 437480 39306 437532 39312
rect 430488 39024 430540 39030
rect 430488 38966 430540 38972
rect 431408 39024 431460 39030
rect 431408 38966 431460 38972
rect 431868 39024 431920 39030
rect 431868 38966 431920 38972
rect 432420 39024 432472 39030
rect 432420 38966 432472 38972
rect 433248 39024 433300 39030
rect 433248 38966 433300 38972
rect 433432 39024 433484 39030
rect 433432 38966 433484 38972
rect 434628 39024 434680 39030
rect 434628 38966 434680 38972
rect 435456 39024 435508 39030
rect 435456 38966 435508 38972
rect 436008 39024 436060 39030
rect 436008 38966 436060 38972
rect 436468 39024 436520 39030
rect 436468 38966 436520 38972
rect 437388 39024 437440 39030
rect 437388 38966 437440 38972
rect 428464 4072 428516 4078
rect 428464 4014 428516 4020
rect 430396 4072 430448 4078
rect 430396 4014 430448 4020
rect 427268 3732 427320 3738
rect 427268 3674 427320 3680
rect 427728 3732 427780 3738
rect 427728 3674 427780 3680
rect 426348 3460 426400 3466
rect 426348 3402 426400 3408
rect 424968 3188 425020 3194
rect 424968 3130 425020 3136
rect 426164 2984 426216 2990
rect 426164 2926 426216 2932
rect 424968 2916 425020 2922
rect 424968 2858 425020 2864
rect 424980 480 425008 2858
rect 426176 480 426204 2926
rect 427280 480 427308 3674
rect 428476 480 428504 4014
rect 430500 3262 430528 38966
rect 431880 4826 431908 38966
rect 431868 4820 431920 4826
rect 431868 4762 431920 4768
rect 433260 4146 433288 38966
rect 430856 4140 430908 4146
rect 430856 4082 430908 4088
rect 433248 4140 433300 4146
rect 433248 4082 433300 4088
rect 429660 3256 429712 3262
rect 429660 3198 429712 3204
rect 430488 3256 430540 3262
rect 430488 3198 430540 3204
rect 429672 480 429700 3198
rect 430868 480 430896 4082
rect 433248 3800 433300 3806
rect 433248 3742 433300 3748
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 432064 480 432092 3334
rect 433260 480 433288 3742
rect 434444 3052 434496 3058
rect 434444 2994 434496 3000
rect 434456 480 434484 2994
rect 434640 2990 434668 38966
rect 436020 3806 436048 38966
rect 436744 3936 436796 3942
rect 436744 3878 436796 3884
rect 436008 3800 436060 3806
rect 436008 3742 436060 3748
rect 435548 3324 435600 3330
rect 435548 3266 435600 3272
rect 434628 2984 434680 2990
rect 434628 2926 434680 2932
rect 435560 480 435588 3266
rect 436756 480 436784 3878
rect 437400 3398 437428 38966
rect 438780 3942 438808 41806
rect 439608 39030 439636 41806
rect 440620 39030 440648 41806
rect 441632 39030 441660 41806
rect 439596 39024 439648 39030
rect 439596 38966 439648 38972
rect 440148 39024 440200 39030
rect 440148 38966 440200 38972
rect 440608 39024 440660 39030
rect 440608 38966 440660 38972
rect 441528 39024 441580 39030
rect 441528 38966 441580 38972
rect 441620 39024 441672 39030
rect 441620 38966 441672 38972
rect 438768 3936 438820 3942
rect 438768 3878 438820 3884
rect 439136 3868 439188 3874
rect 439136 3810 439188 3816
rect 437940 3596 437992 3602
rect 437940 3538 437992 3544
rect 437388 3392 437440 3398
rect 437388 3334 437440 3340
rect 437952 480 437980 3538
rect 439148 480 439176 3810
rect 440160 3330 440188 38966
rect 441540 4010 441568 38966
rect 440332 4004 440384 4010
rect 440332 3946 440384 3952
rect 441528 4004 441580 4010
rect 441528 3946 441580 3952
rect 440148 3324 440200 3330
rect 440148 3266 440200 3272
rect 440344 480 440372 3946
rect 442828 3602 442856 41806
rect 443552 39432 443604 39438
rect 443552 39374 443604 39380
rect 442908 39024 442960 39030
rect 442908 38966 442960 38972
rect 442920 3874 442948 38966
rect 443564 35894 443592 39374
rect 443656 39030 443684 41806
rect 443644 39024 443696 39030
rect 443644 38966 443696 38972
rect 444288 39024 444340 39030
rect 444288 38966 444340 38972
rect 443564 35866 443684 35894
rect 443656 4962 443684 35866
rect 443644 4956 443696 4962
rect 443644 4898 443696 4904
rect 442908 3868 442960 3874
rect 442908 3810 442960 3816
rect 442816 3596 442868 3602
rect 442816 3538 442868 3544
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 441540 480 441568 3470
rect 443828 3188 443880 3194
rect 443828 3130 443880 3136
rect 442632 3120 442684 3126
rect 442632 3062 442684 3068
rect 442644 480 442672 3062
rect 443840 480 443868 3130
rect 444300 3058 444328 38966
rect 444668 38962 444696 41806
rect 445588 41806 445662 41834
rect 446646 41834 446674 42092
rect 447658 41834 447686 42092
rect 448670 41834 448698 42092
rect 449682 41834 449710 42092
rect 450694 41834 450722 42092
rect 451706 41834 451734 42092
rect 452718 41834 452746 42092
rect 453822 41834 453850 42092
rect 454834 41834 454862 42092
rect 455846 41834 455874 42092
rect 456858 41834 456886 42092
rect 457870 41834 457898 42092
rect 458882 41834 458910 42092
rect 459894 41834 459922 42092
rect 460906 41834 460934 42092
rect 461918 41834 461946 42092
rect 462930 41834 462958 42092
rect 463942 41834 463970 42092
rect 464954 41834 464982 42092
rect 465966 41834 465994 42092
rect 466978 41834 467006 42092
rect 467990 41834 468018 42092
rect 469094 41834 469122 42092
rect 470106 41834 470134 42092
rect 471118 41834 471146 42092
rect 472130 41834 472158 42092
rect 473142 41834 473170 42092
rect 474154 41834 474182 42092
rect 475166 41834 475194 42092
rect 476178 41834 476206 42092
rect 477190 41834 477218 42092
rect 478202 41834 478230 42092
rect 479214 41834 479242 42092
rect 480226 41834 480254 42092
rect 481238 41834 481266 42092
rect 482250 41834 482278 42092
rect 483262 41834 483290 42092
rect 484366 41834 484394 42092
rect 485378 41834 485406 42092
rect 486390 41834 486418 42092
rect 487402 41834 487430 42092
rect 488414 41834 488442 42092
rect 489426 41834 489454 42092
rect 490438 41834 490466 42092
rect 491450 41834 491478 42092
rect 492462 41834 492490 42092
rect 493474 41834 493502 42092
rect 494486 41834 494514 42092
rect 495498 41834 495526 42092
rect 496510 41834 496538 42092
rect 497522 41834 497550 42092
rect 498534 41834 498562 42092
rect 499638 41834 499666 42092
rect 500650 41834 500678 42092
rect 501662 41834 501690 42092
rect 502674 41834 502702 42092
rect 503686 41834 503714 42092
rect 504698 41834 504726 42092
rect 505710 41834 505738 42092
rect 506722 41834 506750 42092
rect 507734 41834 507762 42092
rect 446646 41806 447088 41834
rect 447658 41806 447732 41834
rect 448670 41806 448744 41834
rect 449682 41806 449756 41834
rect 450694 41806 450768 41834
rect 451706 41806 451780 41834
rect 452718 41806 452792 41834
rect 453822 41806 453988 41834
rect 454834 41806 454908 41834
rect 455846 41806 455920 41834
rect 456858 41806 456932 41834
rect 457870 41806 458128 41834
rect 458882 41806 458956 41834
rect 459894 41806 459968 41834
rect 460906 41806 460980 41834
rect 461918 41806 462176 41834
rect 462930 41806 463004 41834
rect 463942 41806 464016 41834
rect 464954 41806 465028 41834
rect 465966 41806 466408 41834
rect 466978 41806 467052 41834
rect 467990 41806 468064 41834
rect 469094 41806 469168 41834
rect 470106 41806 470548 41834
rect 471118 41806 471192 41834
rect 472130 41806 472204 41834
rect 473142 41806 473308 41834
rect 474154 41806 474228 41834
rect 475166 41806 475240 41834
rect 476178 41806 476252 41834
rect 477190 41806 477264 41834
rect 478202 41806 478276 41834
rect 479214 41806 479288 41834
rect 480226 41806 480300 41834
rect 481238 41806 481588 41834
rect 482250 41806 482324 41834
rect 483262 41806 483336 41834
rect 484366 41806 484440 41834
rect 485378 41806 485728 41834
rect 486390 41806 486464 41834
rect 487402 41806 487476 41834
rect 488414 41806 488488 41834
rect 489426 41806 489868 41834
rect 490438 41806 490512 41834
rect 491450 41806 491524 41834
rect 492462 41806 492536 41834
rect 493474 41806 493548 41834
rect 494486 41806 494560 41834
rect 495498 41806 495572 41834
rect 496510 41806 496768 41834
rect 497522 41806 497596 41834
rect 498534 41806 498608 41834
rect 499638 41806 499712 41834
rect 500650 41806 500908 41834
rect 501662 41806 501736 41834
rect 502674 41806 502748 41834
rect 503686 41806 503760 41834
rect 504698 41806 505048 41834
rect 505710 41806 505784 41834
rect 506722 41806 506796 41834
rect 444656 38956 444708 38962
rect 444656 38898 444708 38904
rect 445024 3664 445076 3670
rect 445024 3606 445076 3612
rect 444288 3052 444340 3058
rect 444288 2994 444340 3000
rect 445036 480 445064 3606
rect 445588 3534 445616 41806
rect 445668 38956 445720 38962
rect 445668 38898 445720 38904
rect 445680 3670 445708 38898
rect 445668 3664 445720 3670
rect 445668 3606 445720 3612
rect 445576 3528 445628 3534
rect 445576 3470 445628 3476
rect 446220 3460 446272 3466
rect 446220 3402 446272 3408
rect 446232 480 446260 3402
rect 447060 2854 447088 41806
rect 447704 39030 447732 41806
rect 448716 39030 448744 41806
rect 447692 39024 447744 39030
rect 447692 38966 447744 38972
rect 448428 39024 448480 39030
rect 448428 38966 448480 38972
rect 448704 39024 448756 39030
rect 448704 38966 448756 38972
rect 448440 3738 448468 38966
rect 448612 4888 448664 4894
rect 448612 4830 448664 4836
rect 447416 3732 447468 3738
rect 447416 3674 447468 3680
rect 448428 3732 448480 3738
rect 448428 3674 448480 3680
rect 447048 2848 447100 2854
rect 447048 2790 447100 2796
rect 447428 480 447456 3674
rect 448624 480 448652 4830
rect 449728 3466 449756 41806
rect 450740 39030 450768 41806
rect 451752 39030 451780 41806
rect 452764 39030 452792 41806
rect 449808 39024 449860 39030
rect 449808 38966 449860 38972
rect 450728 39024 450780 39030
rect 450728 38966 450780 38972
rect 451188 39024 451240 39030
rect 451188 38966 451240 38972
rect 451740 39024 451792 39030
rect 451740 38966 451792 38972
rect 452568 39024 452620 39030
rect 452568 38966 452620 38972
rect 452752 39024 452804 39030
rect 452752 38966 452804 38972
rect 453856 39024 453908 39030
rect 453856 38966 453908 38972
rect 449716 3460 449768 3466
rect 449716 3402 449768 3408
rect 449820 3346 449848 38966
rect 450912 4072 450964 4078
rect 450912 4014 450964 4020
rect 449728 3318 449848 3346
rect 449728 3126 449756 3318
rect 449808 3256 449860 3262
rect 449808 3198 449860 3204
rect 449716 3120 449768 3126
rect 449716 3062 449768 3068
rect 449820 480 449848 3198
rect 450924 480 450952 4014
rect 451200 3194 451228 38966
rect 452108 4820 452160 4826
rect 452108 4762 452160 4768
rect 451188 3188 451240 3194
rect 451188 3130 451240 3136
rect 452120 480 452148 4762
rect 452580 2922 452608 38966
rect 453304 4140 453356 4146
rect 453304 4082 453356 4088
rect 452568 2916 452620 2922
rect 452568 2858 452620 2864
rect 453316 480 453344 4082
rect 453868 3262 453896 38966
rect 453960 4078 453988 41806
rect 454684 39364 454736 39370
rect 454684 39306 454736 39312
rect 454696 5574 454724 39306
rect 454880 39030 454908 41806
rect 455892 39370 455920 41806
rect 455880 39364 455932 39370
rect 455880 39306 455932 39312
rect 456904 39030 456932 41806
rect 454868 39024 454920 39030
rect 454868 38966 454920 38972
rect 455328 39024 455380 39030
rect 455328 38966 455380 38972
rect 456892 39024 456944 39030
rect 456892 38966 456944 38972
rect 457996 39024 458048 39030
rect 457996 38966 458048 38972
rect 454684 5568 454736 5574
rect 454684 5510 454736 5516
rect 455340 4146 455368 38966
rect 455696 4956 455748 4962
rect 455696 4898 455748 4904
rect 455328 4140 455380 4146
rect 455328 4082 455380 4088
rect 453948 4072 454000 4078
rect 453948 4014 454000 4020
rect 453856 3256 453908 3262
rect 453856 3198 453908 3204
rect 454500 2984 454552 2990
rect 454500 2926 454552 2932
rect 454512 480 454540 2926
rect 455708 480 455736 4898
rect 458008 3806 458036 38966
rect 456892 3800 456944 3806
rect 456892 3742 456944 3748
rect 457996 3800 458048 3806
rect 457996 3742 458048 3748
rect 456904 480 456932 3742
rect 458100 3398 458128 41806
rect 458928 39438 458956 41806
rect 458916 39432 458968 39438
rect 458916 39374 458968 39380
rect 459940 39030 459968 41806
rect 460952 39030 460980 41806
rect 459928 39024 459980 39030
rect 459928 38966 459980 38972
rect 460848 39024 460900 39030
rect 460848 38966 460900 38972
rect 460940 39024 460992 39030
rect 460940 38966 460992 38972
rect 459192 5568 459244 5574
rect 459192 5510 459244 5516
rect 457996 3392 458048 3398
rect 457996 3334 458048 3340
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458008 1714 458036 3334
rect 458008 1686 458128 1714
rect 458100 480 458128 1686
rect 459204 480 459232 5510
rect 460388 3936 460440 3942
rect 460388 3878 460440 3884
rect 460400 480 460428 3878
rect 460860 2990 460888 38966
rect 462148 4962 462176 41806
rect 462976 39030 463004 41806
rect 462228 39024 462280 39030
rect 462228 38966 462280 38972
rect 462964 39024 463016 39030
rect 462964 38966 463016 38972
rect 463608 39024 463660 39030
rect 463608 38966 463660 38972
rect 462136 4956 462188 4962
rect 462136 4898 462188 4904
rect 462240 3330 462268 38966
rect 463620 4010 463648 38966
rect 463988 38962 464016 41806
rect 465000 39642 465028 41806
rect 464988 39636 465040 39642
rect 464988 39578 465040 39584
rect 465724 39364 465776 39370
rect 465724 39306 465776 39312
rect 463976 38956 464028 38962
rect 463976 38898 464028 38904
rect 464988 38956 465040 38962
rect 464988 38898 465040 38904
rect 462780 4004 462832 4010
rect 462780 3946 462832 3952
rect 463608 4004 463660 4010
rect 463608 3946 463660 3952
rect 461584 3324 461636 3330
rect 461584 3266 461636 3272
rect 462228 3324 462280 3330
rect 462228 3266 462280 3272
rect 460848 2984 460900 2990
rect 460848 2926 460900 2932
rect 461596 480 461624 3266
rect 462792 480 462820 3946
rect 465000 3942 465028 38898
rect 465736 5030 465764 39306
rect 465724 5024 465776 5030
rect 465724 4966 465776 4972
rect 464988 3936 465040 3942
rect 464988 3878 465040 3884
rect 463976 3868 464028 3874
rect 463976 3810 464028 3816
rect 463988 480 464016 3810
rect 465172 3596 465224 3602
rect 465172 3538 465224 3544
rect 465184 480 465212 3538
rect 466380 3058 466408 41806
rect 467024 39030 467052 41806
rect 468036 39030 468064 41806
rect 467012 39024 467064 39030
rect 467012 38966 467064 38972
rect 467748 39024 467800 39030
rect 467748 38966 467800 38972
rect 468024 39024 468076 39030
rect 468024 38966 468076 38972
rect 469036 39024 469088 39030
rect 469036 38966 469088 38972
rect 467760 3874 467788 38966
rect 469048 4894 469076 38966
rect 469036 4888 469088 4894
rect 469036 4830 469088 4836
rect 467748 3868 467800 3874
rect 467748 3810 467800 3816
rect 469140 3670 469168 41806
rect 467472 3664 467524 3670
rect 467472 3606 467524 3612
rect 469128 3664 469180 3670
rect 469128 3606 469180 3612
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466368 3052 466420 3058
rect 466368 2994 466420 3000
rect 466288 480 466316 2994
rect 467484 480 467512 3606
rect 470520 3534 470548 41806
rect 471164 39030 471192 41806
rect 471152 39024 471204 39030
rect 471152 38966 471204 38972
rect 471888 39024 471940 39030
rect 471888 38966 471940 38972
rect 471900 4826 471928 38966
rect 472176 38758 472204 41806
rect 472164 38752 472216 38758
rect 472164 38694 472216 38700
rect 473176 38752 473228 38758
rect 473176 38694 473228 38700
rect 471888 4820 471940 4826
rect 471888 4762 471940 4768
rect 473188 3738 473216 38694
rect 471060 3732 471112 3738
rect 471060 3674 471112 3680
rect 473176 3732 473228 3738
rect 473176 3674 473228 3680
rect 468668 3528 468720 3534
rect 468668 3470 468720 3476
rect 470508 3528 470560 3534
rect 470508 3470 470560 3476
rect 468680 480 468708 3470
rect 469864 2848 469916 2854
rect 469864 2790 469916 2796
rect 469876 480 469904 2790
rect 471072 480 471100 3674
rect 473280 3602 473308 41806
rect 474200 39370 474228 41806
rect 474188 39364 474240 39370
rect 474188 39306 474240 39312
rect 475212 39030 475240 41806
rect 476224 39030 476252 41806
rect 477236 39574 477264 41806
rect 477224 39568 477276 39574
rect 477224 39510 477276 39516
rect 478248 39030 478276 41806
rect 479260 39030 479288 41806
rect 480272 39506 480300 41806
rect 480260 39500 480312 39506
rect 480260 39442 480312 39448
rect 475200 39024 475252 39030
rect 475200 38966 475252 38972
rect 476028 39024 476080 39030
rect 476028 38966 476080 38972
rect 476212 39024 476264 39030
rect 476212 38966 476264 38972
rect 477408 39024 477460 39030
rect 477408 38966 477460 38972
rect 478236 39024 478288 39030
rect 478236 38966 478288 38972
rect 478788 39024 478840 39030
rect 478788 38966 478840 38972
rect 479248 39024 479300 39030
rect 479248 38966 479300 38972
rect 480168 39024 480220 39030
rect 480168 38966 480220 38972
rect 473268 3596 473320 3602
rect 473268 3538 473320 3544
rect 473452 3460 473504 3466
rect 473452 3402 473504 3408
rect 472256 3120 472308 3126
rect 472256 3062 472308 3068
rect 472268 480 472296 3062
rect 473464 480 473492 3402
rect 476040 3194 476068 38966
rect 477420 3466 477448 38966
rect 478144 4072 478196 4078
rect 478144 4014 478196 4020
rect 477408 3460 477460 3466
rect 477408 3402 477460 3408
rect 476948 3256 477000 3262
rect 476948 3198 477000 3204
rect 474556 3188 474608 3194
rect 474556 3130 474608 3136
rect 476028 3188 476080 3194
rect 476028 3130 476080 3136
rect 474568 480 474596 3130
rect 475752 2916 475804 2922
rect 475752 2858 475804 2864
rect 475764 480 475792 2858
rect 476960 480 476988 3198
rect 478156 480 478184 4014
rect 478800 3262 478828 38966
rect 479340 4140 479392 4146
rect 479340 4082 479392 4088
rect 478788 3256 478840 3262
rect 478788 3198 478840 3204
rect 479352 480 479380 4082
rect 480180 3126 480208 38966
rect 480536 5024 480588 5030
rect 480536 4966 480588 4972
rect 480168 3120 480220 3126
rect 480168 3062 480220 3068
rect 480548 480 480576 4966
rect 481560 4146 481588 41806
rect 482296 39030 482324 41806
rect 483308 39438 483336 41806
rect 483020 39432 483072 39438
rect 483020 39374 483072 39380
rect 483296 39432 483348 39438
rect 483296 39374 483348 39380
rect 482284 39024 482336 39030
rect 482284 38966 482336 38972
rect 482928 39024 482980 39030
rect 482928 38966 482980 38972
rect 481548 4140 481600 4146
rect 481548 4082 481600 4088
rect 481732 3800 481784 3806
rect 481732 3742 481784 3748
rect 481744 480 481772 3742
rect 482940 3398 482968 38966
rect 483032 16574 483060 39374
rect 484412 39030 484440 41806
rect 484400 39024 484452 39030
rect 484400 38966 484452 38972
rect 485596 39024 485648 39030
rect 485596 38966 485648 38972
rect 483032 16546 484072 16574
rect 482836 3392 482888 3398
rect 482836 3334 482888 3340
rect 482928 3392 482980 3398
rect 482928 3334 482980 3340
rect 482848 480 482876 3334
rect 484044 480 484072 16546
rect 485608 4078 485636 38966
rect 485596 4072 485648 4078
rect 485596 4014 485648 4020
rect 485700 3806 485728 41806
rect 486436 39030 486464 41806
rect 487448 39030 487476 41806
rect 488460 39710 488488 41806
rect 488448 39704 488500 39710
rect 488448 39646 488500 39652
rect 486424 39024 486476 39030
rect 486424 38966 486476 38972
rect 487068 39024 487120 39030
rect 487068 38966 487120 38972
rect 487436 39024 487488 39030
rect 487436 38966 487488 38972
rect 488448 39024 488500 39030
rect 488448 38966 488500 38972
rect 487080 5098 487108 38966
rect 487068 5092 487120 5098
rect 487068 5034 487120 5040
rect 487620 4956 487672 4962
rect 487620 4898 487672 4904
rect 485688 3800 485740 3806
rect 485688 3742 485740 3748
rect 486424 3324 486476 3330
rect 486424 3266 486476 3272
rect 485228 2984 485280 2990
rect 485228 2926 485280 2932
rect 485240 480 485268 2926
rect 486436 480 486464 3266
rect 487632 480 487660 4898
rect 488460 3330 488488 38966
rect 489840 5030 489868 41806
rect 490012 39636 490064 39642
rect 490012 39578 490064 39584
rect 490024 16574 490052 39578
rect 490484 38826 490512 41806
rect 491496 39642 491524 41806
rect 491484 39636 491536 39642
rect 491484 39578 491536 39584
rect 492508 39030 492536 41806
rect 492496 39024 492548 39030
rect 492496 38966 492548 38972
rect 493324 39024 493376 39030
rect 493324 38966 493376 38972
rect 490472 38820 490524 38826
rect 490472 38762 490524 38768
rect 491208 38820 491260 38826
rect 491208 38762 491260 38768
rect 490024 16546 490696 16574
rect 489828 5024 489880 5030
rect 489828 4966 489880 4972
rect 488816 4004 488868 4010
rect 488816 3946 488868 3952
rect 488448 3324 488500 3330
rect 488448 3266 488500 3272
rect 488828 480 488856 3946
rect 489920 3936 489972 3942
rect 489920 3878 489972 3884
rect 489932 480 489960 3878
rect 490668 490 490696 16546
rect 491220 4010 491248 38762
rect 493336 4962 493364 38966
rect 493520 38758 493548 41806
rect 494532 39030 494560 41806
rect 495544 39982 495572 41806
rect 495532 39976 495584 39982
rect 495532 39918 495584 39924
rect 494520 39024 494572 39030
rect 494520 38966 494572 38972
rect 495348 39024 495400 39030
rect 495348 38966 495400 38972
rect 493508 38752 493560 38758
rect 493508 38694 493560 38700
rect 493968 38752 494020 38758
rect 493968 38694 494020 38700
rect 493324 4956 493376 4962
rect 493324 4898 493376 4904
rect 491208 4004 491260 4010
rect 491208 3946 491260 3952
rect 493980 3942 494008 38694
rect 494704 4888 494756 4894
rect 494704 4830 494756 4836
rect 493968 3936 494020 3942
rect 493968 3878 494020 3884
rect 493508 3868 493560 3874
rect 493508 3810 493560 3816
rect 492312 3052 492364 3058
rect 492312 2994 492364 3000
rect 490944 598 491156 626
rect 490944 490 490972 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 462 490972 490
rect 491128 480 491156 598
rect 492324 480 492352 2994
rect 493520 480 493548 3810
rect 494716 480 494744 4830
rect 495360 3874 495388 38966
rect 495348 3868 495400 3874
rect 495348 3810 495400 3816
rect 496740 3670 496768 41806
rect 497464 39704 497516 39710
rect 497464 39646 497516 39652
rect 495900 3664 495952 3670
rect 495900 3606 495952 3612
rect 496728 3664 496780 3670
rect 496728 3606 496780 3612
rect 495912 480 495940 3606
rect 497096 3528 497148 3534
rect 497096 3470 497148 3476
rect 497108 480 497136 3470
rect 497476 2922 497504 39646
rect 497568 39030 497596 41806
rect 498580 39778 498608 41806
rect 498568 39772 498620 39778
rect 498568 39714 498620 39720
rect 497556 39024 497608 39030
rect 497556 38966 497608 38972
rect 498108 39024 498160 39030
rect 498108 38966 498160 38972
rect 498120 3534 498148 38966
rect 499684 38962 499712 41806
rect 499672 38956 499724 38962
rect 499672 38898 499724 38904
rect 500776 38956 500828 38962
rect 500776 38898 500828 38904
rect 498200 4820 498252 4826
rect 498200 4762 498252 4768
rect 498108 3528 498160 3534
rect 498108 3470 498160 3476
rect 497464 2916 497516 2922
rect 497464 2858 497516 2864
rect 498212 480 498240 4762
rect 499396 3732 499448 3738
rect 499396 3674 499448 3680
rect 499408 480 499436 3674
rect 500788 3602 500816 38898
rect 500880 3738 500908 41806
rect 501708 39846 501736 41806
rect 501696 39840 501748 39846
rect 501696 39782 501748 39788
rect 500960 39296 501012 39302
rect 500960 39238 501012 39244
rect 500972 16574 501000 39238
rect 502720 39030 502748 41806
rect 503732 39574 503760 41806
rect 502984 39568 503036 39574
rect 502984 39510 503036 39516
rect 503720 39568 503772 39574
rect 503720 39510 503772 39516
rect 502708 39024 502760 39030
rect 502708 38966 502760 38972
rect 500972 16546 501368 16574
rect 500868 3732 500920 3738
rect 500868 3674 500920 3680
rect 500592 3596 500644 3602
rect 500592 3538 500644 3544
rect 500776 3596 500828 3602
rect 500776 3538 500828 3544
rect 500604 480 500632 3538
rect 501340 490 501368 16546
rect 502996 4214 503024 39510
rect 503628 39024 503680 39030
rect 503628 38966 503680 38972
rect 502984 4208 503036 4214
rect 502984 4150 503036 4156
rect 502984 3188 503036 3194
rect 502984 3130 503036 3136
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 3130
rect 503640 2990 503668 38966
rect 505020 4894 505048 41806
rect 505756 39030 505784 41806
rect 506768 39030 506796 41806
rect 507688 41806 507762 41834
rect 508746 41834 508774 42092
rect 509758 41834 509786 42092
rect 510770 41834 510798 42092
rect 511782 41834 511810 42092
rect 512794 41834 512822 42092
rect 513806 41834 513834 42092
rect 514910 41834 514938 42092
rect 515922 41834 515950 42092
rect 516934 41834 516962 42092
rect 517946 41834 517974 42092
rect 518958 41834 518986 42092
rect 519970 41834 519998 42092
rect 520982 41834 521010 42092
rect 521994 41834 522022 42092
rect 523006 41834 523034 42092
rect 524018 41834 524046 42092
rect 525030 41834 525058 42092
rect 526042 41834 526070 42092
rect 527054 41834 527082 42092
rect 528066 41834 528094 42092
rect 529078 41834 529106 42092
rect 530182 41834 530210 42092
rect 531194 41834 531222 42092
rect 508746 41806 509188 41834
rect 509758 41806 509832 41834
rect 510770 41806 510844 41834
rect 511782 41806 511948 41834
rect 512794 41806 512868 41834
rect 513806 41806 513880 41834
rect 514910 41806 514984 41834
rect 515922 41806 515996 41834
rect 516934 41806 517008 41834
rect 517946 41806 518020 41834
rect 518958 41806 519032 41834
rect 519970 41806 520044 41834
rect 520982 41806 521056 41834
rect 521994 41806 522068 41834
rect 523006 41806 523080 41834
rect 524018 41806 524368 41834
rect 525030 41806 525104 41834
rect 526042 41806 526116 41834
rect 527054 41806 527128 41834
rect 528066 41806 528140 41834
rect 529078 41806 529152 41834
rect 530182 41806 530256 41834
rect 505744 39024 505796 39030
rect 505744 38966 505796 38972
rect 506388 39024 506440 39030
rect 506388 38966 506440 38972
rect 506756 39024 506808 39030
rect 506756 38966 506808 38972
rect 505008 4888 505060 4894
rect 505008 4830 505060 4836
rect 505376 4208 505428 4214
rect 505376 4150 505428 4156
rect 504180 3460 504232 3466
rect 504180 3402 504232 3408
rect 503628 2984 503680 2990
rect 503628 2926 503680 2932
rect 504192 480 504220 3402
rect 505388 480 505416 4150
rect 506400 3466 506428 38966
rect 507688 4826 507716 41806
rect 507860 39500 507912 39506
rect 507860 39442 507912 39448
rect 507768 39024 507820 39030
rect 507768 38966 507820 38972
rect 507676 4820 507728 4826
rect 507676 4762 507728 4768
rect 506388 3460 506440 3466
rect 506388 3402 506440 3408
rect 506480 3256 506532 3262
rect 506480 3198 506532 3204
rect 506492 480 506520 3198
rect 507780 3194 507808 38966
rect 507872 16574 507900 39442
rect 507872 16546 508912 16574
rect 507768 3188 507820 3194
rect 507768 3130 507820 3136
rect 507676 3120 507728 3126
rect 507676 3062 507728 3068
rect 507688 480 507716 3062
rect 508884 480 508912 16546
rect 509160 3058 509188 41806
rect 509804 40050 509832 41806
rect 509792 40044 509844 40050
rect 509792 39986 509844 39992
rect 510816 39370 510844 41806
rect 510804 39364 510856 39370
rect 510804 39306 510856 39312
rect 510068 4140 510120 4146
rect 510068 4082 510120 4088
rect 509148 3052 509200 3058
rect 509148 2994 509200 3000
rect 510080 480 510108 4082
rect 511920 3398 511948 41806
rect 512840 39710 512868 41806
rect 513852 39982 513880 41806
rect 513840 39976 513892 39982
rect 513840 39918 513892 39924
rect 512828 39704 512880 39710
rect 512828 39646 512880 39652
rect 512644 39636 512696 39642
rect 512644 39578 512696 39584
rect 512000 39432 512052 39438
rect 512000 39374 512052 39380
rect 511264 3392 511316 3398
rect 511264 3334 511316 3340
rect 511908 3392 511960 3398
rect 511908 3334 511960 3340
rect 511276 480 511304 3334
rect 512012 490 512040 39374
rect 512656 3262 512684 39578
rect 514956 39030 514984 41806
rect 515404 39908 515456 39914
rect 515404 39850 515456 39856
rect 514944 39024 514996 39030
rect 514944 38966 514996 38972
rect 515416 5166 515444 39850
rect 515968 39642 515996 41806
rect 515956 39636 516008 39642
rect 515956 39578 516008 39584
rect 516980 39506 517008 41806
rect 516968 39500 517020 39506
rect 516968 39442 517020 39448
rect 517992 39030 518020 41806
rect 518164 39772 518216 39778
rect 518164 39714 518216 39720
rect 516048 39024 516100 39030
rect 516048 38966 516100 38972
rect 517980 39024 518032 39030
rect 517980 38966 518032 38972
rect 515404 5160 515456 5166
rect 515404 5102 515456 5108
rect 515956 5092 516008 5098
rect 515956 5034 516008 5040
rect 513564 4072 513616 4078
rect 513564 4014 513616 4020
rect 512644 3256 512696 3262
rect 512644 3198 512696 3204
rect 512288 598 512500 626
rect 512288 490 512316 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 462 512316 490
rect 512472 480 512500 598
rect 513576 480 513604 4014
rect 514760 3800 514812 3806
rect 514760 3742 514812 3748
rect 514772 480 514800 3742
rect 515968 480 515996 5034
rect 516060 3126 516088 38966
rect 518176 5098 518204 39714
rect 519004 39030 519032 41806
rect 520016 39438 520044 41806
rect 520004 39432 520056 39438
rect 520004 39374 520056 39380
rect 518808 39024 518860 39030
rect 518808 38966 518860 38972
rect 518992 39024 519044 39030
rect 518992 38966 519044 38972
rect 520188 39024 520240 39030
rect 520188 38966 520240 38972
rect 518164 5092 518216 5098
rect 518164 5034 518216 5040
rect 518820 4146 518848 38966
rect 519544 5024 519596 5030
rect 519544 4966 519596 4972
rect 518808 4140 518860 4146
rect 518808 4082 518860 4088
rect 517152 3324 517204 3330
rect 517152 3266 517204 3272
rect 516048 3120 516100 3126
rect 516048 3062 516100 3068
rect 517164 480 517192 3266
rect 518348 2916 518400 2922
rect 518348 2858 518400 2864
rect 518360 480 518388 2858
rect 519556 480 519584 4966
rect 520200 3330 520228 38966
rect 521028 38826 521056 41806
rect 522040 39030 522068 41806
rect 523052 39574 523080 41806
rect 522304 39568 522356 39574
rect 522304 39510 522356 39516
rect 523040 39568 523092 39574
rect 523040 39510 523092 39516
rect 522028 39024 522080 39030
rect 522028 38966 522080 38972
rect 521016 38820 521068 38826
rect 521016 38762 521068 38768
rect 521568 38820 521620 38826
rect 521568 38762 521620 38768
rect 521580 4010 521608 38762
rect 520740 4004 520792 4010
rect 520740 3946 520792 3952
rect 521568 4004 521620 4010
rect 521568 3946 521620 3952
rect 520188 3324 520240 3330
rect 520188 3266 520240 3272
rect 520752 480 520780 3946
rect 521844 3256 521896 3262
rect 521844 3198 521896 3204
rect 521856 480 521884 3198
rect 522316 2922 522344 39510
rect 522948 39024 523000 39030
rect 522948 38966 523000 38972
rect 522960 3262 522988 38966
rect 523040 4956 523092 4962
rect 523040 4898 523092 4904
rect 522948 3256 523000 3262
rect 522948 3198 523000 3204
rect 522304 2916 522356 2922
rect 522304 2858 522356 2864
rect 523052 480 523080 4898
rect 524340 3942 524368 41806
rect 524972 39976 525024 39982
rect 524972 39918 525024 39924
rect 524984 35894 525012 39918
rect 525076 39030 525104 41806
rect 526088 39778 526116 41806
rect 526076 39772 526128 39778
rect 526076 39714 526128 39720
rect 525064 39024 525116 39030
rect 525064 38966 525116 38972
rect 525708 39024 525760 39030
rect 525708 38966 525760 38972
rect 524984 35866 525104 35894
rect 525076 4962 525104 35866
rect 525064 4956 525116 4962
rect 525064 4898 525116 4904
rect 525720 4078 525748 38966
rect 526628 5160 526680 5166
rect 526628 5102 526680 5108
rect 525708 4072 525760 4078
rect 525708 4014 525760 4020
rect 524236 3936 524288 3942
rect 524236 3878 524288 3884
rect 524328 3936 524380 3942
rect 524328 3878 524380 3884
rect 524248 480 524276 3878
rect 525432 3868 525484 3874
rect 525432 3810 525484 3816
rect 525444 480 525472 3810
rect 526640 480 526668 5102
rect 527100 3806 527128 41806
rect 528112 39302 528140 41806
rect 528100 39296 528152 39302
rect 528100 39238 528152 39244
rect 529124 39030 529152 41806
rect 530228 39030 530256 41806
rect 531148 41806 531222 41834
rect 532206 41834 532234 42092
rect 533218 41834 533246 42092
rect 534230 41834 534258 42092
rect 535242 41834 535270 42092
rect 536254 41834 536282 42092
rect 537266 41834 537294 42092
rect 538278 41834 538306 42092
rect 539290 41834 539318 42092
rect 540302 41834 540330 42092
rect 541314 41834 541342 42092
rect 542326 41834 542354 42092
rect 543352 42078 543688 42106
rect 532206 41806 532280 41834
rect 533218 41806 533292 41834
rect 534230 41806 534304 41834
rect 535242 41806 535316 41834
rect 536254 41806 536328 41834
rect 537266 41806 537340 41834
rect 538278 41806 538352 41834
rect 539290 41806 539548 41834
rect 540302 41806 540376 41834
rect 541314 41806 541388 41834
rect 542326 41806 542400 41834
rect 529112 39024 529164 39030
rect 529112 38966 529164 38972
rect 529848 39024 529900 39030
rect 529848 38966 529900 38972
rect 530216 39024 530268 39030
rect 530216 38966 530268 38972
rect 529860 6186 529888 38966
rect 529848 6180 529900 6186
rect 529848 6122 529900 6128
rect 530124 5092 530176 5098
rect 530124 5034 530176 5040
rect 527088 3800 527140 3806
rect 527088 3742 527140 3748
rect 527824 3664 527876 3670
rect 527824 3606 527876 3612
rect 527836 480 527864 3606
rect 529020 3528 529072 3534
rect 529020 3470 529072 3476
rect 529032 480 529060 3470
rect 530136 480 530164 5034
rect 531148 3534 531176 41806
rect 532252 39982 532280 41806
rect 532240 39976 532292 39982
rect 532240 39918 532292 39924
rect 532700 39840 532752 39846
rect 532700 39782 532752 39788
rect 531228 39024 531280 39030
rect 531228 38966 531280 38972
rect 531240 3874 531268 38966
rect 532712 16574 532740 39782
rect 533264 39030 533292 41806
rect 534276 39234 534304 41806
rect 535288 39846 535316 41806
rect 535276 39840 535328 39846
rect 535276 39782 535328 39788
rect 534264 39228 534316 39234
rect 534264 39170 534316 39176
rect 533252 39024 533304 39030
rect 533252 38966 533304 38972
rect 533988 39024 534040 39030
rect 533988 38966 534040 38972
rect 532712 16546 533752 16574
rect 531228 3868 531280 3874
rect 531228 3810 531280 3816
rect 532516 3732 532568 3738
rect 532516 3674 532568 3680
rect 531320 3596 531372 3602
rect 531320 3538 531372 3544
rect 531136 3528 531188 3534
rect 531136 3470 531188 3476
rect 531332 480 531360 3538
rect 532528 480 532556 3674
rect 533724 480 533752 16546
rect 534000 3738 534028 38966
rect 536300 38894 536328 41806
rect 537312 39030 537340 41806
rect 538324 40050 538352 41806
rect 538312 40044 538364 40050
rect 538312 39986 538364 39992
rect 537300 39024 537352 39030
rect 537300 38966 537352 38972
rect 538128 39024 538180 39030
rect 538128 38966 538180 38972
rect 536288 38888 536340 38894
rect 536288 38830 536340 38836
rect 536748 38888 536800 38894
rect 536748 38830 536800 38836
rect 533988 3732 534040 3738
rect 533988 3674 534040 3680
rect 536760 3670 536788 38830
rect 537208 4888 537260 4894
rect 537208 4830 537260 4836
rect 536748 3664 536800 3670
rect 536748 3606 536800 3612
rect 534908 2984 534960 2990
rect 534908 2926 534960 2932
rect 534920 480 534948 2926
rect 536104 2916 536156 2922
rect 536104 2858 536156 2864
rect 536116 480 536144 2858
rect 537220 480 537248 4830
rect 538140 3602 538168 38966
rect 538128 3596 538180 3602
rect 538128 3538 538180 3544
rect 538404 3460 538456 3466
rect 538404 3402 538456 3408
rect 538416 480 538444 3402
rect 539520 2990 539548 41806
rect 540244 39296 540296 39302
rect 540244 39238 540296 39244
rect 539600 3188 539652 3194
rect 539600 3130 539652 3136
rect 539508 2984 539560 2990
rect 539508 2926 539560 2932
rect 539612 480 539640 3130
rect 540256 2922 540284 39238
rect 540348 39030 540376 41806
rect 540428 39908 540480 39914
rect 540428 39850 540480 39856
rect 540336 39024 540388 39030
rect 540336 38966 540388 38972
rect 540440 26234 540468 39850
rect 541360 39710 541388 41806
rect 542372 39914 542400 41806
rect 542360 39908 542412 39914
rect 542360 39850 542412 39856
rect 541348 39704 541400 39710
rect 541348 39646 541400 39652
rect 543660 39370 543688 42078
rect 544384 39636 544436 39642
rect 544384 39578 544436 39584
rect 543004 39364 543056 39370
rect 543004 39306 543056 39312
rect 543648 39364 543700 39370
rect 543648 39306 543700 39312
rect 541624 39228 541676 39234
rect 541624 39170 541676 39176
rect 540348 26206 540468 26234
rect 540348 3466 540376 26206
rect 540796 4820 540848 4826
rect 540796 4762 540848 4768
rect 540336 3460 540388 3466
rect 540336 3402 540388 3408
rect 540244 2916 540296 2922
rect 540244 2858 540296 2864
rect 540808 480 540836 4762
rect 541636 2854 541664 39170
rect 543016 4214 543044 39306
rect 544396 16574 544424 39578
rect 545764 39024 545816 39030
rect 545764 38966 545816 38972
rect 544396 16546 544516 16574
rect 543004 4208 543056 4214
rect 543004 4150 543056 4156
rect 544384 4208 544436 4214
rect 544384 4150 544436 4156
rect 543188 3460 543240 3466
rect 543188 3402 543240 3408
rect 541992 3052 542044 3058
rect 541992 2994 542044 3000
rect 541624 2848 541676 2854
rect 541624 2790 541676 2796
rect 542004 480 542032 2994
rect 543200 480 543228 3402
rect 544396 480 544424 4150
rect 544488 3466 544516 16546
rect 544476 3460 544528 3466
rect 544476 3402 544528 3408
rect 545488 3392 545540 3398
rect 545488 3334 545540 3340
rect 545500 480 545528 3334
rect 545776 2990 545804 38966
rect 547156 6866 547184 545255
rect 547248 313274 547276 545974
rect 547236 313268 547288 313274
rect 547236 313210 547288 313216
rect 548536 86970 548564 546722
rect 548628 511970 548656 547742
rect 551376 547120 551428 547126
rect 551376 547062 551428 547068
rect 551282 546816 551338 546825
rect 551282 546751 551338 546760
rect 548616 511964 548668 511970
rect 548616 511906 548668 511912
rect 548524 86964 548576 86970
rect 548524 86906 548576 86912
rect 548616 39908 548668 39914
rect 548616 39850 548668 39856
rect 548524 39704 548576 39710
rect 548524 39646 548576 39652
rect 547236 39296 547288 39302
rect 547236 39238 547288 39244
rect 547144 6860 547196 6866
rect 547144 6802 547196 6808
rect 546684 3460 546736 3466
rect 546684 3402 546736 3408
rect 545764 2984 545816 2990
rect 545764 2926 545816 2932
rect 546696 480 546724 3402
rect 547248 3398 547276 39238
rect 547880 4956 547932 4962
rect 547880 4898 547932 4904
rect 547236 3392 547288 3398
rect 547236 3334 547288 3340
rect 547892 480 547920 4898
rect 548536 3194 548564 39646
rect 548524 3188 548576 3194
rect 548524 3130 548576 3136
rect 548628 3058 548656 39850
rect 550640 39500 550692 39506
rect 550640 39442 550692 39448
rect 550652 16574 550680 39442
rect 551296 20670 551324 546751
rect 551388 167006 551416 547062
rect 554056 525774 554084 549102
rect 565176 549024 565228 549030
rect 565176 548966 565228 548972
rect 561036 548752 561088 548758
rect 561036 548694 561088 548700
rect 558184 548004 558236 548010
rect 558184 547946 558236 547952
rect 556896 547256 556948 547262
rect 556896 547198 556948 547204
rect 555516 547188 555568 547194
rect 555516 547130 555568 547136
rect 555422 546680 555478 546689
rect 555422 546615 555478 546624
rect 554044 525768 554096 525774
rect 554044 525710 554096 525716
rect 551376 167000 551428 167006
rect 551376 166942 551428 166948
rect 554780 39432 554832 39438
rect 554780 39374 554832 39380
rect 551284 20664 551336 20670
rect 551284 20606 551336 20612
rect 554792 16574 554820 39374
rect 555436 33114 555464 546615
rect 555528 206990 555556 547130
rect 556804 546576 556856 546582
rect 556804 546518 556856 546524
rect 555516 206984 555568 206990
rect 555516 206926 555568 206932
rect 556816 73166 556844 546518
rect 556908 245614 556936 547198
rect 556896 245608 556948 245614
rect 556896 245550 556948 245556
rect 558196 113150 558224 547946
rect 558276 547324 558328 547330
rect 558276 547266 558328 547272
rect 558288 299470 558316 547266
rect 560944 546848 560996 546854
rect 560944 546790 560996 546796
rect 558276 299464 558328 299470
rect 558276 299406 558328 299412
rect 560956 153202 560984 546790
rect 561048 353258 561076 548694
rect 562324 548276 562376 548282
rect 562324 548218 562376 548224
rect 561036 353252 561088 353258
rect 561036 353194 561088 353200
rect 562336 193186 562364 548218
rect 562416 546100 562468 546106
rect 562416 546042 562468 546048
rect 562428 405686 562456 546042
rect 565084 545556 565136 545562
rect 565084 545498 565136 545504
rect 562416 405680 562468 405686
rect 562416 405622 562468 405628
rect 565096 233238 565124 545498
rect 565188 485790 565216 548966
rect 576216 548956 576268 548962
rect 576216 548898 576268 548904
rect 574836 548820 574888 548826
rect 574836 548762 574888 548768
rect 573456 548684 573508 548690
rect 573456 548626 573508 548632
rect 569316 545692 569368 545698
rect 569316 545634 569368 545640
rect 566556 545624 566608 545630
rect 566556 545566 566608 545572
rect 566464 545148 566516 545154
rect 566464 545090 566516 545096
rect 565176 485784 565228 485790
rect 565176 485726 565228 485732
rect 565084 233232 565136 233238
rect 565084 233174 565136 233180
rect 562324 193180 562376 193186
rect 562324 193122 562376 193128
rect 560944 153196 560996 153202
rect 560944 153138 560996 153144
rect 558184 113144 558236 113150
rect 558184 113086 558236 113092
rect 556804 73160 556856 73166
rect 556804 73102 556856 73108
rect 566476 60722 566504 545090
rect 566568 273222 566596 545566
rect 569224 545216 569276 545222
rect 569224 545158 569276 545164
rect 566556 273216 566608 273222
rect 566556 273158 566608 273164
rect 569236 100706 569264 545158
rect 569328 325650 569356 545634
rect 573364 545352 573416 545358
rect 573364 545294 573416 545300
rect 569316 325644 569368 325650
rect 569316 325586 569368 325592
rect 573376 139398 573404 545294
rect 573468 379506 573496 548626
rect 574744 545420 574796 545426
rect 574744 545362 574796 545368
rect 573456 379500 573508 379506
rect 573456 379442 573508 379448
rect 574756 179382 574784 545362
rect 574848 431934 574876 548762
rect 576124 545488 576176 545494
rect 576124 545430 576176 545436
rect 574836 431928 574888 431934
rect 574836 431870 574888 431876
rect 576136 219434 576164 545430
rect 576228 471986 576256 548898
rect 580448 547596 580500 547602
rect 580448 547538 580500 547544
rect 580264 546440 580316 546446
rect 580264 546382 580316 546388
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580172 525768 580224 525774
rect 580172 525710 580224 525716
rect 580184 524521 580212 525710
rect 580170 524512 580226 524521
rect 580170 524447 580226 524456
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 576216 471980 576268 471986
rect 576216 471922 576268 471928
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 580276 258913 580304 546382
rect 580356 545760 580408 545766
rect 580356 545702 580408 545708
rect 580368 365129 580396 545702
rect 580460 418305 580488 547538
rect 580446 418296 580502 418305
rect 580446 418231 580502 418240
rect 580354 365120 580410 365129
rect 580354 365055 580410 365064
rect 580262 258904 580318 258913
rect 580262 258839 580318 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 576124 219428 576176 219434
rect 576124 219370 576176 219376
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 574744 179376 574796 179382
rect 574744 179318 574796 179324
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 573364 139392 573416 139398
rect 580172 139392 580224 139398
rect 573364 139334 573416 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 569224 100700 569276 100706
rect 569224 100642 569276 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 566464 60716 566516 60722
rect 566464 60658 566516 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 565084 40044 565136 40050
rect 565084 39986 565136 39992
rect 560944 39976 560996 39982
rect 560944 39918 560996 39924
rect 558184 39772 558236 39778
rect 558184 39714 558236 39720
rect 556804 39568 556856 39574
rect 556804 39510 556856 39516
rect 555424 33108 555476 33114
rect 555424 33050 555476 33056
rect 550652 16546 551048 16574
rect 554792 16546 555004 16574
rect 550272 3392 550324 3398
rect 550272 3334 550324 3340
rect 549076 3120 549128 3126
rect 549076 3062 549128 3068
rect 548616 3052 548668 3058
rect 548616 2994 548668 3000
rect 549088 480 549116 3062
rect 550284 480 550312 3334
rect 551020 490 551048 16546
rect 552664 4140 552716 4146
rect 552664 4082 552716 4088
rect 551296 598 551508 626
rect 551296 490 551324 598
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 462 551324 490
rect 551480 480 551508 598
rect 552676 480 552704 4082
rect 553768 3324 553820 3330
rect 553768 3266 553820 3272
rect 553780 480 553808 3266
rect 554976 480 555004 16546
rect 556816 5642 556844 39510
rect 556804 5636 556856 5642
rect 556804 5578 556856 5584
rect 558196 5574 558224 39714
rect 560956 5642 560984 39918
rect 562324 39840 562376 39846
rect 562324 39782 562376 39788
rect 562336 6254 562364 39782
rect 562324 6248 562376 6254
rect 562324 6190 562376 6196
rect 565096 6186 565124 39986
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 572720 6248 572772 6254
rect 572720 6190 572772 6196
rect 565084 6180 565136 6186
rect 565084 6122 565136 6128
rect 565636 6112 565688 6118
rect 565636 6054 565688 6060
rect 558552 5636 558604 5642
rect 558552 5578 558604 5584
rect 560944 5636 560996 5642
rect 560944 5578 560996 5584
rect 558184 5568 558236 5574
rect 558184 5510 558236 5516
rect 556160 4004 556212 4010
rect 556160 3946 556212 3952
rect 556172 480 556200 3946
rect 557356 3188 557408 3194
rect 557356 3130 557408 3136
rect 557368 480 557396 3130
rect 558564 480 558592 5578
rect 562048 5568 562100 5574
rect 562048 5510 562100 5516
rect 560852 4072 560904 4078
rect 560852 4014 560904 4020
rect 559748 3936 559800 3942
rect 559748 3878 559800 3884
rect 559760 480 559788 3878
rect 560864 480 560892 4014
rect 562060 480 562088 5510
rect 563244 3800 563296 3806
rect 563244 3742 563296 3748
rect 563256 480 563284 3742
rect 564440 2916 564492 2922
rect 564440 2858 564492 2864
rect 564452 480 564480 2858
rect 565648 480 565676 6054
rect 569132 5636 569184 5642
rect 569132 5578 569184 5584
rect 566832 3868 566884 3874
rect 566832 3810 566884 3816
rect 566844 480 566872 3810
rect 568028 3528 568080 3534
rect 568028 3470 568080 3476
rect 568040 480 568068 3470
rect 569144 480 569172 5578
rect 570328 3732 570380 3738
rect 570328 3674 570380 3680
rect 570340 480 570368 3674
rect 571524 2984 571576 2990
rect 571524 2926 571576 2932
rect 571536 480 571564 2926
rect 572732 480 572760 6190
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 573916 3664 573968 3670
rect 573916 3606 573968 3612
rect 573928 480 573956 3606
rect 575112 3596 575164 3602
rect 575112 3538 575164 3544
rect 575124 480 575152 3538
rect 576320 480 576348 6122
rect 577412 3460 577464 3466
rect 577412 3402 577464 3408
rect 577424 480 577452 3402
rect 578608 3392 578660 3398
rect 578608 3334 578660 3340
rect 578620 480 578648 3334
rect 581000 3188 581052 3194
rect 581000 3130 581052 3136
rect 581012 480 581040 3130
rect 582196 3052 582248 3058
rect 582196 2994 582248 3000
rect 583392 3052 583444 3058
rect 583392 2994 583444 3000
rect 582208 480 582236 2994
rect 583404 480 583432 2994
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 7562 547984 7618 548040
rect 3514 547848 3570 547904
rect 3422 545672 3478 545728
rect 3330 527856 3386 527912
rect 3146 514800 3202 514856
rect 2962 501744 3018 501800
rect 3238 475632 3294 475688
rect 3054 462576 3110 462632
rect 3330 449520 3386 449576
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 2962 410488 3018 410544
rect 3330 397432 3386 397488
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 2778 267144 2834 267200
rect 3146 254088 3202 254144
rect 3238 241032 3294 241088
rect 3330 214956 3332 214976
rect 3332 214956 3384 214976
rect 3384 214956 3386 214976
rect 3330 214920 3386 214956
rect 3054 201864 3110 201920
rect 3146 188808 3202 188864
rect 3330 162832 3386 162888
rect 3330 136720 3386 136776
rect 3146 110608 3202 110664
rect 3238 97552 3294 97608
rect 3330 84632 3386 84688
rect 2778 71612 2780 71632
rect 2780 71612 2832 71632
rect 2832 71612 2834 71632
rect 2778 71576 2834 71612
rect 3606 149776 3662 149832
rect 3514 58520 3570 58576
rect 14462 546488 14518 546544
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 15842 545128 15898 545184
rect 18602 548120 18658 548176
rect 53194 546760 53250 546816
rect 48778 546624 48834 546680
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 510618 548120 510674 548176
rect 523682 547984 523738 548040
rect 528098 547848 528154 547904
rect 532698 546488 532754 546544
rect 471518 545672 471574 545728
rect 44454 545400 44510 545456
rect 536930 545400 536986 545456
rect 547142 545264 547198 545320
rect 551282 546760 551338 546816
rect 555422 546624 555478 546680
rect 580170 537784 580226 537840
rect 580170 524456 580226 524512
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 431568 580226 431624
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 351872 580226 351928
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 579618 298696 579674 298752
rect 579894 272176 579950 272232
rect 580446 418240 580502 418296
rect 580354 365064 580410 365120
rect 580262 258848 580318 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect 18597 548178 18663 548181
rect 510613 548178 510679 548181
rect 18597 548176 510679 548178
rect 18597 548120 18602 548176
rect 18658 548120 510618 548176
rect 510674 548120 510679 548176
rect 18597 548118 510679 548120
rect 18597 548115 18663 548118
rect 510613 548115 510679 548118
rect 7557 548042 7623 548045
rect 523677 548042 523743 548045
rect 7557 548040 523743 548042
rect 7557 547984 7562 548040
rect 7618 547984 523682 548040
rect 523738 547984 523743 548040
rect 7557 547982 523743 547984
rect 7557 547979 7623 547982
rect 523677 547979 523743 547982
rect 3509 547906 3575 547909
rect 528093 547906 528159 547909
rect 3509 547904 528159 547906
rect 3509 547848 3514 547904
rect 3570 547848 528098 547904
rect 528154 547848 528159 547904
rect 3509 547846 528159 547848
rect 3509 547843 3575 547846
rect 528093 547843 528159 547846
rect 53189 546818 53255 546821
rect 551277 546818 551343 546821
rect 53189 546816 551343 546818
rect 53189 546760 53194 546816
rect 53250 546760 551282 546816
rect 551338 546760 551343 546816
rect 53189 546758 551343 546760
rect 53189 546755 53255 546758
rect 551277 546755 551343 546758
rect 48773 546682 48839 546685
rect 555417 546682 555483 546685
rect 48773 546680 555483 546682
rect 48773 546624 48778 546680
rect 48834 546624 555422 546680
rect 555478 546624 555483 546680
rect 48773 546622 555483 546624
rect 48773 546619 48839 546622
rect 555417 546619 555483 546622
rect 14457 546546 14523 546549
rect 532693 546546 532759 546549
rect 14457 546544 532759 546546
rect 14457 546488 14462 546544
rect 14518 546488 532698 546544
rect 532754 546488 532759 546544
rect 14457 546486 532759 546488
rect 14457 546483 14523 546486
rect 532693 546483 532759 546486
rect 3417 545730 3483 545733
rect 471513 545730 471579 545733
rect 3417 545728 471579 545730
rect 3417 545672 3422 545728
rect 3478 545672 471518 545728
rect 471574 545672 471579 545728
rect 3417 545670 471579 545672
rect 3417 545667 3483 545670
rect 471513 545667 471579 545670
rect 528510 545534 538230 545594
rect 44449 545458 44515 545461
rect 44449 545456 45570 545458
rect 44449 545400 44454 545456
rect 44510 545400 45570 545456
rect 44449 545398 45570 545400
rect 44449 545395 44515 545398
rect 45510 545322 45570 545398
rect 528510 545322 528570 545534
rect 536925 545458 536991 545461
rect 45510 545262 528570 545322
rect 532742 545456 536991 545458
rect 532742 545400 536930 545456
rect 536986 545400 536991 545456
rect 532742 545398 536991 545400
rect 15837 545186 15903 545189
rect 532742 545186 532802 545398
rect 536925 545395 536991 545398
rect 538170 545322 538230 545534
rect 547137 545322 547203 545325
rect 538170 545320 547203 545322
rect 538170 545264 547142 545320
rect 547198 545264 547203 545320
rect 538170 545262 547203 545264
rect 547137 545259 547203 545262
rect 15837 545184 532802 545186
rect 15837 545128 15842 545184
rect 15898 545128 532802 545184
rect 15837 545126 532802 545128
rect 15837 545123 15903 545126
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3141 514858 3207 514861
rect -960 514856 3207 514858
rect -960 514800 3146 514856
rect 3202 514800 3207 514856
rect -960 514798 3207 514800
rect -960 514708 480 514798
rect 3141 514795 3207 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2957 501802 3023 501805
rect -960 501800 3023 501802
rect -960 501744 2962 501800
rect 3018 501744 3023 501800
rect -960 501742 3023 501744
rect -960 501652 480 501742
rect 2957 501739 3023 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3233 475690 3299 475693
rect -960 475688 3299 475690
rect -960 475632 3238 475688
rect 3294 475632 3299 475688
rect -960 475630 3299 475632
rect -960 475540 480 475630
rect 3233 475627 3299 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3049 462634 3115 462637
rect -960 462632 3115 462634
rect -960 462576 3054 462632
rect 3110 462576 3115 462632
rect -960 462574 3115 462576
rect -960 462484 480 462574
rect 3049 462571 3115 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580441 418298 580507 418301
rect 583520 418298 584960 418388
rect 580441 418296 584960 418298
rect 580441 418240 580446 418296
rect 580502 418240 584960 418296
rect 580441 418238 584960 418240
rect 580441 418235 580507 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580349 365122 580415 365125
rect 583520 365122 584960 365212
rect 580349 365120 584960 365122
rect 580349 365064 580354 365120
rect 580410 365064 584960 365120
rect 580349 365062 584960 365064
rect 580349 365059 580415 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2773 267202 2839 267205
rect -960 267200 2839 267202
rect -960 267144 2778 267200
rect 2834 267144 2839 267200
rect -960 267142 2839 267144
rect -960 267052 480 267142
rect 2773 267139 2839 267142
rect 580257 258906 580323 258909
rect 583520 258906 584960 258996
rect 580257 258904 584960 258906
rect 580257 258848 580262 258904
rect 580318 258848 584960 258904
rect 580257 258846 584960 258848
rect 580257 258843 580323 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 2773 71634 2839 71637
rect -960 71632 2839 71634
rect -960 71576 2778 71632
rect 2834 71576 2839 71632
rect -960 71574 2839 71576
rect -960 71484 480 71574
rect 2773 71571 2839 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 548086 42134 582618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 548086 45854 550338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 548086 49574 554058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 548086 56414 560898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 548086 60134 564618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 548086 63854 568338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 548086 67574 572058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 548086 74414 578898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 548086 78134 582618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 548086 81854 550338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 548086 85574 554058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 548086 92414 560898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 548086 96134 564618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 548086 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 548086 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 548086 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 548086 114134 582618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 548086 117854 550338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 548086 121574 554058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 548086 128414 560898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 548086 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 548086 135854 568338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 548086 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 548086 146414 578898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 548086 150134 582618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 548086 153854 550338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 548086 157574 554058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 548086 164414 560898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 548086 168134 564618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 548086 171854 568338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 548086 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 548086 182414 578898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 548086 186134 582618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 548086 189854 550338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 548086 193574 554058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 548086 200414 560898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 548086 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 548086 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 548086 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 548086 218414 578898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 548086 222134 582618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 548086 225854 550338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 548086 229574 554058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 548086 236414 560898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 548086 240134 564618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 548086 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 548086 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 548086 254414 578898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 548086 258134 582618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 548086 261854 550338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 548086 265574 554058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 548086 272414 560898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 548086 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 548086 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 548086 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 548086 290414 578898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 548086 294134 582618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 548086 297854 550338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 548086 301574 554058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 548086 308414 560898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 548086 312134 564618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 548086 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 548086 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 548086 326414 578898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 548086 330134 582618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 548086 333854 550338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 548086 337574 554058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 548086 344414 560898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 548086 348134 564618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 548086 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 548086 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 548086 362414 578898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 548086 366134 582618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 548086 369854 550338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 548086 373574 554058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 548086 380414 560898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 548086 384134 564618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 548086 387854 568338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 548086 391574 572058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 548086 398414 578898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 548086 402134 582618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 548086 405854 550338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 548086 409574 554058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 548086 416414 560898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 548086 420134 564618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 548086 423854 568338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 548086 427574 572058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 548086 434414 578898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 548086 438134 582618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 548086 441854 550338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 548086 445574 554058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 548086 452414 560898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 548086 456134 564618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 548086 459854 568338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 548086 463574 572058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 548086 470414 578898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 548086 474134 582618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 548086 477854 550338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 548086 481574 554058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 548086 488414 560898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 548086 492134 564618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 548086 495854 568338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 548086 499574 572058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 548086 506414 578898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 548086 510134 582618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 548086 513854 550338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 548086 517574 554058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 548086 524414 560898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 548086 528134 564618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 548086 531854 568338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 548086 535574 572058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 548086 542414 578898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 548086 546134 582618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 46208 543454 46528 543486
rect 46208 543218 46250 543454
rect 46486 543218 46528 543454
rect 46208 543134 46528 543218
rect 46208 542898 46250 543134
rect 46486 542898 46528 543134
rect 46208 542866 46528 542898
rect 76928 543454 77248 543486
rect 76928 543218 76970 543454
rect 77206 543218 77248 543454
rect 76928 543134 77248 543218
rect 76928 542898 76970 543134
rect 77206 542898 77248 543134
rect 76928 542866 77248 542898
rect 107648 543454 107968 543486
rect 107648 543218 107690 543454
rect 107926 543218 107968 543454
rect 107648 543134 107968 543218
rect 107648 542898 107690 543134
rect 107926 542898 107968 543134
rect 107648 542866 107968 542898
rect 138368 543454 138688 543486
rect 138368 543218 138410 543454
rect 138646 543218 138688 543454
rect 138368 543134 138688 543218
rect 138368 542898 138410 543134
rect 138646 542898 138688 543134
rect 138368 542866 138688 542898
rect 169088 543454 169408 543486
rect 169088 543218 169130 543454
rect 169366 543218 169408 543454
rect 169088 543134 169408 543218
rect 169088 542898 169130 543134
rect 169366 542898 169408 543134
rect 169088 542866 169408 542898
rect 199808 543454 200128 543486
rect 199808 543218 199850 543454
rect 200086 543218 200128 543454
rect 199808 543134 200128 543218
rect 199808 542898 199850 543134
rect 200086 542898 200128 543134
rect 199808 542866 200128 542898
rect 230528 543454 230848 543486
rect 230528 543218 230570 543454
rect 230806 543218 230848 543454
rect 230528 543134 230848 543218
rect 230528 542898 230570 543134
rect 230806 542898 230848 543134
rect 230528 542866 230848 542898
rect 261248 543454 261568 543486
rect 261248 543218 261290 543454
rect 261526 543218 261568 543454
rect 261248 543134 261568 543218
rect 261248 542898 261290 543134
rect 261526 542898 261568 543134
rect 261248 542866 261568 542898
rect 291968 543454 292288 543486
rect 291968 543218 292010 543454
rect 292246 543218 292288 543454
rect 291968 543134 292288 543218
rect 291968 542898 292010 543134
rect 292246 542898 292288 543134
rect 291968 542866 292288 542898
rect 322688 543454 323008 543486
rect 322688 543218 322730 543454
rect 322966 543218 323008 543454
rect 322688 543134 323008 543218
rect 322688 542898 322730 543134
rect 322966 542898 323008 543134
rect 322688 542866 323008 542898
rect 353408 543454 353728 543486
rect 353408 543218 353450 543454
rect 353686 543218 353728 543454
rect 353408 543134 353728 543218
rect 353408 542898 353450 543134
rect 353686 542898 353728 543134
rect 353408 542866 353728 542898
rect 384128 543454 384448 543486
rect 384128 543218 384170 543454
rect 384406 543218 384448 543454
rect 384128 543134 384448 543218
rect 384128 542898 384170 543134
rect 384406 542898 384448 543134
rect 384128 542866 384448 542898
rect 414848 543454 415168 543486
rect 414848 543218 414890 543454
rect 415126 543218 415168 543454
rect 414848 543134 415168 543218
rect 414848 542898 414890 543134
rect 415126 542898 415168 543134
rect 414848 542866 415168 542898
rect 445568 543454 445888 543486
rect 445568 543218 445610 543454
rect 445846 543218 445888 543454
rect 445568 543134 445888 543218
rect 445568 542898 445610 543134
rect 445846 542898 445888 543134
rect 445568 542866 445888 542898
rect 476288 543454 476608 543486
rect 476288 543218 476330 543454
rect 476566 543218 476608 543454
rect 476288 543134 476608 543218
rect 476288 542898 476330 543134
rect 476566 542898 476608 543134
rect 476288 542866 476608 542898
rect 507008 543454 507328 543486
rect 507008 543218 507050 543454
rect 507286 543218 507328 543454
rect 507008 543134 507328 543218
rect 507008 542898 507050 543134
rect 507286 542898 507328 543134
rect 507008 542866 507328 542898
rect 537728 543454 538048 543486
rect 537728 543218 537770 543454
rect 538006 543218 538048 543454
rect 537728 543134 538048 543218
rect 537728 542898 537770 543134
rect 538006 542898 538048 543134
rect 537728 542866 538048 542898
rect 61568 525454 61888 525486
rect 61568 525218 61610 525454
rect 61846 525218 61888 525454
rect 61568 525134 61888 525218
rect 61568 524898 61610 525134
rect 61846 524898 61888 525134
rect 61568 524866 61888 524898
rect 92288 525454 92608 525486
rect 92288 525218 92330 525454
rect 92566 525218 92608 525454
rect 92288 525134 92608 525218
rect 92288 524898 92330 525134
rect 92566 524898 92608 525134
rect 92288 524866 92608 524898
rect 123008 525454 123328 525486
rect 123008 525218 123050 525454
rect 123286 525218 123328 525454
rect 123008 525134 123328 525218
rect 123008 524898 123050 525134
rect 123286 524898 123328 525134
rect 123008 524866 123328 524898
rect 153728 525454 154048 525486
rect 153728 525218 153770 525454
rect 154006 525218 154048 525454
rect 153728 525134 154048 525218
rect 153728 524898 153770 525134
rect 154006 524898 154048 525134
rect 153728 524866 154048 524898
rect 184448 525454 184768 525486
rect 184448 525218 184490 525454
rect 184726 525218 184768 525454
rect 184448 525134 184768 525218
rect 184448 524898 184490 525134
rect 184726 524898 184768 525134
rect 184448 524866 184768 524898
rect 215168 525454 215488 525486
rect 215168 525218 215210 525454
rect 215446 525218 215488 525454
rect 215168 525134 215488 525218
rect 215168 524898 215210 525134
rect 215446 524898 215488 525134
rect 215168 524866 215488 524898
rect 245888 525454 246208 525486
rect 245888 525218 245930 525454
rect 246166 525218 246208 525454
rect 245888 525134 246208 525218
rect 245888 524898 245930 525134
rect 246166 524898 246208 525134
rect 245888 524866 246208 524898
rect 276608 525454 276928 525486
rect 276608 525218 276650 525454
rect 276886 525218 276928 525454
rect 276608 525134 276928 525218
rect 276608 524898 276650 525134
rect 276886 524898 276928 525134
rect 276608 524866 276928 524898
rect 307328 525454 307648 525486
rect 307328 525218 307370 525454
rect 307606 525218 307648 525454
rect 307328 525134 307648 525218
rect 307328 524898 307370 525134
rect 307606 524898 307648 525134
rect 307328 524866 307648 524898
rect 338048 525454 338368 525486
rect 338048 525218 338090 525454
rect 338326 525218 338368 525454
rect 338048 525134 338368 525218
rect 338048 524898 338090 525134
rect 338326 524898 338368 525134
rect 338048 524866 338368 524898
rect 368768 525454 369088 525486
rect 368768 525218 368810 525454
rect 369046 525218 369088 525454
rect 368768 525134 369088 525218
rect 368768 524898 368810 525134
rect 369046 524898 369088 525134
rect 368768 524866 369088 524898
rect 399488 525454 399808 525486
rect 399488 525218 399530 525454
rect 399766 525218 399808 525454
rect 399488 525134 399808 525218
rect 399488 524898 399530 525134
rect 399766 524898 399808 525134
rect 399488 524866 399808 524898
rect 430208 525454 430528 525486
rect 430208 525218 430250 525454
rect 430486 525218 430528 525454
rect 430208 525134 430528 525218
rect 430208 524898 430250 525134
rect 430486 524898 430528 525134
rect 430208 524866 430528 524898
rect 460928 525454 461248 525486
rect 460928 525218 460970 525454
rect 461206 525218 461248 525454
rect 460928 525134 461248 525218
rect 460928 524898 460970 525134
rect 461206 524898 461248 525134
rect 460928 524866 461248 524898
rect 491648 525454 491968 525486
rect 491648 525218 491690 525454
rect 491926 525218 491968 525454
rect 491648 525134 491968 525218
rect 491648 524898 491690 525134
rect 491926 524898 491968 525134
rect 491648 524866 491968 524898
rect 522368 525454 522688 525486
rect 522368 525218 522410 525454
rect 522646 525218 522688 525454
rect 522368 525134 522688 525218
rect 522368 524898 522410 525134
rect 522646 524898 522688 525134
rect 522368 524866 522688 524898
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 46208 507454 46528 507486
rect 46208 507218 46250 507454
rect 46486 507218 46528 507454
rect 46208 507134 46528 507218
rect 46208 506898 46250 507134
rect 46486 506898 46528 507134
rect 46208 506866 46528 506898
rect 76928 507454 77248 507486
rect 76928 507218 76970 507454
rect 77206 507218 77248 507454
rect 76928 507134 77248 507218
rect 76928 506898 76970 507134
rect 77206 506898 77248 507134
rect 76928 506866 77248 506898
rect 107648 507454 107968 507486
rect 107648 507218 107690 507454
rect 107926 507218 107968 507454
rect 107648 507134 107968 507218
rect 107648 506898 107690 507134
rect 107926 506898 107968 507134
rect 107648 506866 107968 506898
rect 138368 507454 138688 507486
rect 138368 507218 138410 507454
rect 138646 507218 138688 507454
rect 138368 507134 138688 507218
rect 138368 506898 138410 507134
rect 138646 506898 138688 507134
rect 138368 506866 138688 506898
rect 169088 507454 169408 507486
rect 169088 507218 169130 507454
rect 169366 507218 169408 507454
rect 169088 507134 169408 507218
rect 169088 506898 169130 507134
rect 169366 506898 169408 507134
rect 169088 506866 169408 506898
rect 199808 507454 200128 507486
rect 199808 507218 199850 507454
rect 200086 507218 200128 507454
rect 199808 507134 200128 507218
rect 199808 506898 199850 507134
rect 200086 506898 200128 507134
rect 199808 506866 200128 506898
rect 230528 507454 230848 507486
rect 230528 507218 230570 507454
rect 230806 507218 230848 507454
rect 230528 507134 230848 507218
rect 230528 506898 230570 507134
rect 230806 506898 230848 507134
rect 230528 506866 230848 506898
rect 261248 507454 261568 507486
rect 261248 507218 261290 507454
rect 261526 507218 261568 507454
rect 261248 507134 261568 507218
rect 261248 506898 261290 507134
rect 261526 506898 261568 507134
rect 261248 506866 261568 506898
rect 291968 507454 292288 507486
rect 291968 507218 292010 507454
rect 292246 507218 292288 507454
rect 291968 507134 292288 507218
rect 291968 506898 292010 507134
rect 292246 506898 292288 507134
rect 291968 506866 292288 506898
rect 322688 507454 323008 507486
rect 322688 507218 322730 507454
rect 322966 507218 323008 507454
rect 322688 507134 323008 507218
rect 322688 506898 322730 507134
rect 322966 506898 323008 507134
rect 322688 506866 323008 506898
rect 353408 507454 353728 507486
rect 353408 507218 353450 507454
rect 353686 507218 353728 507454
rect 353408 507134 353728 507218
rect 353408 506898 353450 507134
rect 353686 506898 353728 507134
rect 353408 506866 353728 506898
rect 384128 507454 384448 507486
rect 384128 507218 384170 507454
rect 384406 507218 384448 507454
rect 384128 507134 384448 507218
rect 384128 506898 384170 507134
rect 384406 506898 384448 507134
rect 384128 506866 384448 506898
rect 414848 507454 415168 507486
rect 414848 507218 414890 507454
rect 415126 507218 415168 507454
rect 414848 507134 415168 507218
rect 414848 506898 414890 507134
rect 415126 506898 415168 507134
rect 414848 506866 415168 506898
rect 445568 507454 445888 507486
rect 445568 507218 445610 507454
rect 445846 507218 445888 507454
rect 445568 507134 445888 507218
rect 445568 506898 445610 507134
rect 445846 506898 445888 507134
rect 445568 506866 445888 506898
rect 476288 507454 476608 507486
rect 476288 507218 476330 507454
rect 476566 507218 476608 507454
rect 476288 507134 476608 507218
rect 476288 506898 476330 507134
rect 476566 506898 476608 507134
rect 476288 506866 476608 506898
rect 507008 507454 507328 507486
rect 507008 507218 507050 507454
rect 507286 507218 507328 507454
rect 507008 507134 507328 507218
rect 507008 506898 507050 507134
rect 507286 506898 507328 507134
rect 507008 506866 507328 506898
rect 537728 507454 538048 507486
rect 537728 507218 537770 507454
rect 538006 507218 538048 507454
rect 537728 507134 538048 507218
rect 537728 506898 537770 507134
rect 538006 506898 538048 507134
rect 537728 506866 538048 506898
rect 61568 489454 61888 489486
rect 61568 489218 61610 489454
rect 61846 489218 61888 489454
rect 61568 489134 61888 489218
rect 61568 488898 61610 489134
rect 61846 488898 61888 489134
rect 61568 488866 61888 488898
rect 92288 489454 92608 489486
rect 92288 489218 92330 489454
rect 92566 489218 92608 489454
rect 92288 489134 92608 489218
rect 92288 488898 92330 489134
rect 92566 488898 92608 489134
rect 92288 488866 92608 488898
rect 123008 489454 123328 489486
rect 123008 489218 123050 489454
rect 123286 489218 123328 489454
rect 123008 489134 123328 489218
rect 123008 488898 123050 489134
rect 123286 488898 123328 489134
rect 123008 488866 123328 488898
rect 153728 489454 154048 489486
rect 153728 489218 153770 489454
rect 154006 489218 154048 489454
rect 153728 489134 154048 489218
rect 153728 488898 153770 489134
rect 154006 488898 154048 489134
rect 153728 488866 154048 488898
rect 184448 489454 184768 489486
rect 184448 489218 184490 489454
rect 184726 489218 184768 489454
rect 184448 489134 184768 489218
rect 184448 488898 184490 489134
rect 184726 488898 184768 489134
rect 184448 488866 184768 488898
rect 215168 489454 215488 489486
rect 215168 489218 215210 489454
rect 215446 489218 215488 489454
rect 215168 489134 215488 489218
rect 215168 488898 215210 489134
rect 215446 488898 215488 489134
rect 215168 488866 215488 488898
rect 245888 489454 246208 489486
rect 245888 489218 245930 489454
rect 246166 489218 246208 489454
rect 245888 489134 246208 489218
rect 245888 488898 245930 489134
rect 246166 488898 246208 489134
rect 245888 488866 246208 488898
rect 276608 489454 276928 489486
rect 276608 489218 276650 489454
rect 276886 489218 276928 489454
rect 276608 489134 276928 489218
rect 276608 488898 276650 489134
rect 276886 488898 276928 489134
rect 276608 488866 276928 488898
rect 307328 489454 307648 489486
rect 307328 489218 307370 489454
rect 307606 489218 307648 489454
rect 307328 489134 307648 489218
rect 307328 488898 307370 489134
rect 307606 488898 307648 489134
rect 307328 488866 307648 488898
rect 338048 489454 338368 489486
rect 338048 489218 338090 489454
rect 338326 489218 338368 489454
rect 338048 489134 338368 489218
rect 338048 488898 338090 489134
rect 338326 488898 338368 489134
rect 338048 488866 338368 488898
rect 368768 489454 369088 489486
rect 368768 489218 368810 489454
rect 369046 489218 369088 489454
rect 368768 489134 369088 489218
rect 368768 488898 368810 489134
rect 369046 488898 369088 489134
rect 368768 488866 369088 488898
rect 399488 489454 399808 489486
rect 399488 489218 399530 489454
rect 399766 489218 399808 489454
rect 399488 489134 399808 489218
rect 399488 488898 399530 489134
rect 399766 488898 399808 489134
rect 399488 488866 399808 488898
rect 430208 489454 430528 489486
rect 430208 489218 430250 489454
rect 430486 489218 430528 489454
rect 430208 489134 430528 489218
rect 430208 488898 430250 489134
rect 430486 488898 430528 489134
rect 430208 488866 430528 488898
rect 460928 489454 461248 489486
rect 460928 489218 460970 489454
rect 461206 489218 461248 489454
rect 460928 489134 461248 489218
rect 460928 488898 460970 489134
rect 461206 488898 461248 489134
rect 460928 488866 461248 488898
rect 491648 489454 491968 489486
rect 491648 489218 491690 489454
rect 491926 489218 491968 489454
rect 491648 489134 491968 489218
rect 491648 488898 491690 489134
rect 491926 488898 491968 489134
rect 491648 488866 491968 488898
rect 522368 489454 522688 489486
rect 522368 489218 522410 489454
rect 522646 489218 522688 489454
rect 522368 489134 522688 489218
rect 522368 488898 522410 489134
rect 522646 488898 522688 489134
rect 522368 488866 522688 488898
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 46208 471454 46528 471486
rect 46208 471218 46250 471454
rect 46486 471218 46528 471454
rect 46208 471134 46528 471218
rect 46208 470898 46250 471134
rect 46486 470898 46528 471134
rect 46208 470866 46528 470898
rect 76928 471454 77248 471486
rect 76928 471218 76970 471454
rect 77206 471218 77248 471454
rect 76928 471134 77248 471218
rect 76928 470898 76970 471134
rect 77206 470898 77248 471134
rect 76928 470866 77248 470898
rect 107648 471454 107968 471486
rect 107648 471218 107690 471454
rect 107926 471218 107968 471454
rect 107648 471134 107968 471218
rect 107648 470898 107690 471134
rect 107926 470898 107968 471134
rect 107648 470866 107968 470898
rect 138368 471454 138688 471486
rect 138368 471218 138410 471454
rect 138646 471218 138688 471454
rect 138368 471134 138688 471218
rect 138368 470898 138410 471134
rect 138646 470898 138688 471134
rect 138368 470866 138688 470898
rect 169088 471454 169408 471486
rect 169088 471218 169130 471454
rect 169366 471218 169408 471454
rect 169088 471134 169408 471218
rect 169088 470898 169130 471134
rect 169366 470898 169408 471134
rect 169088 470866 169408 470898
rect 199808 471454 200128 471486
rect 199808 471218 199850 471454
rect 200086 471218 200128 471454
rect 199808 471134 200128 471218
rect 199808 470898 199850 471134
rect 200086 470898 200128 471134
rect 199808 470866 200128 470898
rect 230528 471454 230848 471486
rect 230528 471218 230570 471454
rect 230806 471218 230848 471454
rect 230528 471134 230848 471218
rect 230528 470898 230570 471134
rect 230806 470898 230848 471134
rect 230528 470866 230848 470898
rect 261248 471454 261568 471486
rect 261248 471218 261290 471454
rect 261526 471218 261568 471454
rect 261248 471134 261568 471218
rect 261248 470898 261290 471134
rect 261526 470898 261568 471134
rect 261248 470866 261568 470898
rect 291968 471454 292288 471486
rect 291968 471218 292010 471454
rect 292246 471218 292288 471454
rect 291968 471134 292288 471218
rect 291968 470898 292010 471134
rect 292246 470898 292288 471134
rect 291968 470866 292288 470898
rect 322688 471454 323008 471486
rect 322688 471218 322730 471454
rect 322966 471218 323008 471454
rect 322688 471134 323008 471218
rect 322688 470898 322730 471134
rect 322966 470898 323008 471134
rect 322688 470866 323008 470898
rect 353408 471454 353728 471486
rect 353408 471218 353450 471454
rect 353686 471218 353728 471454
rect 353408 471134 353728 471218
rect 353408 470898 353450 471134
rect 353686 470898 353728 471134
rect 353408 470866 353728 470898
rect 384128 471454 384448 471486
rect 384128 471218 384170 471454
rect 384406 471218 384448 471454
rect 384128 471134 384448 471218
rect 384128 470898 384170 471134
rect 384406 470898 384448 471134
rect 384128 470866 384448 470898
rect 414848 471454 415168 471486
rect 414848 471218 414890 471454
rect 415126 471218 415168 471454
rect 414848 471134 415168 471218
rect 414848 470898 414890 471134
rect 415126 470898 415168 471134
rect 414848 470866 415168 470898
rect 445568 471454 445888 471486
rect 445568 471218 445610 471454
rect 445846 471218 445888 471454
rect 445568 471134 445888 471218
rect 445568 470898 445610 471134
rect 445846 470898 445888 471134
rect 445568 470866 445888 470898
rect 476288 471454 476608 471486
rect 476288 471218 476330 471454
rect 476566 471218 476608 471454
rect 476288 471134 476608 471218
rect 476288 470898 476330 471134
rect 476566 470898 476608 471134
rect 476288 470866 476608 470898
rect 507008 471454 507328 471486
rect 507008 471218 507050 471454
rect 507286 471218 507328 471454
rect 507008 471134 507328 471218
rect 507008 470898 507050 471134
rect 507286 470898 507328 471134
rect 507008 470866 507328 470898
rect 537728 471454 538048 471486
rect 537728 471218 537770 471454
rect 538006 471218 538048 471454
rect 537728 471134 538048 471218
rect 537728 470898 537770 471134
rect 538006 470898 538048 471134
rect 537728 470866 538048 470898
rect 61568 453454 61888 453486
rect 61568 453218 61610 453454
rect 61846 453218 61888 453454
rect 61568 453134 61888 453218
rect 61568 452898 61610 453134
rect 61846 452898 61888 453134
rect 61568 452866 61888 452898
rect 92288 453454 92608 453486
rect 92288 453218 92330 453454
rect 92566 453218 92608 453454
rect 92288 453134 92608 453218
rect 92288 452898 92330 453134
rect 92566 452898 92608 453134
rect 92288 452866 92608 452898
rect 123008 453454 123328 453486
rect 123008 453218 123050 453454
rect 123286 453218 123328 453454
rect 123008 453134 123328 453218
rect 123008 452898 123050 453134
rect 123286 452898 123328 453134
rect 123008 452866 123328 452898
rect 153728 453454 154048 453486
rect 153728 453218 153770 453454
rect 154006 453218 154048 453454
rect 153728 453134 154048 453218
rect 153728 452898 153770 453134
rect 154006 452898 154048 453134
rect 153728 452866 154048 452898
rect 184448 453454 184768 453486
rect 184448 453218 184490 453454
rect 184726 453218 184768 453454
rect 184448 453134 184768 453218
rect 184448 452898 184490 453134
rect 184726 452898 184768 453134
rect 184448 452866 184768 452898
rect 215168 453454 215488 453486
rect 215168 453218 215210 453454
rect 215446 453218 215488 453454
rect 215168 453134 215488 453218
rect 215168 452898 215210 453134
rect 215446 452898 215488 453134
rect 215168 452866 215488 452898
rect 245888 453454 246208 453486
rect 245888 453218 245930 453454
rect 246166 453218 246208 453454
rect 245888 453134 246208 453218
rect 245888 452898 245930 453134
rect 246166 452898 246208 453134
rect 245888 452866 246208 452898
rect 276608 453454 276928 453486
rect 276608 453218 276650 453454
rect 276886 453218 276928 453454
rect 276608 453134 276928 453218
rect 276608 452898 276650 453134
rect 276886 452898 276928 453134
rect 276608 452866 276928 452898
rect 307328 453454 307648 453486
rect 307328 453218 307370 453454
rect 307606 453218 307648 453454
rect 307328 453134 307648 453218
rect 307328 452898 307370 453134
rect 307606 452898 307648 453134
rect 307328 452866 307648 452898
rect 338048 453454 338368 453486
rect 338048 453218 338090 453454
rect 338326 453218 338368 453454
rect 338048 453134 338368 453218
rect 338048 452898 338090 453134
rect 338326 452898 338368 453134
rect 338048 452866 338368 452898
rect 368768 453454 369088 453486
rect 368768 453218 368810 453454
rect 369046 453218 369088 453454
rect 368768 453134 369088 453218
rect 368768 452898 368810 453134
rect 369046 452898 369088 453134
rect 368768 452866 369088 452898
rect 399488 453454 399808 453486
rect 399488 453218 399530 453454
rect 399766 453218 399808 453454
rect 399488 453134 399808 453218
rect 399488 452898 399530 453134
rect 399766 452898 399808 453134
rect 399488 452866 399808 452898
rect 430208 453454 430528 453486
rect 430208 453218 430250 453454
rect 430486 453218 430528 453454
rect 430208 453134 430528 453218
rect 430208 452898 430250 453134
rect 430486 452898 430528 453134
rect 430208 452866 430528 452898
rect 460928 453454 461248 453486
rect 460928 453218 460970 453454
rect 461206 453218 461248 453454
rect 460928 453134 461248 453218
rect 460928 452898 460970 453134
rect 461206 452898 461248 453134
rect 460928 452866 461248 452898
rect 491648 453454 491968 453486
rect 491648 453218 491690 453454
rect 491926 453218 491968 453454
rect 491648 453134 491968 453218
rect 491648 452898 491690 453134
rect 491926 452898 491968 453134
rect 491648 452866 491968 452898
rect 522368 453454 522688 453486
rect 522368 453218 522410 453454
rect 522646 453218 522688 453454
rect 522368 453134 522688 453218
rect 522368 452898 522410 453134
rect 522646 452898 522688 453134
rect 522368 452866 522688 452898
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 46208 435454 46528 435486
rect 46208 435218 46250 435454
rect 46486 435218 46528 435454
rect 46208 435134 46528 435218
rect 46208 434898 46250 435134
rect 46486 434898 46528 435134
rect 46208 434866 46528 434898
rect 76928 435454 77248 435486
rect 76928 435218 76970 435454
rect 77206 435218 77248 435454
rect 76928 435134 77248 435218
rect 76928 434898 76970 435134
rect 77206 434898 77248 435134
rect 76928 434866 77248 434898
rect 107648 435454 107968 435486
rect 107648 435218 107690 435454
rect 107926 435218 107968 435454
rect 107648 435134 107968 435218
rect 107648 434898 107690 435134
rect 107926 434898 107968 435134
rect 107648 434866 107968 434898
rect 138368 435454 138688 435486
rect 138368 435218 138410 435454
rect 138646 435218 138688 435454
rect 138368 435134 138688 435218
rect 138368 434898 138410 435134
rect 138646 434898 138688 435134
rect 138368 434866 138688 434898
rect 169088 435454 169408 435486
rect 169088 435218 169130 435454
rect 169366 435218 169408 435454
rect 169088 435134 169408 435218
rect 169088 434898 169130 435134
rect 169366 434898 169408 435134
rect 169088 434866 169408 434898
rect 199808 435454 200128 435486
rect 199808 435218 199850 435454
rect 200086 435218 200128 435454
rect 199808 435134 200128 435218
rect 199808 434898 199850 435134
rect 200086 434898 200128 435134
rect 199808 434866 200128 434898
rect 230528 435454 230848 435486
rect 230528 435218 230570 435454
rect 230806 435218 230848 435454
rect 230528 435134 230848 435218
rect 230528 434898 230570 435134
rect 230806 434898 230848 435134
rect 230528 434866 230848 434898
rect 261248 435454 261568 435486
rect 261248 435218 261290 435454
rect 261526 435218 261568 435454
rect 261248 435134 261568 435218
rect 261248 434898 261290 435134
rect 261526 434898 261568 435134
rect 261248 434866 261568 434898
rect 291968 435454 292288 435486
rect 291968 435218 292010 435454
rect 292246 435218 292288 435454
rect 291968 435134 292288 435218
rect 291968 434898 292010 435134
rect 292246 434898 292288 435134
rect 291968 434866 292288 434898
rect 322688 435454 323008 435486
rect 322688 435218 322730 435454
rect 322966 435218 323008 435454
rect 322688 435134 323008 435218
rect 322688 434898 322730 435134
rect 322966 434898 323008 435134
rect 322688 434866 323008 434898
rect 353408 435454 353728 435486
rect 353408 435218 353450 435454
rect 353686 435218 353728 435454
rect 353408 435134 353728 435218
rect 353408 434898 353450 435134
rect 353686 434898 353728 435134
rect 353408 434866 353728 434898
rect 384128 435454 384448 435486
rect 384128 435218 384170 435454
rect 384406 435218 384448 435454
rect 384128 435134 384448 435218
rect 384128 434898 384170 435134
rect 384406 434898 384448 435134
rect 384128 434866 384448 434898
rect 414848 435454 415168 435486
rect 414848 435218 414890 435454
rect 415126 435218 415168 435454
rect 414848 435134 415168 435218
rect 414848 434898 414890 435134
rect 415126 434898 415168 435134
rect 414848 434866 415168 434898
rect 445568 435454 445888 435486
rect 445568 435218 445610 435454
rect 445846 435218 445888 435454
rect 445568 435134 445888 435218
rect 445568 434898 445610 435134
rect 445846 434898 445888 435134
rect 445568 434866 445888 434898
rect 476288 435454 476608 435486
rect 476288 435218 476330 435454
rect 476566 435218 476608 435454
rect 476288 435134 476608 435218
rect 476288 434898 476330 435134
rect 476566 434898 476608 435134
rect 476288 434866 476608 434898
rect 507008 435454 507328 435486
rect 507008 435218 507050 435454
rect 507286 435218 507328 435454
rect 507008 435134 507328 435218
rect 507008 434898 507050 435134
rect 507286 434898 507328 435134
rect 507008 434866 507328 434898
rect 537728 435454 538048 435486
rect 537728 435218 537770 435454
rect 538006 435218 538048 435454
rect 537728 435134 538048 435218
rect 537728 434898 537770 435134
rect 538006 434898 538048 435134
rect 537728 434866 538048 434898
rect 61568 417454 61888 417486
rect 61568 417218 61610 417454
rect 61846 417218 61888 417454
rect 61568 417134 61888 417218
rect 61568 416898 61610 417134
rect 61846 416898 61888 417134
rect 61568 416866 61888 416898
rect 92288 417454 92608 417486
rect 92288 417218 92330 417454
rect 92566 417218 92608 417454
rect 92288 417134 92608 417218
rect 92288 416898 92330 417134
rect 92566 416898 92608 417134
rect 92288 416866 92608 416898
rect 123008 417454 123328 417486
rect 123008 417218 123050 417454
rect 123286 417218 123328 417454
rect 123008 417134 123328 417218
rect 123008 416898 123050 417134
rect 123286 416898 123328 417134
rect 123008 416866 123328 416898
rect 153728 417454 154048 417486
rect 153728 417218 153770 417454
rect 154006 417218 154048 417454
rect 153728 417134 154048 417218
rect 153728 416898 153770 417134
rect 154006 416898 154048 417134
rect 153728 416866 154048 416898
rect 184448 417454 184768 417486
rect 184448 417218 184490 417454
rect 184726 417218 184768 417454
rect 184448 417134 184768 417218
rect 184448 416898 184490 417134
rect 184726 416898 184768 417134
rect 184448 416866 184768 416898
rect 215168 417454 215488 417486
rect 215168 417218 215210 417454
rect 215446 417218 215488 417454
rect 215168 417134 215488 417218
rect 215168 416898 215210 417134
rect 215446 416898 215488 417134
rect 215168 416866 215488 416898
rect 245888 417454 246208 417486
rect 245888 417218 245930 417454
rect 246166 417218 246208 417454
rect 245888 417134 246208 417218
rect 245888 416898 245930 417134
rect 246166 416898 246208 417134
rect 245888 416866 246208 416898
rect 276608 417454 276928 417486
rect 276608 417218 276650 417454
rect 276886 417218 276928 417454
rect 276608 417134 276928 417218
rect 276608 416898 276650 417134
rect 276886 416898 276928 417134
rect 276608 416866 276928 416898
rect 307328 417454 307648 417486
rect 307328 417218 307370 417454
rect 307606 417218 307648 417454
rect 307328 417134 307648 417218
rect 307328 416898 307370 417134
rect 307606 416898 307648 417134
rect 307328 416866 307648 416898
rect 338048 417454 338368 417486
rect 338048 417218 338090 417454
rect 338326 417218 338368 417454
rect 338048 417134 338368 417218
rect 338048 416898 338090 417134
rect 338326 416898 338368 417134
rect 338048 416866 338368 416898
rect 368768 417454 369088 417486
rect 368768 417218 368810 417454
rect 369046 417218 369088 417454
rect 368768 417134 369088 417218
rect 368768 416898 368810 417134
rect 369046 416898 369088 417134
rect 368768 416866 369088 416898
rect 399488 417454 399808 417486
rect 399488 417218 399530 417454
rect 399766 417218 399808 417454
rect 399488 417134 399808 417218
rect 399488 416898 399530 417134
rect 399766 416898 399808 417134
rect 399488 416866 399808 416898
rect 430208 417454 430528 417486
rect 430208 417218 430250 417454
rect 430486 417218 430528 417454
rect 430208 417134 430528 417218
rect 430208 416898 430250 417134
rect 430486 416898 430528 417134
rect 430208 416866 430528 416898
rect 460928 417454 461248 417486
rect 460928 417218 460970 417454
rect 461206 417218 461248 417454
rect 460928 417134 461248 417218
rect 460928 416898 460970 417134
rect 461206 416898 461248 417134
rect 460928 416866 461248 416898
rect 491648 417454 491968 417486
rect 491648 417218 491690 417454
rect 491926 417218 491968 417454
rect 491648 417134 491968 417218
rect 491648 416898 491690 417134
rect 491926 416898 491968 417134
rect 491648 416866 491968 416898
rect 522368 417454 522688 417486
rect 522368 417218 522410 417454
rect 522646 417218 522688 417454
rect 522368 417134 522688 417218
rect 522368 416898 522410 417134
rect 522646 416898 522688 417134
rect 522368 416866 522688 416898
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 46208 399454 46528 399486
rect 46208 399218 46250 399454
rect 46486 399218 46528 399454
rect 46208 399134 46528 399218
rect 46208 398898 46250 399134
rect 46486 398898 46528 399134
rect 46208 398866 46528 398898
rect 76928 399454 77248 399486
rect 76928 399218 76970 399454
rect 77206 399218 77248 399454
rect 76928 399134 77248 399218
rect 76928 398898 76970 399134
rect 77206 398898 77248 399134
rect 76928 398866 77248 398898
rect 107648 399454 107968 399486
rect 107648 399218 107690 399454
rect 107926 399218 107968 399454
rect 107648 399134 107968 399218
rect 107648 398898 107690 399134
rect 107926 398898 107968 399134
rect 107648 398866 107968 398898
rect 138368 399454 138688 399486
rect 138368 399218 138410 399454
rect 138646 399218 138688 399454
rect 138368 399134 138688 399218
rect 138368 398898 138410 399134
rect 138646 398898 138688 399134
rect 138368 398866 138688 398898
rect 169088 399454 169408 399486
rect 169088 399218 169130 399454
rect 169366 399218 169408 399454
rect 169088 399134 169408 399218
rect 169088 398898 169130 399134
rect 169366 398898 169408 399134
rect 169088 398866 169408 398898
rect 199808 399454 200128 399486
rect 199808 399218 199850 399454
rect 200086 399218 200128 399454
rect 199808 399134 200128 399218
rect 199808 398898 199850 399134
rect 200086 398898 200128 399134
rect 199808 398866 200128 398898
rect 230528 399454 230848 399486
rect 230528 399218 230570 399454
rect 230806 399218 230848 399454
rect 230528 399134 230848 399218
rect 230528 398898 230570 399134
rect 230806 398898 230848 399134
rect 230528 398866 230848 398898
rect 261248 399454 261568 399486
rect 261248 399218 261290 399454
rect 261526 399218 261568 399454
rect 261248 399134 261568 399218
rect 261248 398898 261290 399134
rect 261526 398898 261568 399134
rect 261248 398866 261568 398898
rect 291968 399454 292288 399486
rect 291968 399218 292010 399454
rect 292246 399218 292288 399454
rect 291968 399134 292288 399218
rect 291968 398898 292010 399134
rect 292246 398898 292288 399134
rect 291968 398866 292288 398898
rect 322688 399454 323008 399486
rect 322688 399218 322730 399454
rect 322966 399218 323008 399454
rect 322688 399134 323008 399218
rect 322688 398898 322730 399134
rect 322966 398898 323008 399134
rect 322688 398866 323008 398898
rect 353408 399454 353728 399486
rect 353408 399218 353450 399454
rect 353686 399218 353728 399454
rect 353408 399134 353728 399218
rect 353408 398898 353450 399134
rect 353686 398898 353728 399134
rect 353408 398866 353728 398898
rect 384128 399454 384448 399486
rect 384128 399218 384170 399454
rect 384406 399218 384448 399454
rect 384128 399134 384448 399218
rect 384128 398898 384170 399134
rect 384406 398898 384448 399134
rect 384128 398866 384448 398898
rect 414848 399454 415168 399486
rect 414848 399218 414890 399454
rect 415126 399218 415168 399454
rect 414848 399134 415168 399218
rect 414848 398898 414890 399134
rect 415126 398898 415168 399134
rect 414848 398866 415168 398898
rect 445568 399454 445888 399486
rect 445568 399218 445610 399454
rect 445846 399218 445888 399454
rect 445568 399134 445888 399218
rect 445568 398898 445610 399134
rect 445846 398898 445888 399134
rect 445568 398866 445888 398898
rect 476288 399454 476608 399486
rect 476288 399218 476330 399454
rect 476566 399218 476608 399454
rect 476288 399134 476608 399218
rect 476288 398898 476330 399134
rect 476566 398898 476608 399134
rect 476288 398866 476608 398898
rect 507008 399454 507328 399486
rect 507008 399218 507050 399454
rect 507286 399218 507328 399454
rect 507008 399134 507328 399218
rect 507008 398898 507050 399134
rect 507286 398898 507328 399134
rect 507008 398866 507328 398898
rect 537728 399454 538048 399486
rect 537728 399218 537770 399454
rect 538006 399218 538048 399454
rect 537728 399134 538048 399218
rect 537728 398898 537770 399134
rect 538006 398898 538048 399134
rect 537728 398866 538048 398898
rect 61568 381454 61888 381486
rect 61568 381218 61610 381454
rect 61846 381218 61888 381454
rect 61568 381134 61888 381218
rect 61568 380898 61610 381134
rect 61846 380898 61888 381134
rect 61568 380866 61888 380898
rect 92288 381454 92608 381486
rect 92288 381218 92330 381454
rect 92566 381218 92608 381454
rect 92288 381134 92608 381218
rect 92288 380898 92330 381134
rect 92566 380898 92608 381134
rect 92288 380866 92608 380898
rect 123008 381454 123328 381486
rect 123008 381218 123050 381454
rect 123286 381218 123328 381454
rect 123008 381134 123328 381218
rect 123008 380898 123050 381134
rect 123286 380898 123328 381134
rect 123008 380866 123328 380898
rect 153728 381454 154048 381486
rect 153728 381218 153770 381454
rect 154006 381218 154048 381454
rect 153728 381134 154048 381218
rect 153728 380898 153770 381134
rect 154006 380898 154048 381134
rect 153728 380866 154048 380898
rect 184448 381454 184768 381486
rect 184448 381218 184490 381454
rect 184726 381218 184768 381454
rect 184448 381134 184768 381218
rect 184448 380898 184490 381134
rect 184726 380898 184768 381134
rect 184448 380866 184768 380898
rect 215168 381454 215488 381486
rect 215168 381218 215210 381454
rect 215446 381218 215488 381454
rect 215168 381134 215488 381218
rect 215168 380898 215210 381134
rect 215446 380898 215488 381134
rect 215168 380866 215488 380898
rect 245888 381454 246208 381486
rect 245888 381218 245930 381454
rect 246166 381218 246208 381454
rect 245888 381134 246208 381218
rect 245888 380898 245930 381134
rect 246166 380898 246208 381134
rect 245888 380866 246208 380898
rect 276608 381454 276928 381486
rect 276608 381218 276650 381454
rect 276886 381218 276928 381454
rect 276608 381134 276928 381218
rect 276608 380898 276650 381134
rect 276886 380898 276928 381134
rect 276608 380866 276928 380898
rect 307328 381454 307648 381486
rect 307328 381218 307370 381454
rect 307606 381218 307648 381454
rect 307328 381134 307648 381218
rect 307328 380898 307370 381134
rect 307606 380898 307648 381134
rect 307328 380866 307648 380898
rect 338048 381454 338368 381486
rect 338048 381218 338090 381454
rect 338326 381218 338368 381454
rect 338048 381134 338368 381218
rect 338048 380898 338090 381134
rect 338326 380898 338368 381134
rect 338048 380866 338368 380898
rect 368768 381454 369088 381486
rect 368768 381218 368810 381454
rect 369046 381218 369088 381454
rect 368768 381134 369088 381218
rect 368768 380898 368810 381134
rect 369046 380898 369088 381134
rect 368768 380866 369088 380898
rect 399488 381454 399808 381486
rect 399488 381218 399530 381454
rect 399766 381218 399808 381454
rect 399488 381134 399808 381218
rect 399488 380898 399530 381134
rect 399766 380898 399808 381134
rect 399488 380866 399808 380898
rect 430208 381454 430528 381486
rect 430208 381218 430250 381454
rect 430486 381218 430528 381454
rect 430208 381134 430528 381218
rect 430208 380898 430250 381134
rect 430486 380898 430528 381134
rect 430208 380866 430528 380898
rect 460928 381454 461248 381486
rect 460928 381218 460970 381454
rect 461206 381218 461248 381454
rect 460928 381134 461248 381218
rect 460928 380898 460970 381134
rect 461206 380898 461248 381134
rect 460928 380866 461248 380898
rect 491648 381454 491968 381486
rect 491648 381218 491690 381454
rect 491926 381218 491968 381454
rect 491648 381134 491968 381218
rect 491648 380898 491690 381134
rect 491926 380898 491968 381134
rect 491648 380866 491968 380898
rect 522368 381454 522688 381486
rect 522368 381218 522410 381454
rect 522646 381218 522688 381454
rect 522368 381134 522688 381218
rect 522368 380898 522410 381134
rect 522646 380898 522688 381134
rect 522368 380866 522688 380898
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 46208 363454 46528 363486
rect 46208 363218 46250 363454
rect 46486 363218 46528 363454
rect 46208 363134 46528 363218
rect 46208 362898 46250 363134
rect 46486 362898 46528 363134
rect 46208 362866 46528 362898
rect 76928 363454 77248 363486
rect 76928 363218 76970 363454
rect 77206 363218 77248 363454
rect 76928 363134 77248 363218
rect 76928 362898 76970 363134
rect 77206 362898 77248 363134
rect 76928 362866 77248 362898
rect 107648 363454 107968 363486
rect 107648 363218 107690 363454
rect 107926 363218 107968 363454
rect 107648 363134 107968 363218
rect 107648 362898 107690 363134
rect 107926 362898 107968 363134
rect 107648 362866 107968 362898
rect 138368 363454 138688 363486
rect 138368 363218 138410 363454
rect 138646 363218 138688 363454
rect 138368 363134 138688 363218
rect 138368 362898 138410 363134
rect 138646 362898 138688 363134
rect 138368 362866 138688 362898
rect 169088 363454 169408 363486
rect 169088 363218 169130 363454
rect 169366 363218 169408 363454
rect 169088 363134 169408 363218
rect 169088 362898 169130 363134
rect 169366 362898 169408 363134
rect 169088 362866 169408 362898
rect 199808 363454 200128 363486
rect 199808 363218 199850 363454
rect 200086 363218 200128 363454
rect 199808 363134 200128 363218
rect 199808 362898 199850 363134
rect 200086 362898 200128 363134
rect 199808 362866 200128 362898
rect 230528 363454 230848 363486
rect 230528 363218 230570 363454
rect 230806 363218 230848 363454
rect 230528 363134 230848 363218
rect 230528 362898 230570 363134
rect 230806 362898 230848 363134
rect 230528 362866 230848 362898
rect 261248 363454 261568 363486
rect 261248 363218 261290 363454
rect 261526 363218 261568 363454
rect 261248 363134 261568 363218
rect 261248 362898 261290 363134
rect 261526 362898 261568 363134
rect 261248 362866 261568 362898
rect 291968 363454 292288 363486
rect 291968 363218 292010 363454
rect 292246 363218 292288 363454
rect 291968 363134 292288 363218
rect 291968 362898 292010 363134
rect 292246 362898 292288 363134
rect 291968 362866 292288 362898
rect 322688 363454 323008 363486
rect 322688 363218 322730 363454
rect 322966 363218 323008 363454
rect 322688 363134 323008 363218
rect 322688 362898 322730 363134
rect 322966 362898 323008 363134
rect 322688 362866 323008 362898
rect 353408 363454 353728 363486
rect 353408 363218 353450 363454
rect 353686 363218 353728 363454
rect 353408 363134 353728 363218
rect 353408 362898 353450 363134
rect 353686 362898 353728 363134
rect 353408 362866 353728 362898
rect 384128 363454 384448 363486
rect 384128 363218 384170 363454
rect 384406 363218 384448 363454
rect 384128 363134 384448 363218
rect 384128 362898 384170 363134
rect 384406 362898 384448 363134
rect 384128 362866 384448 362898
rect 414848 363454 415168 363486
rect 414848 363218 414890 363454
rect 415126 363218 415168 363454
rect 414848 363134 415168 363218
rect 414848 362898 414890 363134
rect 415126 362898 415168 363134
rect 414848 362866 415168 362898
rect 445568 363454 445888 363486
rect 445568 363218 445610 363454
rect 445846 363218 445888 363454
rect 445568 363134 445888 363218
rect 445568 362898 445610 363134
rect 445846 362898 445888 363134
rect 445568 362866 445888 362898
rect 476288 363454 476608 363486
rect 476288 363218 476330 363454
rect 476566 363218 476608 363454
rect 476288 363134 476608 363218
rect 476288 362898 476330 363134
rect 476566 362898 476608 363134
rect 476288 362866 476608 362898
rect 507008 363454 507328 363486
rect 507008 363218 507050 363454
rect 507286 363218 507328 363454
rect 507008 363134 507328 363218
rect 507008 362898 507050 363134
rect 507286 362898 507328 363134
rect 507008 362866 507328 362898
rect 537728 363454 538048 363486
rect 537728 363218 537770 363454
rect 538006 363218 538048 363454
rect 537728 363134 538048 363218
rect 537728 362898 537770 363134
rect 538006 362898 538048 363134
rect 537728 362866 538048 362898
rect 61568 345454 61888 345486
rect 61568 345218 61610 345454
rect 61846 345218 61888 345454
rect 61568 345134 61888 345218
rect 61568 344898 61610 345134
rect 61846 344898 61888 345134
rect 61568 344866 61888 344898
rect 92288 345454 92608 345486
rect 92288 345218 92330 345454
rect 92566 345218 92608 345454
rect 92288 345134 92608 345218
rect 92288 344898 92330 345134
rect 92566 344898 92608 345134
rect 92288 344866 92608 344898
rect 123008 345454 123328 345486
rect 123008 345218 123050 345454
rect 123286 345218 123328 345454
rect 123008 345134 123328 345218
rect 123008 344898 123050 345134
rect 123286 344898 123328 345134
rect 123008 344866 123328 344898
rect 153728 345454 154048 345486
rect 153728 345218 153770 345454
rect 154006 345218 154048 345454
rect 153728 345134 154048 345218
rect 153728 344898 153770 345134
rect 154006 344898 154048 345134
rect 153728 344866 154048 344898
rect 184448 345454 184768 345486
rect 184448 345218 184490 345454
rect 184726 345218 184768 345454
rect 184448 345134 184768 345218
rect 184448 344898 184490 345134
rect 184726 344898 184768 345134
rect 184448 344866 184768 344898
rect 215168 345454 215488 345486
rect 215168 345218 215210 345454
rect 215446 345218 215488 345454
rect 215168 345134 215488 345218
rect 215168 344898 215210 345134
rect 215446 344898 215488 345134
rect 215168 344866 215488 344898
rect 245888 345454 246208 345486
rect 245888 345218 245930 345454
rect 246166 345218 246208 345454
rect 245888 345134 246208 345218
rect 245888 344898 245930 345134
rect 246166 344898 246208 345134
rect 245888 344866 246208 344898
rect 276608 345454 276928 345486
rect 276608 345218 276650 345454
rect 276886 345218 276928 345454
rect 276608 345134 276928 345218
rect 276608 344898 276650 345134
rect 276886 344898 276928 345134
rect 276608 344866 276928 344898
rect 307328 345454 307648 345486
rect 307328 345218 307370 345454
rect 307606 345218 307648 345454
rect 307328 345134 307648 345218
rect 307328 344898 307370 345134
rect 307606 344898 307648 345134
rect 307328 344866 307648 344898
rect 338048 345454 338368 345486
rect 338048 345218 338090 345454
rect 338326 345218 338368 345454
rect 338048 345134 338368 345218
rect 338048 344898 338090 345134
rect 338326 344898 338368 345134
rect 338048 344866 338368 344898
rect 368768 345454 369088 345486
rect 368768 345218 368810 345454
rect 369046 345218 369088 345454
rect 368768 345134 369088 345218
rect 368768 344898 368810 345134
rect 369046 344898 369088 345134
rect 368768 344866 369088 344898
rect 399488 345454 399808 345486
rect 399488 345218 399530 345454
rect 399766 345218 399808 345454
rect 399488 345134 399808 345218
rect 399488 344898 399530 345134
rect 399766 344898 399808 345134
rect 399488 344866 399808 344898
rect 430208 345454 430528 345486
rect 430208 345218 430250 345454
rect 430486 345218 430528 345454
rect 430208 345134 430528 345218
rect 430208 344898 430250 345134
rect 430486 344898 430528 345134
rect 430208 344866 430528 344898
rect 460928 345454 461248 345486
rect 460928 345218 460970 345454
rect 461206 345218 461248 345454
rect 460928 345134 461248 345218
rect 460928 344898 460970 345134
rect 461206 344898 461248 345134
rect 460928 344866 461248 344898
rect 491648 345454 491968 345486
rect 491648 345218 491690 345454
rect 491926 345218 491968 345454
rect 491648 345134 491968 345218
rect 491648 344898 491690 345134
rect 491926 344898 491968 345134
rect 491648 344866 491968 344898
rect 522368 345454 522688 345486
rect 522368 345218 522410 345454
rect 522646 345218 522688 345454
rect 522368 345134 522688 345218
rect 522368 344898 522410 345134
rect 522646 344898 522688 345134
rect 522368 344866 522688 344898
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 46208 327454 46528 327486
rect 46208 327218 46250 327454
rect 46486 327218 46528 327454
rect 46208 327134 46528 327218
rect 46208 326898 46250 327134
rect 46486 326898 46528 327134
rect 46208 326866 46528 326898
rect 76928 327454 77248 327486
rect 76928 327218 76970 327454
rect 77206 327218 77248 327454
rect 76928 327134 77248 327218
rect 76928 326898 76970 327134
rect 77206 326898 77248 327134
rect 76928 326866 77248 326898
rect 107648 327454 107968 327486
rect 107648 327218 107690 327454
rect 107926 327218 107968 327454
rect 107648 327134 107968 327218
rect 107648 326898 107690 327134
rect 107926 326898 107968 327134
rect 107648 326866 107968 326898
rect 138368 327454 138688 327486
rect 138368 327218 138410 327454
rect 138646 327218 138688 327454
rect 138368 327134 138688 327218
rect 138368 326898 138410 327134
rect 138646 326898 138688 327134
rect 138368 326866 138688 326898
rect 169088 327454 169408 327486
rect 169088 327218 169130 327454
rect 169366 327218 169408 327454
rect 169088 327134 169408 327218
rect 169088 326898 169130 327134
rect 169366 326898 169408 327134
rect 169088 326866 169408 326898
rect 199808 327454 200128 327486
rect 199808 327218 199850 327454
rect 200086 327218 200128 327454
rect 199808 327134 200128 327218
rect 199808 326898 199850 327134
rect 200086 326898 200128 327134
rect 199808 326866 200128 326898
rect 230528 327454 230848 327486
rect 230528 327218 230570 327454
rect 230806 327218 230848 327454
rect 230528 327134 230848 327218
rect 230528 326898 230570 327134
rect 230806 326898 230848 327134
rect 230528 326866 230848 326898
rect 261248 327454 261568 327486
rect 261248 327218 261290 327454
rect 261526 327218 261568 327454
rect 261248 327134 261568 327218
rect 261248 326898 261290 327134
rect 261526 326898 261568 327134
rect 261248 326866 261568 326898
rect 291968 327454 292288 327486
rect 291968 327218 292010 327454
rect 292246 327218 292288 327454
rect 291968 327134 292288 327218
rect 291968 326898 292010 327134
rect 292246 326898 292288 327134
rect 291968 326866 292288 326898
rect 322688 327454 323008 327486
rect 322688 327218 322730 327454
rect 322966 327218 323008 327454
rect 322688 327134 323008 327218
rect 322688 326898 322730 327134
rect 322966 326898 323008 327134
rect 322688 326866 323008 326898
rect 353408 327454 353728 327486
rect 353408 327218 353450 327454
rect 353686 327218 353728 327454
rect 353408 327134 353728 327218
rect 353408 326898 353450 327134
rect 353686 326898 353728 327134
rect 353408 326866 353728 326898
rect 384128 327454 384448 327486
rect 384128 327218 384170 327454
rect 384406 327218 384448 327454
rect 384128 327134 384448 327218
rect 384128 326898 384170 327134
rect 384406 326898 384448 327134
rect 384128 326866 384448 326898
rect 414848 327454 415168 327486
rect 414848 327218 414890 327454
rect 415126 327218 415168 327454
rect 414848 327134 415168 327218
rect 414848 326898 414890 327134
rect 415126 326898 415168 327134
rect 414848 326866 415168 326898
rect 445568 327454 445888 327486
rect 445568 327218 445610 327454
rect 445846 327218 445888 327454
rect 445568 327134 445888 327218
rect 445568 326898 445610 327134
rect 445846 326898 445888 327134
rect 445568 326866 445888 326898
rect 476288 327454 476608 327486
rect 476288 327218 476330 327454
rect 476566 327218 476608 327454
rect 476288 327134 476608 327218
rect 476288 326898 476330 327134
rect 476566 326898 476608 327134
rect 476288 326866 476608 326898
rect 507008 327454 507328 327486
rect 507008 327218 507050 327454
rect 507286 327218 507328 327454
rect 507008 327134 507328 327218
rect 507008 326898 507050 327134
rect 507286 326898 507328 327134
rect 507008 326866 507328 326898
rect 537728 327454 538048 327486
rect 537728 327218 537770 327454
rect 538006 327218 538048 327454
rect 537728 327134 538048 327218
rect 537728 326898 537770 327134
rect 538006 326898 538048 327134
rect 537728 326866 538048 326898
rect 61568 309454 61888 309486
rect 61568 309218 61610 309454
rect 61846 309218 61888 309454
rect 61568 309134 61888 309218
rect 61568 308898 61610 309134
rect 61846 308898 61888 309134
rect 61568 308866 61888 308898
rect 92288 309454 92608 309486
rect 92288 309218 92330 309454
rect 92566 309218 92608 309454
rect 92288 309134 92608 309218
rect 92288 308898 92330 309134
rect 92566 308898 92608 309134
rect 92288 308866 92608 308898
rect 123008 309454 123328 309486
rect 123008 309218 123050 309454
rect 123286 309218 123328 309454
rect 123008 309134 123328 309218
rect 123008 308898 123050 309134
rect 123286 308898 123328 309134
rect 123008 308866 123328 308898
rect 153728 309454 154048 309486
rect 153728 309218 153770 309454
rect 154006 309218 154048 309454
rect 153728 309134 154048 309218
rect 153728 308898 153770 309134
rect 154006 308898 154048 309134
rect 153728 308866 154048 308898
rect 184448 309454 184768 309486
rect 184448 309218 184490 309454
rect 184726 309218 184768 309454
rect 184448 309134 184768 309218
rect 184448 308898 184490 309134
rect 184726 308898 184768 309134
rect 184448 308866 184768 308898
rect 215168 309454 215488 309486
rect 215168 309218 215210 309454
rect 215446 309218 215488 309454
rect 215168 309134 215488 309218
rect 215168 308898 215210 309134
rect 215446 308898 215488 309134
rect 215168 308866 215488 308898
rect 245888 309454 246208 309486
rect 245888 309218 245930 309454
rect 246166 309218 246208 309454
rect 245888 309134 246208 309218
rect 245888 308898 245930 309134
rect 246166 308898 246208 309134
rect 245888 308866 246208 308898
rect 276608 309454 276928 309486
rect 276608 309218 276650 309454
rect 276886 309218 276928 309454
rect 276608 309134 276928 309218
rect 276608 308898 276650 309134
rect 276886 308898 276928 309134
rect 276608 308866 276928 308898
rect 307328 309454 307648 309486
rect 307328 309218 307370 309454
rect 307606 309218 307648 309454
rect 307328 309134 307648 309218
rect 307328 308898 307370 309134
rect 307606 308898 307648 309134
rect 307328 308866 307648 308898
rect 338048 309454 338368 309486
rect 338048 309218 338090 309454
rect 338326 309218 338368 309454
rect 338048 309134 338368 309218
rect 338048 308898 338090 309134
rect 338326 308898 338368 309134
rect 338048 308866 338368 308898
rect 368768 309454 369088 309486
rect 368768 309218 368810 309454
rect 369046 309218 369088 309454
rect 368768 309134 369088 309218
rect 368768 308898 368810 309134
rect 369046 308898 369088 309134
rect 368768 308866 369088 308898
rect 399488 309454 399808 309486
rect 399488 309218 399530 309454
rect 399766 309218 399808 309454
rect 399488 309134 399808 309218
rect 399488 308898 399530 309134
rect 399766 308898 399808 309134
rect 399488 308866 399808 308898
rect 430208 309454 430528 309486
rect 430208 309218 430250 309454
rect 430486 309218 430528 309454
rect 430208 309134 430528 309218
rect 430208 308898 430250 309134
rect 430486 308898 430528 309134
rect 430208 308866 430528 308898
rect 460928 309454 461248 309486
rect 460928 309218 460970 309454
rect 461206 309218 461248 309454
rect 460928 309134 461248 309218
rect 460928 308898 460970 309134
rect 461206 308898 461248 309134
rect 460928 308866 461248 308898
rect 491648 309454 491968 309486
rect 491648 309218 491690 309454
rect 491926 309218 491968 309454
rect 491648 309134 491968 309218
rect 491648 308898 491690 309134
rect 491926 308898 491968 309134
rect 491648 308866 491968 308898
rect 522368 309454 522688 309486
rect 522368 309218 522410 309454
rect 522646 309218 522688 309454
rect 522368 309134 522688 309218
rect 522368 308898 522410 309134
rect 522646 308898 522688 309134
rect 522368 308866 522688 308898
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 46208 291454 46528 291486
rect 46208 291218 46250 291454
rect 46486 291218 46528 291454
rect 46208 291134 46528 291218
rect 46208 290898 46250 291134
rect 46486 290898 46528 291134
rect 46208 290866 46528 290898
rect 76928 291454 77248 291486
rect 76928 291218 76970 291454
rect 77206 291218 77248 291454
rect 76928 291134 77248 291218
rect 76928 290898 76970 291134
rect 77206 290898 77248 291134
rect 76928 290866 77248 290898
rect 107648 291454 107968 291486
rect 107648 291218 107690 291454
rect 107926 291218 107968 291454
rect 107648 291134 107968 291218
rect 107648 290898 107690 291134
rect 107926 290898 107968 291134
rect 107648 290866 107968 290898
rect 138368 291454 138688 291486
rect 138368 291218 138410 291454
rect 138646 291218 138688 291454
rect 138368 291134 138688 291218
rect 138368 290898 138410 291134
rect 138646 290898 138688 291134
rect 138368 290866 138688 290898
rect 169088 291454 169408 291486
rect 169088 291218 169130 291454
rect 169366 291218 169408 291454
rect 169088 291134 169408 291218
rect 169088 290898 169130 291134
rect 169366 290898 169408 291134
rect 169088 290866 169408 290898
rect 199808 291454 200128 291486
rect 199808 291218 199850 291454
rect 200086 291218 200128 291454
rect 199808 291134 200128 291218
rect 199808 290898 199850 291134
rect 200086 290898 200128 291134
rect 199808 290866 200128 290898
rect 230528 291454 230848 291486
rect 230528 291218 230570 291454
rect 230806 291218 230848 291454
rect 230528 291134 230848 291218
rect 230528 290898 230570 291134
rect 230806 290898 230848 291134
rect 230528 290866 230848 290898
rect 261248 291454 261568 291486
rect 261248 291218 261290 291454
rect 261526 291218 261568 291454
rect 261248 291134 261568 291218
rect 261248 290898 261290 291134
rect 261526 290898 261568 291134
rect 261248 290866 261568 290898
rect 291968 291454 292288 291486
rect 291968 291218 292010 291454
rect 292246 291218 292288 291454
rect 291968 291134 292288 291218
rect 291968 290898 292010 291134
rect 292246 290898 292288 291134
rect 291968 290866 292288 290898
rect 322688 291454 323008 291486
rect 322688 291218 322730 291454
rect 322966 291218 323008 291454
rect 322688 291134 323008 291218
rect 322688 290898 322730 291134
rect 322966 290898 323008 291134
rect 322688 290866 323008 290898
rect 353408 291454 353728 291486
rect 353408 291218 353450 291454
rect 353686 291218 353728 291454
rect 353408 291134 353728 291218
rect 353408 290898 353450 291134
rect 353686 290898 353728 291134
rect 353408 290866 353728 290898
rect 384128 291454 384448 291486
rect 384128 291218 384170 291454
rect 384406 291218 384448 291454
rect 384128 291134 384448 291218
rect 384128 290898 384170 291134
rect 384406 290898 384448 291134
rect 384128 290866 384448 290898
rect 414848 291454 415168 291486
rect 414848 291218 414890 291454
rect 415126 291218 415168 291454
rect 414848 291134 415168 291218
rect 414848 290898 414890 291134
rect 415126 290898 415168 291134
rect 414848 290866 415168 290898
rect 445568 291454 445888 291486
rect 445568 291218 445610 291454
rect 445846 291218 445888 291454
rect 445568 291134 445888 291218
rect 445568 290898 445610 291134
rect 445846 290898 445888 291134
rect 445568 290866 445888 290898
rect 476288 291454 476608 291486
rect 476288 291218 476330 291454
rect 476566 291218 476608 291454
rect 476288 291134 476608 291218
rect 476288 290898 476330 291134
rect 476566 290898 476608 291134
rect 476288 290866 476608 290898
rect 507008 291454 507328 291486
rect 507008 291218 507050 291454
rect 507286 291218 507328 291454
rect 507008 291134 507328 291218
rect 507008 290898 507050 291134
rect 507286 290898 507328 291134
rect 507008 290866 507328 290898
rect 537728 291454 538048 291486
rect 537728 291218 537770 291454
rect 538006 291218 538048 291454
rect 537728 291134 538048 291218
rect 537728 290898 537770 291134
rect 538006 290898 538048 291134
rect 537728 290866 538048 290898
rect 61568 273454 61888 273486
rect 61568 273218 61610 273454
rect 61846 273218 61888 273454
rect 61568 273134 61888 273218
rect 61568 272898 61610 273134
rect 61846 272898 61888 273134
rect 61568 272866 61888 272898
rect 92288 273454 92608 273486
rect 92288 273218 92330 273454
rect 92566 273218 92608 273454
rect 92288 273134 92608 273218
rect 92288 272898 92330 273134
rect 92566 272898 92608 273134
rect 92288 272866 92608 272898
rect 123008 273454 123328 273486
rect 123008 273218 123050 273454
rect 123286 273218 123328 273454
rect 123008 273134 123328 273218
rect 123008 272898 123050 273134
rect 123286 272898 123328 273134
rect 123008 272866 123328 272898
rect 153728 273454 154048 273486
rect 153728 273218 153770 273454
rect 154006 273218 154048 273454
rect 153728 273134 154048 273218
rect 153728 272898 153770 273134
rect 154006 272898 154048 273134
rect 153728 272866 154048 272898
rect 184448 273454 184768 273486
rect 184448 273218 184490 273454
rect 184726 273218 184768 273454
rect 184448 273134 184768 273218
rect 184448 272898 184490 273134
rect 184726 272898 184768 273134
rect 184448 272866 184768 272898
rect 215168 273454 215488 273486
rect 215168 273218 215210 273454
rect 215446 273218 215488 273454
rect 215168 273134 215488 273218
rect 215168 272898 215210 273134
rect 215446 272898 215488 273134
rect 215168 272866 215488 272898
rect 245888 273454 246208 273486
rect 245888 273218 245930 273454
rect 246166 273218 246208 273454
rect 245888 273134 246208 273218
rect 245888 272898 245930 273134
rect 246166 272898 246208 273134
rect 245888 272866 246208 272898
rect 276608 273454 276928 273486
rect 276608 273218 276650 273454
rect 276886 273218 276928 273454
rect 276608 273134 276928 273218
rect 276608 272898 276650 273134
rect 276886 272898 276928 273134
rect 276608 272866 276928 272898
rect 307328 273454 307648 273486
rect 307328 273218 307370 273454
rect 307606 273218 307648 273454
rect 307328 273134 307648 273218
rect 307328 272898 307370 273134
rect 307606 272898 307648 273134
rect 307328 272866 307648 272898
rect 338048 273454 338368 273486
rect 338048 273218 338090 273454
rect 338326 273218 338368 273454
rect 338048 273134 338368 273218
rect 338048 272898 338090 273134
rect 338326 272898 338368 273134
rect 338048 272866 338368 272898
rect 368768 273454 369088 273486
rect 368768 273218 368810 273454
rect 369046 273218 369088 273454
rect 368768 273134 369088 273218
rect 368768 272898 368810 273134
rect 369046 272898 369088 273134
rect 368768 272866 369088 272898
rect 399488 273454 399808 273486
rect 399488 273218 399530 273454
rect 399766 273218 399808 273454
rect 399488 273134 399808 273218
rect 399488 272898 399530 273134
rect 399766 272898 399808 273134
rect 399488 272866 399808 272898
rect 430208 273454 430528 273486
rect 430208 273218 430250 273454
rect 430486 273218 430528 273454
rect 430208 273134 430528 273218
rect 430208 272898 430250 273134
rect 430486 272898 430528 273134
rect 430208 272866 430528 272898
rect 460928 273454 461248 273486
rect 460928 273218 460970 273454
rect 461206 273218 461248 273454
rect 460928 273134 461248 273218
rect 460928 272898 460970 273134
rect 461206 272898 461248 273134
rect 460928 272866 461248 272898
rect 491648 273454 491968 273486
rect 491648 273218 491690 273454
rect 491926 273218 491968 273454
rect 491648 273134 491968 273218
rect 491648 272898 491690 273134
rect 491926 272898 491968 273134
rect 491648 272866 491968 272898
rect 522368 273454 522688 273486
rect 522368 273218 522410 273454
rect 522646 273218 522688 273454
rect 522368 273134 522688 273218
rect 522368 272898 522410 273134
rect 522646 272898 522688 273134
rect 522368 272866 522688 272898
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 46208 255454 46528 255486
rect 46208 255218 46250 255454
rect 46486 255218 46528 255454
rect 46208 255134 46528 255218
rect 46208 254898 46250 255134
rect 46486 254898 46528 255134
rect 46208 254866 46528 254898
rect 76928 255454 77248 255486
rect 76928 255218 76970 255454
rect 77206 255218 77248 255454
rect 76928 255134 77248 255218
rect 76928 254898 76970 255134
rect 77206 254898 77248 255134
rect 76928 254866 77248 254898
rect 107648 255454 107968 255486
rect 107648 255218 107690 255454
rect 107926 255218 107968 255454
rect 107648 255134 107968 255218
rect 107648 254898 107690 255134
rect 107926 254898 107968 255134
rect 107648 254866 107968 254898
rect 138368 255454 138688 255486
rect 138368 255218 138410 255454
rect 138646 255218 138688 255454
rect 138368 255134 138688 255218
rect 138368 254898 138410 255134
rect 138646 254898 138688 255134
rect 138368 254866 138688 254898
rect 169088 255454 169408 255486
rect 169088 255218 169130 255454
rect 169366 255218 169408 255454
rect 169088 255134 169408 255218
rect 169088 254898 169130 255134
rect 169366 254898 169408 255134
rect 169088 254866 169408 254898
rect 199808 255454 200128 255486
rect 199808 255218 199850 255454
rect 200086 255218 200128 255454
rect 199808 255134 200128 255218
rect 199808 254898 199850 255134
rect 200086 254898 200128 255134
rect 199808 254866 200128 254898
rect 230528 255454 230848 255486
rect 230528 255218 230570 255454
rect 230806 255218 230848 255454
rect 230528 255134 230848 255218
rect 230528 254898 230570 255134
rect 230806 254898 230848 255134
rect 230528 254866 230848 254898
rect 261248 255454 261568 255486
rect 261248 255218 261290 255454
rect 261526 255218 261568 255454
rect 261248 255134 261568 255218
rect 261248 254898 261290 255134
rect 261526 254898 261568 255134
rect 261248 254866 261568 254898
rect 291968 255454 292288 255486
rect 291968 255218 292010 255454
rect 292246 255218 292288 255454
rect 291968 255134 292288 255218
rect 291968 254898 292010 255134
rect 292246 254898 292288 255134
rect 291968 254866 292288 254898
rect 322688 255454 323008 255486
rect 322688 255218 322730 255454
rect 322966 255218 323008 255454
rect 322688 255134 323008 255218
rect 322688 254898 322730 255134
rect 322966 254898 323008 255134
rect 322688 254866 323008 254898
rect 353408 255454 353728 255486
rect 353408 255218 353450 255454
rect 353686 255218 353728 255454
rect 353408 255134 353728 255218
rect 353408 254898 353450 255134
rect 353686 254898 353728 255134
rect 353408 254866 353728 254898
rect 384128 255454 384448 255486
rect 384128 255218 384170 255454
rect 384406 255218 384448 255454
rect 384128 255134 384448 255218
rect 384128 254898 384170 255134
rect 384406 254898 384448 255134
rect 384128 254866 384448 254898
rect 414848 255454 415168 255486
rect 414848 255218 414890 255454
rect 415126 255218 415168 255454
rect 414848 255134 415168 255218
rect 414848 254898 414890 255134
rect 415126 254898 415168 255134
rect 414848 254866 415168 254898
rect 445568 255454 445888 255486
rect 445568 255218 445610 255454
rect 445846 255218 445888 255454
rect 445568 255134 445888 255218
rect 445568 254898 445610 255134
rect 445846 254898 445888 255134
rect 445568 254866 445888 254898
rect 476288 255454 476608 255486
rect 476288 255218 476330 255454
rect 476566 255218 476608 255454
rect 476288 255134 476608 255218
rect 476288 254898 476330 255134
rect 476566 254898 476608 255134
rect 476288 254866 476608 254898
rect 507008 255454 507328 255486
rect 507008 255218 507050 255454
rect 507286 255218 507328 255454
rect 507008 255134 507328 255218
rect 507008 254898 507050 255134
rect 507286 254898 507328 255134
rect 507008 254866 507328 254898
rect 537728 255454 538048 255486
rect 537728 255218 537770 255454
rect 538006 255218 538048 255454
rect 537728 255134 538048 255218
rect 537728 254898 537770 255134
rect 538006 254898 538048 255134
rect 537728 254866 538048 254898
rect 61568 237454 61888 237486
rect 61568 237218 61610 237454
rect 61846 237218 61888 237454
rect 61568 237134 61888 237218
rect 61568 236898 61610 237134
rect 61846 236898 61888 237134
rect 61568 236866 61888 236898
rect 92288 237454 92608 237486
rect 92288 237218 92330 237454
rect 92566 237218 92608 237454
rect 92288 237134 92608 237218
rect 92288 236898 92330 237134
rect 92566 236898 92608 237134
rect 92288 236866 92608 236898
rect 123008 237454 123328 237486
rect 123008 237218 123050 237454
rect 123286 237218 123328 237454
rect 123008 237134 123328 237218
rect 123008 236898 123050 237134
rect 123286 236898 123328 237134
rect 123008 236866 123328 236898
rect 153728 237454 154048 237486
rect 153728 237218 153770 237454
rect 154006 237218 154048 237454
rect 153728 237134 154048 237218
rect 153728 236898 153770 237134
rect 154006 236898 154048 237134
rect 153728 236866 154048 236898
rect 184448 237454 184768 237486
rect 184448 237218 184490 237454
rect 184726 237218 184768 237454
rect 184448 237134 184768 237218
rect 184448 236898 184490 237134
rect 184726 236898 184768 237134
rect 184448 236866 184768 236898
rect 215168 237454 215488 237486
rect 215168 237218 215210 237454
rect 215446 237218 215488 237454
rect 215168 237134 215488 237218
rect 215168 236898 215210 237134
rect 215446 236898 215488 237134
rect 215168 236866 215488 236898
rect 245888 237454 246208 237486
rect 245888 237218 245930 237454
rect 246166 237218 246208 237454
rect 245888 237134 246208 237218
rect 245888 236898 245930 237134
rect 246166 236898 246208 237134
rect 245888 236866 246208 236898
rect 276608 237454 276928 237486
rect 276608 237218 276650 237454
rect 276886 237218 276928 237454
rect 276608 237134 276928 237218
rect 276608 236898 276650 237134
rect 276886 236898 276928 237134
rect 276608 236866 276928 236898
rect 307328 237454 307648 237486
rect 307328 237218 307370 237454
rect 307606 237218 307648 237454
rect 307328 237134 307648 237218
rect 307328 236898 307370 237134
rect 307606 236898 307648 237134
rect 307328 236866 307648 236898
rect 338048 237454 338368 237486
rect 338048 237218 338090 237454
rect 338326 237218 338368 237454
rect 338048 237134 338368 237218
rect 338048 236898 338090 237134
rect 338326 236898 338368 237134
rect 338048 236866 338368 236898
rect 368768 237454 369088 237486
rect 368768 237218 368810 237454
rect 369046 237218 369088 237454
rect 368768 237134 369088 237218
rect 368768 236898 368810 237134
rect 369046 236898 369088 237134
rect 368768 236866 369088 236898
rect 399488 237454 399808 237486
rect 399488 237218 399530 237454
rect 399766 237218 399808 237454
rect 399488 237134 399808 237218
rect 399488 236898 399530 237134
rect 399766 236898 399808 237134
rect 399488 236866 399808 236898
rect 430208 237454 430528 237486
rect 430208 237218 430250 237454
rect 430486 237218 430528 237454
rect 430208 237134 430528 237218
rect 430208 236898 430250 237134
rect 430486 236898 430528 237134
rect 430208 236866 430528 236898
rect 460928 237454 461248 237486
rect 460928 237218 460970 237454
rect 461206 237218 461248 237454
rect 460928 237134 461248 237218
rect 460928 236898 460970 237134
rect 461206 236898 461248 237134
rect 460928 236866 461248 236898
rect 491648 237454 491968 237486
rect 491648 237218 491690 237454
rect 491926 237218 491968 237454
rect 491648 237134 491968 237218
rect 491648 236898 491690 237134
rect 491926 236898 491968 237134
rect 491648 236866 491968 236898
rect 522368 237454 522688 237486
rect 522368 237218 522410 237454
rect 522646 237218 522688 237454
rect 522368 237134 522688 237218
rect 522368 236898 522410 237134
rect 522646 236898 522688 237134
rect 522368 236866 522688 236898
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 46208 219454 46528 219486
rect 46208 219218 46250 219454
rect 46486 219218 46528 219454
rect 46208 219134 46528 219218
rect 46208 218898 46250 219134
rect 46486 218898 46528 219134
rect 46208 218866 46528 218898
rect 76928 219454 77248 219486
rect 76928 219218 76970 219454
rect 77206 219218 77248 219454
rect 76928 219134 77248 219218
rect 76928 218898 76970 219134
rect 77206 218898 77248 219134
rect 76928 218866 77248 218898
rect 107648 219454 107968 219486
rect 107648 219218 107690 219454
rect 107926 219218 107968 219454
rect 107648 219134 107968 219218
rect 107648 218898 107690 219134
rect 107926 218898 107968 219134
rect 107648 218866 107968 218898
rect 138368 219454 138688 219486
rect 138368 219218 138410 219454
rect 138646 219218 138688 219454
rect 138368 219134 138688 219218
rect 138368 218898 138410 219134
rect 138646 218898 138688 219134
rect 138368 218866 138688 218898
rect 169088 219454 169408 219486
rect 169088 219218 169130 219454
rect 169366 219218 169408 219454
rect 169088 219134 169408 219218
rect 169088 218898 169130 219134
rect 169366 218898 169408 219134
rect 169088 218866 169408 218898
rect 199808 219454 200128 219486
rect 199808 219218 199850 219454
rect 200086 219218 200128 219454
rect 199808 219134 200128 219218
rect 199808 218898 199850 219134
rect 200086 218898 200128 219134
rect 199808 218866 200128 218898
rect 230528 219454 230848 219486
rect 230528 219218 230570 219454
rect 230806 219218 230848 219454
rect 230528 219134 230848 219218
rect 230528 218898 230570 219134
rect 230806 218898 230848 219134
rect 230528 218866 230848 218898
rect 261248 219454 261568 219486
rect 261248 219218 261290 219454
rect 261526 219218 261568 219454
rect 261248 219134 261568 219218
rect 261248 218898 261290 219134
rect 261526 218898 261568 219134
rect 261248 218866 261568 218898
rect 291968 219454 292288 219486
rect 291968 219218 292010 219454
rect 292246 219218 292288 219454
rect 291968 219134 292288 219218
rect 291968 218898 292010 219134
rect 292246 218898 292288 219134
rect 291968 218866 292288 218898
rect 322688 219454 323008 219486
rect 322688 219218 322730 219454
rect 322966 219218 323008 219454
rect 322688 219134 323008 219218
rect 322688 218898 322730 219134
rect 322966 218898 323008 219134
rect 322688 218866 323008 218898
rect 353408 219454 353728 219486
rect 353408 219218 353450 219454
rect 353686 219218 353728 219454
rect 353408 219134 353728 219218
rect 353408 218898 353450 219134
rect 353686 218898 353728 219134
rect 353408 218866 353728 218898
rect 384128 219454 384448 219486
rect 384128 219218 384170 219454
rect 384406 219218 384448 219454
rect 384128 219134 384448 219218
rect 384128 218898 384170 219134
rect 384406 218898 384448 219134
rect 384128 218866 384448 218898
rect 414848 219454 415168 219486
rect 414848 219218 414890 219454
rect 415126 219218 415168 219454
rect 414848 219134 415168 219218
rect 414848 218898 414890 219134
rect 415126 218898 415168 219134
rect 414848 218866 415168 218898
rect 445568 219454 445888 219486
rect 445568 219218 445610 219454
rect 445846 219218 445888 219454
rect 445568 219134 445888 219218
rect 445568 218898 445610 219134
rect 445846 218898 445888 219134
rect 445568 218866 445888 218898
rect 476288 219454 476608 219486
rect 476288 219218 476330 219454
rect 476566 219218 476608 219454
rect 476288 219134 476608 219218
rect 476288 218898 476330 219134
rect 476566 218898 476608 219134
rect 476288 218866 476608 218898
rect 507008 219454 507328 219486
rect 507008 219218 507050 219454
rect 507286 219218 507328 219454
rect 507008 219134 507328 219218
rect 507008 218898 507050 219134
rect 507286 218898 507328 219134
rect 507008 218866 507328 218898
rect 537728 219454 538048 219486
rect 537728 219218 537770 219454
rect 538006 219218 538048 219454
rect 537728 219134 538048 219218
rect 537728 218898 537770 219134
rect 538006 218898 538048 219134
rect 537728 218866 538048 218898
rect 61568 201454 61888 201486
rect 61568 201218 61610 201454
rect 61846 201218 61888 201454
rect 61568 201134 61888 201218
rect 61568 200898 61610 201134
rect 61846 200898 61888 201134
rect 61568 200866 61888 200898
rect 92288 201454 92608 201486
rect 92288 201218 92330 201454
rect 92566 201218 92608 201454
rect 92288 201134 92608 201218
rect 92288 200898 92330 201134
rect 92566 200898 92608 201134
rect 92288 200866 92608 200898
rect 123008 201454 123328 201486
rect 123008 201218 123050 201454
rect 123286 201218 123328 201454
rect 123008 201134 123328 201218
rect 123008 200898 123050 201134
rect 123286 200898 123328 201134
rect 123008 200866 123328 200898
rect 153728 201454 154048 201486
rect 153728 201218 153770 201454
rect 154006 201218 154048 201454
rect 153728 201134 154048 201218
rect 153728 200898 153770 201134
rect 154006 200898 154048 201134
rect 153728 200866 154048 200898
rect 184448 201454 184768 201486
rect 184448 201218 184490 201454
rect 184726 201218 184768 201454
rect 184448 201134 184768 201218
rect 184448 200898 184490 201134
rect 184726 200898 184768 201134
rect 184448 200866 184768 200898
rect 215168 201454 215488 201486
rect 215168 201218 215210 201454
rect 215446 201218 215488 201454
rect 215168 201134 215488 201218
rect 215168 200898 215210 201134
rect 215446 200898 215488 201134
rect 215168 200866 215488 200898
rect 245888 201454 246208 201486
rect 245888 201218 245930 201454
rect 246166 201218 246208 201454
rect 245888 201134 246208 201218
rect 245888 200898 245930 201134
rect 246166 200898 246208 201134
rect 245888 200866 246208 200898
rect 276608 201454 276928 201486
rect 276608 201218 276650 201454
rect 276886 201218 276928 201454
rect 276608 201134 276928 201218
rect 276608 200898 276650 201134
rect 276886 200898 276928 201134
rect 276608 200866 276928 200898
rect 307328 201454 307648 201486
rect 307328 201218 307370 201454
rect 307606 201218 307648 201454
rect 307328 201134 307648 201218
rect 307328 200898 307370 201134
rect 307606 200898 307648 201134
rect 307328 200866 307648 200898
rect 338048 201454 338368 201486
rect 338048 201218 338090 201454
rect 338326 201218 338368 201454
rect 338048 201134 338368 201218
rect 338048 200898 338090 201134
rect 338326 200898 338368 201134
rect 338048 200866 338368 200898
rect 368768 201454 369088 201486
rect 368768 201218 368810 201454
rect 369046 201218 369088 201454
rect 368768 201134 369088 201218
rect 368768 200898 368810 201134
rect 369046 200898 369088 201134
rect 368768 200866 369088 200898
rect 399488 201454 399808 201486
rect 399488 201218 399530 201454
rect 399766 201218 399808 201454
rect 399488 201134 399808 201218
rect 399488 200898 399530 201134
rect 399766 200898 399808 201134
rect 399488 200866 399808 200898
rect 430208 201454 430528 201486
rect 430208 201218 430250 201454
rect 430486 201218 430528 201454
rect 430208 201134 430528 201218
rect 430208 200898 430250 201134
rect 430486 200898 430528 201134
rect 430208 200866 430528 200898
rect 460928 201454 461248 201486
rect 460928 201218 460970 201454
rect 461206 201218 461248 201454
rect 460928 201134 461248 201218
rect 460928 200898 460970 201134
rect 461206 200898 461248 201134
rect 460928 200866 461248 200898
rect 491648 201454 491968 201486
rect 491648 201218 491690 201454
rect 491926 201218 491968 201454
rect 491648 201134 491968 201218
rect 491648 200898 491690 201134
rect 491926 200898 491968 201134
rect 491648 200866 491968 200898
rect 522368 201454 522688 201486
rect 522368 201218 522410 201454
rect 522646 201218 522688 201454
rect 522368 201134 522688 201218
rect 522368 200898 522410 201134
rect 522646 200898 522688 201134
rect 522368 200866 522688 200898
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 46208 183454 46528 183486
rect 46208 183218 46250 183454
rect 46486 183218 46528 183454
rect 46208 183134 46528 183218
rect 46208 182898 46250 183134
rect 46486 182898 46528 183134
rect 46208 182866 46528 182898
rect 76928 183454 77248 183486
rect 76928 183218 76970 183454
rect 77206 183218 77248 183454
rect 76928 183134 77248 183218
rect 76928 182898 76970 183134
rect 77206 182898 77248 183134
rect 76928 182866 77248 182898
rect 107648 183454 107968 183486
rect 107648 183218 107690 183454
rect 107926 183218 107968 183454
rect 107648 183134 107968 183218
rect 107648 182898 107690 183134
rect 107926 182898 107968 183134
rect 107648 182866 107968 182898
rect 138368 183454 138688 183486
rect 138368 183218 138410 183454
rect 138646 183218 138688 183454
rect 138368 183134 138688 183218
rect 138368 182898 138410 183134
rect 138646 182898 138688 183134
rect 138368 182866 138688 182898
rect 169088 183454 169408 183486
rect 169088 183218 169130 183454
rect 169366 183218 169408 183454
rect 169088 183134 169408 183218
rect 169088 182898 169130 183134
rect 169366 182898 169408 183134
rect 169088 182866 169408 182898
rect 199808 183454 200128 183486
rect 199808 183218 199850 183454
rect 200086 183218 200128 183454
rect 199808 183134 200128 183218
rect 199808 182898 199850 183134
rect 200086 182898 200128 183134
rect 199808 182866 200128 182898
rect 230528 183454 230848 183486
rect 230528 183218 230570 183454
rect 230806 183218 230848 183454
rect 230528 183134 230848 183218
rect 230528 182898 230570 183134
rect 230806 182898 230848 183134
rect 230528 182866 230848 182898
rect 261248 183454 261568 183486
rect 261248 183218 261290 183454
rect 261526 183218 261568 183454
rect 261248 183134 261568 183218
rect 261248 182898 261290 183134
rect 261526 182898 261568 183134
rect 261248 182866 261568 182898
rect 291968 183454 292288 183486
rect 291968 183218 292010 183454
rect 292246 183218 292288 183454
rect 291968 183134 292288 183218
rect 291968 182898 292010 183134
rect 292246 182898 292288 183134
rect 291968 182866 292288 182898
rect 322688 183454 323008 183486
rect 322688 183218 322730 183454
rect 322966 183218 323008 183454
rect 322688 183134 323008 183218
rect 322688 182898 322730 183134
rect 322966 182898 323008 183134
rect 322688 182866 323008 182898
rect 353408 183454 353728 183486
rect 353408 183218 353450 183454
rect 353686 183218 353728 183454
rect 353408 183134 353728 183218
rect 353408 182898 353450 183134
rect 353686 182898 353728 183134
rect 353408 182866 353728 182898
rect 384128 183454 384448 183486
rect 384128 183218 384170 183454
rect 384406 183218 384448 183454
rect 384128 183134 384448 183218
rect 384128 182898 384170 183134
rect 384406 182898 384448 183134
rect 384128 182866 384448 182898
rect 414848 183454 415168 183486
rect 414848 183218 414890 183454
rect 415126 183218 415168 183454
rect 414848 183134 415168 183218
rect 414848 182898 414890 183134
rect 415126 182898 415168 183134
rect 414848 182866 415168 182898
rect 445568 183454 445888 183486
rect 445568 183218 445610 183454
rect 445846 183218 445888 183454
rect 445568 183134 445888 183218
rect 445568 182898 445610 183134
rect 445846 182898 445888 183134
rect 445568 182866 445888 182898
rect 476288 183454 476608 183486
rect 476288 183218 476330 183454
rect 476566 183218 476608 183454
rect 476288 183134 476608 183218
rect 476288 182898 476330 183134
rect 476566 182898 476608 183134
rect 476288 182866 476608 182898
rect 507008 183454 507328 183486
rect 507008 183218 507050 183454
rect 507286 183218 507328 183454
rect 507008 183134 507328 183218
rect 507008 182898 507050 183134
rect 507286 182898 507328 183134
rect 507008 182866 507328 182898
rect 537728 183454 538048 183486
rect 537728 183218 537770 183454
rect 538006 183218 538048 183454
rect 537728 183134 538048 183218
rect 537728 182898 537770 183134
rect 538006 182898 538048 183134
rect 537728 182866 538048 182898
rect 61568 165454 61888 165486
rect 61568 165218 61610 165454
rect 61846 165218 61888 165454
rect 61568 165134 61888 165218
rect 61568 164898 61610 165134
rect 61846 164898 61888 165134
rect 61568 164866 61888 164898
rect 92288 165454 92608 165486
rect 92288 165218 92330 165454
rect 92566 165218 92608 165454
rect 92288 165134 92608 165218
rect 92288 164898 92330 165134
rect 92566 164898 92608 165134
rect 92288 164866 92608 164898
rect 123008 165454 123328 165486
rect 123008 165218 123050 165454
rect 123286 165218 123328 165454
rect 123008 165134 123328 165218
rect 123008 164898 123050 165134
rect 123286 164898 123328 165134
rect 123008 164866 123328 164898
rect 153728 165454 154048 165486
rect 153728 165218 153770 165454
rect 154006 165218 154048 165454
rect 153728 165134 154048 165218
rect 153728 164898 153770 165134
rect 154006 164898 154048 165134
rect 153728 164866 154048 164898
rect 184448 165454 184768 165486
rect 184448 165218 184490 165454
rect 184726 165218 184768 165454
rect 184448 165134 184768 165218
rect 184448 164898 184490 165134
rect 184726 164898 184768 165134
rect 184448 164866 184768 164898
rect 215168 165454 215488 165486
rect 215168 165218 215210 165454
rect 215446 165218 215488 165454
rect 215168 165134 215488 165218
rect 215168 164898 215210 165134
rect 215446 164898 215488 165134
rect 215168 164866 215488 164898
rect 245888 165454 246208 165486
rect 245888 165218 245930 165454
rect 246166 165218 246208 165454
rect 245888 165134 246208 165218
rect 245888 164898 245930 165134
rect 246166 164898 246208 165134
rect 245888 164866 246208 164898
rect 276608 165454 276928 165486
rect 276608 165218 276650 165454
rect 276886 165218 276928 165454
rect 276608 165134 276928 165218
rect 276608 164898 276650 165134
rect 276886 164898 276928 165134
rect 276608 164866 276928 164898
rect 307328 165454 307648 165486
rect 307328 165218 307370 165454
rect 307606 165218 307648 165454
rect 307328 165134 307648 165218
rect 307328 164898 307370 165134
rect 307606 164898 307648 165134
rect 307328 164866 307648 164898
rect 338048 165454 338368 165486
rect 338048 165218 338090 165454
rect 338326 165218 338368 165454
rect 338048 165134 338368 165218
rect 338048 164898 338090 165134
rect 338326 164898 338368 165134
rect 338048 164866 338368 164898
rect 368768 165454 369088 165486
rect 368768 165218 368810 165454
rect 369046 165218 369088 165454
rect 368768 165134 369088 165218
rect 368768 164898 368810 165134
rect 369046 164898 369088 165134
rect 368768 164866 369088 164898
rect 399488 165454 399808 165486
rect 399488 165218 399530 165454
rect 399766 165218 399808 165454
rect 399488 165134 399808 165218
rect 399488 164898 399530 165134
rect 399766 164898 399808 165134
rect 399488 164866 399808 164898
rect 430208 165454 430528 165486
rect 430208 165218 430250 165454
rect 430486 165218 430528 165454
rect 430208 165134 430528 165218
rect 430208 164898 430250 165134
rect 430486 164898 430528 165134
rect 430208 164866 430528 164898
rect 460928 165454 461248 165486
rect 460928 165218 460970 165454
rect 461206 165218 461248 165454
rect 460928 165134 461248 165218
rect 460928 164898 460970 165134
rect 461206 164898 461248 165134
rect 460928 164866 461248 164898
rect 491648 165454 491968 165486
rect 491648 165218 491690 165454
rect 491926 165218 491968 165454
rect 491648 165134 491968 165218
rect 491648 164898 491690 165134
rect 491926 164898 491968 165134
rect 491648 164866 491968 164898
rect 522368 165454 522688 165486
rect 522368 165218 522410 165454
rect 522646 165218 522688 165454
rect 522368 165134 522688 165218
rect 522368 164898 522410 165134
rect 522646 164898 522688 165134
rect 522368 164866 522688 164898
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 46208 147454 46528 147486
rect 46208 147218 46250 147454
rect 46486 147218 46528 147454
rect 46208 147134 46528 147218
rect 46208 146898 46250 147134
rect 46486 146898 46528 147134
rect 46208 146866 46528 146898
rect 76928 147454 77248 147486
rect 76928 147218 76970 147454
rect 77206 147218 77248 147454
rect 76928 147134 77248 147218
rect 76928 146898 76970 147134
rect 77206 146898 77248 147134
rect 76928 146866 77248 146898
rect 107648 147454 107968 147486
rect 107648 147218 107690 147454
rect 107926 147218 107968 147454
rect 107648 147134 107968 147218
rect 107648 146898 107690 147134
rect 107926 146898 107968 147134
rect 107648 146866 107968 146898
rect 138368 147454 138688 147486
rect 138368 147218 138410 147454
rect 138646 147218 138688 147454
rect 138368 147134 138688 147218
rect 138368 146898 138410 147134
rect 138646 146898 138688 147134
rect 138368 146866 138688 146898
rect 169088 147454 169408 147486
rect 169088 147218 169130 147454
rect 169366 147218 169408 147454
rect 169088 147134 169408 147218
rect 169088 146898 169130 147134
rect 169366 146898 169408 147134
rect 169088 146866 169408 146898
rect 199808 147454 200128 147486
rect 199808 147218 199850 147454
rect 200086 147218 200128 147454
rect 199808 147134 200128 147218
rect 199808 146898 199850 147134
rect 200086 146898 200128 147134
rect 199808 146866 200128 146898
rect 230528 147454 230848 147486
rect 230528 147218 230570 147454
rect 230806 147218 230848 147454
rect 230528 147134 230848 147218
rect 230528 146898 230570 147134
rect 230806 146898 230848 147134
rect 230528 146866 230848 146898
rect 261248 147454 261568 147486
rect 261248 147218 261290 147454
rect 261526 147218 261568 147454
rect 261248 147134 261568 147218
rect 261248 146898 261290 147134
rect 261526 146898 261568 147134
rect 261248 146866 261568 146898
rect 291968 147454 292288 147486
rect 291968 147218 292010 147454
rect 292246 147218 292288 147454
rect 291968 147134 292288 147218
rect 291968 146898 292010 147134
rect 292246 146898 292288 147134
rect 291968 146866 292288 146898
rect 322688 147454 323008 147486
rect 322688 147218 322730 147454
rect 322966 147218 323008 147454
rect 322688 147134 323008 147218
rect 322688 146898 322730 147134
rect 322966 146898 323008 147134
rect 322688 146866 323008 146898
rect 353408 147454 353728 147486
rect 353408 147218 353450 147454
rect 353686 147218 353728 147454
rect 353408 147134 353728 147218
rect 353408 146898 353450 147134
rect 353686 146898 353728 147134
rect 353408 146866 353728 146898
rect 384128 147454 384448 147486
rect 384128 147218 384170 147454
rect 384406 147218 384448 147454
rect 384128 147134 384448 147218
rect 384128 146898 384170 147134
rect 384406 146898 384448 147134
rect 384128 146866 384448 146898
rect 414848 147454 415168 147486
rect 414848 147218 414890 147454
rect 415126 147218 415168 147454
rect 414848 147134 415168 147218
rect 414848 146898 414890 147134
rect 415126 146898 415168 147134
rect 414848 146866 415168 146898
rect 445568 147454 445888 147486
rect 445568 147218 445610 147454
rect 445846 147218 445888 147454
rect 445568 147134 445888 147218
rect 445568 146898 445610 147134
rect 445846 146898 445888 147134
rect 445568 146866 445888 146898
rect 476288 147454 476608 147486
rect 476288 147218 476330 147454
rect 476566 147218 476608 147454
rect 476288 147134 476608 147218
rect 476288 146898 476330 147134
rect 476566 146898 476608 147134
rect 476288 146866 476608 146898
rect 507008 147454 507328 147486
rect 507008 147218 507050 147454
rect 507286 147218 507328 147454
rect 507008 147134 507328 147218
rect 507008 146898 507050 147134
rect 507286 146898 507328 147134
rect 507008 146866 507328 146898
rect 537728 147454 538048 147486
rect 537728 147218 537770 147454
rect 538006 147218 538048 147454
rect 537728 147134 538048 147218
rect 537728 146898 537770 147134
rect 538006 146898 538048 147134
rect 537728 146866 538048 146898
rect 61568 129454 61888 129486
rect 61568 129218 61610 129454
rect 61846 129218 61888 129454
rect 61568 129134 61888 129218
rect 61568 128898 61610 129134
rect 61846 128898 61888 129134
rect 61568 128866 61888 128898
rect 92288 129454 92608 129486
rect 92288 129218 92330 129454
rect 92566 129218 92608 129454
rect 92288 129134 92608 129218
rect 92288 128898 92330 129134
rect 92566 128898 92608 129134
rect 92288 128866 92608 128898
rect 123008 129454 123328 129486
rect 123008 129218 123050 129454
rect 123286 129218 123328 129454
rect 123008 129134 123328 129218
rect 123008 128898 123050 129134
rect 123286 128898 123328 129134
rect 123008 128866 123328 128898
rect 153728 129454 154048 129486
rect 153728 129218 153770 129454
rect 154006 129218 154048 129454
rect 153728 129134 154048 129218
rect 153728 128898 153770 129134
rect 154006 128898 154048 129134
rect 153728 128866 154048 128898
rect 184448 129454 184768 129486
rect 184448 129218 184490 129454
rect 184726 129218 184768 129454
rect 184448 129134 184768 129218
rect 184448 128898 184490 129134
rect 184726 128898 184768 129134
rect 184448 128866 184768 128898
rect 215168 129454 215488 129486
rect 215168 129218 215210 129454
rect 215446 129218 215488 129454
rect 215168 129134 215488 129218
rect 215168 128898 215210 129134
rect 215446 128898 215488 129134
rect 215168 128866 215488 128898
rect 245888 129454 246208 129486
rect 245888 129218 245930 129454
rect 246166 129218 246208 129454
rect 245888 129134 246208 129218
rect 245888 128898 245930 129134
rect 246166 128898 246208 129134
rect 245888 128866 246208 128898
rect 276608 129454 276928 129486
rect 276608 129218 276650 129454
rect 276886 129218 276928 129454
rect 276608 129134 276928 129218
rect 276608 128898 276650 129134
rect 276886 128898 276928 129134
rect 276608 128866 276928 128898
rect 307328 129454 307648 129486
rect 307328 129218 307370 129454
rect 307606 129218 307648 129454
rect 307328 129134 307648 129218
rect 307328 128898 307370 129134
rect 307606 128898 307648 129134
rect 307328 128866 307648 128898
rect 338048 129454 338368 129486
rect 338048 129218 338090 129454
rect 338326 129218 338368 129454
rect 338048 129134 338368 129218
rect 338048 128898 338090 129134
rect 338326 128898 338368 129134
rect 338048 128866 338368 128898
rect 368768 129454 369088 129486
rect 368768 129218 368810 129454
rect 369046 129218 369088 129454
rect 368768 129134 369088 129218
rect 368768 128898 368810 129134
rect 369046 128898 369088 129134
rect 368768 128866 369088 128898
rect 399488 129454 399808 129486
rect 399488 129218 399530 129454
rect 399766 129218 399808 129454
rect 399488 129134 399808 129218
rect 399488 128898 399530 129134
rect 399766 128898 399808 129134
rect 399488 128866 399808 128898
rect 430208 129454 430528 129486
rect 430208 129218 430250 129454
rect 430486 129218 430528 129454
rect 430208 129134 430528 129218
rect 430208 128898 430250 129134
rect 430486 128898 430528 129134
rect 430208 128866 430528 128898
rect 460928 129454 461248 129486
rect 460928 129218 460970 129454
rect 461206 129218 461248 129454
rect 460928 129134 461248 129218
rect 460928 128898 460970 129134
rect 461206 128898 461248 129134
rect 460928 128866 461248 128898
rect 491648 129454 491968 129486
rect 491648 129218 491690 129454
rect 491926 129218 491968 129454
rect 491648 129134 491968 129218
rect 491648 128898 491690 129134
rect 491926 128898 491968 129134
rect 491648 128866 491968 128898
rect 522368 129454 522688 129486
rect 522368 129218 522410 129454
rect 522646 129218 522688 129454
rect 522368 129134 522688 129218
rect 522368 128898 522410 129134
rect 522646 128898 522688 129134
rect 522368 128866 522688 128898
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 46208 111454 46528 111486
rect 46208 111218 46250 111454
rect 46486 111218 46528 111454
rect 46208 111134 46528 111218
rect 46208 110898 46250 111134
rect 46486 110898 46528 111134
rect 46208 110866 46528 110898
rect 76928 111454 77248 111486
rect 76928 111218 76970 111454
rect 77206 111218 77248 111454
rect 76928 111134 77248 111218
rect 76928 110898 76970 111134
rect 77206 110898 77248 111134
rect 76928 110866 77248 110898
rect 107648 111454 107968 111486
rect 107648 111218 107690 111454
rect 107926 111218 107968 111454
rect 107648 111134 107968 111218
rect 107648 110898 107690 111134
rect 107926 110898 107968 111134
rect 107648 110866 107968 110898
rect 138368 111454 138688 111486
rect 138368 111218 138410 111454
rect 138646 111218 138688 111454
rect 138368 111134 138688 111218
rect 138368 110898 138410 111134
rect 138646 110898 138688 111134
rect 138368 110866 138688 110898
rect 169088 111454 169408 111486
rect 169088 111218 169130 111454
rect 169366 111218 169408 111454
rect 169088 111134 169408 111218
rect 169088 110898 169130 111134
rect 169366 110898 169408 111134
rect 169088 110866 169408 110898
rect 199808 111454 200128 111486
rect 199808 111218 199850 111454
rect 200086 111218 200128 111454
rect 199808 111134 200128 111218
rect 199808 110898 199850 111134
rect 200086 110898 200128 111134
rect 199808 110866 200128 110898
rect 230528 111454 230848 111486
rect 230528 111218 230570 111454
rect 230806 111218 230848 111454
rect 230528 111134 230848 111218
rect 230528 110898 230570 111134
rect 230806 110898 230848 111134
rect 230528 110866 230848 110898
rect 261248 111454 261568 111486
rect 261248 111218 261290 111454
rect 261526 111218 261568 111454
rect 261248 111134 261568 111218
rect 261248 110898 261290 111134
rect 261526 110898 261568 111134
rect 261248 110866 261568 110898
rect 291968 111454 292288 111486
rect 291968 111218 292010 111454
rect 292246 111218 292288 111454
rect 291968 111134 292288 111218
rect 291968 110898 292010 111134
rect 292246 110898 292288 111134
rect 291968 110866 292288 110898
rect 322688 111454 323008 111486
rect 322688 111218 322730 111454
rect 322966 111218 323008 111454
rect 322688 111134 323008 111218
rect 322688 110898 322730 111134
rect 322966 110898 323008 111134
rect 322688 110866 323008 110898
rect 353408 111454 353728 111486
rect 353408 111218 353450 111454
rect 353686 111218 353728 111454
rect 353408 111134 353728 111218
rect 353408 110898 353450 111134
rect 353686 110898 353728 111134
rect 353408 110866 353728 110898
rect 384128 111454 384448 111486
rect 384128 111218 384170 111454
rect 384406 111218 384448 111454
rect 384128 111134 384448 111218
rect 384128 110898 384170 111134
rect 384406 110898 384448 111134
rect 384128 110866 384448 110898
rect 414848 111454 415168 111486
rect 414848 111218 414890 111454
rect 415126 111218 415168 111454
rect 414848 111134 415168 111218
rect 414848 110898 414890 111134
rect 415126 110898 415168 111134
rect 414848 110866 415168 110898
rect 445568 111454 445888 111486
rect 445568 111218 445610 111454
rect 445846 111218 445888 111454
rect 445568 111134 445888 111218
rect 445568 110898 445610 111134
rect 445846 110898 445888 111134
rect 445568 110866 445888 110898
rect 476288 111454 476608 111486
rect 476288 111218 476330 111454
rect 476566 111218 476608 111454
rect 476288 111134 476608 111218
rect 476288 110898 476330 111134
rect 476566 110898 476608 111134
rect 476288 110866 476608 110898
rect 507008 111454 507328 111486
rect 507008 111218 507050 111454
rect 507286 111218 507328 111454
rect 507008 111134 507328 111218
rect 507008 110898 507050 111134
rect 507286 110898 507328 111134
rect 507008 110866 507328 110898
rect 537728 111454 538048 111486
rect 537728 111218 537770 111454
rect 538006 111218 538048 111454
rect 537728 111134 538048 111218
rect 537728 110898 537770 111134
rect 538006 110898 538048 111134
rect 537728 110866 538048 110898
rect 61568 93454 61888 93486
rect 61568 93218 61610 93454
rect 61846 93218 61888 93454
rect 61568 93134 61888 93218
rect 61568 92898 61610 93134
rect 61846 92898 61888 93134
rect 61568 92866 61888 92898
rect 92288 93454 92608 93486
rect 92288 93218 92330 93454
rect 92566 93218 92608 93454
rect 92288 93134 92608 93218
rect 92288 92898 92330 93134
rect 92566 92898 92608 93134
rect 92288 92866 92608 92898
rect 123008 93454 123328 93486
rect 123008 93218 123050 93454
rect 123286 93218 123328 93454
rect 123008 93134 123328 93218
rect 123008 92898 123050 93134
rect 123286 92898 123328 93134
rect 123008 92866 123328 92898
rect 153728 93454 154048 93486
rect 153728 93218 153770 93454
rect 154006 93218 154048 93454
rect 153728 93134 154048 93218
rect 153728 92898 153770 93134
rect 154006 92898 154048 93134
rect 153728 92866 154048 92898
rect 184448 93454 184768 93486
rect 184448 93218 184490 93454
rect 184726 93218 184768 93454
rect 184448 93134 184768 93218
rect 184448 92898 184490 93134
rect 184726 92898 184768 93134
rect 184448 92866 184768 92898
rect 215168 93454 215488 93486
rect 215168 93218 215210 93454
rect 215446 93218 215488 93454
rect 215168 93134 215488 93218
rect 215168 92898 215210 93134
rect 215446 92898 215488 93134
rect 215168 92866 215488 92898
rect 245888 93454 246208 93486
rect 245888 93218 245930 93454
rect 246166 93218 246208 93454
rect 245888 93134 246208 93218
rect 245888 92898 245930 93134
rect 246166 92898 246208 93134
rect 245888 92866 246208 92898
rect 276608 93454 276928 93486
rect 276608 93218 276650 93454
rect 276886 93218 276928 93454
rect 276608 93134 276928 93218
rect 276608 92898 276650 93134
rect 276886 92898 276928 93134
rect 276608 92866 276928 92898
rect 307328 93454 307648 93486
rect 307328 93218 307370 93454
rect 307606 93218 307648 93454
rect 307328 93134 307648 93218
rect 307328 92898 307370 93134
rect 307606 92898 307648 93134
rect 307328 92866 307648 92898
rect 338048 93454 338368 93486
rect 338048 93218 338090 93454
rect 338326 93218 338368 93454
rect 338048 93134 338368 93218
rect 338048 92898 338090 93134
rect 338326 92898 338368 93134
rect 338048 92866 338368 92898
rect 368768 93454 369088 93486
rect 368768 93218 368810 93454
rect 369046 93218 369088 93454
rect 368768 93134 369088 93218
rect 368768 92898 368810 93134
rect 369046 92898 369088 93134
rect 368768 92866 369088 92898
rect 399488 93454 399808 93486
rect 399488 93218 399530 93454
rect 399766 93218 399808 93454
rect 399488 93134 399808 93218
rect 399488 92898 399530 93134
rect 399766 92898 399808 93134
rect 399488 92866 399808 92898
rect 430208 93454 430528 93486
rect 430208 93218 430250 93454
rect 430486 93218 430528 93454
rect 430208 93134 430528 93218
rect 430208 92898 430250 93134
rect 430486 92898 430528 93134
rect 430208 92866 430528 92898
rect 460928 93454 461248 93486
rect 460928 93218 460970 93454
rect 461206 93218 461248 93454
rect 460928 93134 461248 93218
rect 460928 92898 460970 93134
rect 461206 92898 461248 93134
rect 460928 92866 461248 92898
rect 491648 93454 491968 93486
rect 491648 93218 491690 93454
rect 491926 93218 491968 93454
rect 491648 93134 491968 93218
rect 491648 92898 491690 93134
rect 491926 92898 491968 93134
rect 491648 92866 491968 92898
rect 522368 93454 522688 93486
rect 522368 93218 522410 93454
rect 522646 93218 522688 93454
rect 522368 93134 522688 93218
rect 522368 92898 522410 93134
rect 522646 92898 522688 93134
rect 522368 92866 522688 92898
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 46208 75454 46528 75486
rect 46208 75218 46250 75454
rect 46486 75218 46528 75454
rect 46208 75134 46528 75218
rect 46208 74898 46250 75134
rect 46486 74898 46528 75134
rect 46208 74866 46528 74898
rect 76928 75454 77248 75486
rect 76928 75218 76970 75454
rect 77206 75218 77248 75454
rect 76928 75134 77248 75218
rect 76928 74898 76970 75134
rect 77206 74898 77248 75134
rect 76928 74866 77248 74898
rect 107648 75454 107968 75486
rect 107648 75218 107690 75454
rect 107926 75218 107968 75454
rect 107648 75134 107968 75218
rect 107648 74898 107690 75134
rect 107926 74898 107968 75134
rect 107648 74866 107968 74898
rect 138368 75454 138688 75486
rect 138368 75218 138410 75454
rect 138646 75218 138688 75454
rect 138368 75134 138688 75218
rect 138368 74898 138410 75134
rect 138646 74898 138688 75134
rect 138368 74866 138688 74898
rect 169088 75454 169408 75486
rect 169088 75218 169130 75454
rect 169366 75218 169408 75454
rect 169088 75134 169408 75218
rect 169088 74898 169130 75134
rect 169366 74898 169408 75134
rect 169088 74866 169408 74898
rect 199808 75454 200128 75486
rect 199808 75218 199850 75454
rect 200086 75218 200128 75454
rect 199808 75134 200128 75218
rect 199808 74898 199850 75134
rect 200086 74898 200128 75134
rect 199808 74866 200128 74898
rect 230528 75454 230848 75486
rect 230528 75218 230570 75454
rect 230806 75218 230848 75454
rect 230528 75134 230848 75218
rect 230528 74898 230570 75134
rect 230806 74898 230848 75134
rect 230528 74866 230848 74898
rect 261248 75454 261568 75486
rect 261248 75218 261290 75454
rect 261526 75218 261568 75454
rect 261248 75134 261568 75218
rect 261248 74898 261290 75134
rect 261526 74898 261568 75134
rect 261248 74866 261568 74898
rect 291968 75454 292288 75486
rect 291968 75218 292010 75454
rect 292246 75218 292288 75454
rect 291968 75134 292288 75218
rect 291968 74898 292010 75134
rect 292246 74898 292288 75134
rect 291968 74866 292288 74898
rect 322688 75454 323008 75486
rect 322688 75218 322730 75454
rect 322966 75218 323008 75454
rect 322688 75134 323008 75218
rect 322688 74898 322730 75134
rect 322966 74898 323008 75134
rect 322688 74866 323008 74898
rect 353408 75454 353728 75486
rect 353408 75218 353450 75454
rect 353686 75218 353728 75454
rect 353408 75134 353728 75218
rect 353408 74898 353450 75134
rect 353686 74898 353728 75134
rect 353408 74866 353728 74898
rect 384128 75454 384448 75486
rect 384128 75218 384170 75454
rect 384406 75218 384448 75454
rect 384128 75134 384448 75218
rect 384128 74898 384170 75134
rect 384406 74898 384448 75134
rect 384128 74866 384448 74898
rect 414848 75454 415168 75486
rect 414848 75218 414890 75454
rect 415126 75218 415168 75454
rect 414848 75134 415168 75218
rect 414848 74898 414890 75134
rect 415126 74898 415168 75134
rect 414848 74866 415168 74898
rect 445568 75454 445888 75486
rect 445568 75218 445610 75454
rect 445846 75218 445888 75454
rect 445568 75134 445888 75218
rect 445568 74898 445610 75134
rect 445846 74898 445888 75134
rect 445568 74866 445888 74898
rect 476288 75454 476608 75486
rect 476288 75218 476330 75454
rect 476566 75218 476608 75454
rect 476288 75134 476608 75218
rect 476288 74898 476330 75134
rect 476566 74898 476608 75134
rect 476288 74866 476608 74898
rect 507008 75454 507328 75486
rect 507008 75218 507050 75454
rect 507286 75218 507328 75454
rect 507008 75134 507328 75218
rect 507008 74898 507050 75134
rect 507286 74898 507328 75134
rect 507008 74866 507328 74898
rect 537728 75454 538048 75486
rect 537728 75218 537770 75454
rect 538006 75218 538048 75454
rect 537728 75134 538048 75218
rect 537728 74898 537770 75134
rect 538006 74898 538048 75134
rect 537728 74866 538048 74898
rect 61568 57454 61888 57486
rect 61568 57218 61610 57454
rect 61846 57218 61888 57454
rect 61568 57134 61888 57218
rect 61568 56898 61610 57134
rect 61846 56898 61888 57134
rect 61568 56866 61888 56898
rect 92288 57454 92608 57486
rect 92288 57218 92330 57454
rect 92566 57218 92608 57454
rect 92288 57134 92608 57218
rect 92288 56898 92330 57134
rect 92566 56898 92608 57134
rect 92288 56866 92608 56898
rect 123008 57454 123328 57486
rect 123008 57218 123050 57454
rect 123286 57218 123328 57454
rect 123008 57134 123328 57218
rect 123008 56898 123050 57134
rect 123286 56898 123328 57134
rect 123008 56866 123328 56898
rect 153728 57454 154048 57486
rect 153728 57218 153770 57454
rect 154006 57218 154048 57454
rect 153728 57134 154048 57218
rect 153728 56898 153770 57134
rect 154006 56898 154048 57134
rect 153728 56866 154048 56898
rect 184448 57454 184768 57486
rect 184448 57218 184490 57454
rect 184726 57218 184768 57454
rect 184448 57134 184768 57218
rect 184448 56898 184490 57134
rect 184726 56898 184768 57134
rect 184448 56866 184768 56898
rect 215168 57454 215488 57486
rect 215168 57218 215210 57454
rect 215446 57218 215488 57454
rect 215168 57134 215488 57218
rect 215168 56898 215210 57134
rect 215446 56898 215488 57134
rect 215168 56866 215488 56898
rect 245888 57454 246208 57486
rect 245888 57218 245930 57454
rect 246166 57218 246208 57454
rect 245888 57134 246208 57218
rect 245888 56898 245930 57134
rect 246166 56898 246208 57134
rect 245888 56866 246208 56898
rect 276608 57454 276928 57486
rect 276608 57218 276650 57454
rect 276886 57218 276928 57454
rect 276608 57134 276928 57218
rect 276608 56898 276650 57134
rect 276886 56898 276928 57134
rect 276608 56866 276928 56898
rect 307328 57454 307648 57486
rect 307328 57218 307370 57454
rect 307606 57218 307648 57454
rect 307328 57134 307648 57218
rect 307328 56898 307370 57134
rect 307606 56898 307648 57134
rect 307328 56866 307648 56898
rect 338048 57454 338368 57486
rect 338048 57218 338090 57454
rect 338326 57218 338368 57454
rect 338048 57134 338368 57218
rect 338048 56898 338090 57134
rect 338326 56898 338368 57134
rect 338048 56866 338368 56898
rect 368768 57454 369088 57486
rect 368768 57218 368810 57454
rect 369046 57218 369088 57454
rect 368768 57134 369088 57218
rect 368768 56898 368810 57134
rect 369046 56898 369088 57134
rect 368768 56866 369088 56898
rect 399488 57454 399808 57486
rect 399488 57218 399530 57454
rect 399766 57218 399808 57454
rect 399488 57134 399808 57218
rect 399488 56898 399530 57134
rect 399766 56898 399808 57134
rect 399488 56866 399808 56898
rect 430208 57454 430528 57486
rect 430208 57218 430250 57454
rect 430486 57218 430528 57454
rect 430208 57134 430528 57218
rect 430208 56898 430250 57134
rect 430486 56898 430528 57134
rect 430208 56866 430528 56898
rect 460928 57454 461248 57486
rect 460928 57218 460970 57454
rect 461206 57218 461248 57454
rect 460928 57134 461248 57218
rect 460928 56898 460970 57134
rect 461206 56898 461248 57134
rect 460928 56866 461248 56898
rect 491648 57454 491968 57486
rect 491648 57218 491690 57454
rect 491926 57218 491968 57454
rect 491648 57134 491968 57218
rect 491648 56898 491690 57134
rect 491926 56898 491968 57134
rect 491648 56866 491968 56898
rect 522368 57454 522688 57486
rect 522368 57218 522410 57454
rect 522646 57218 522688 57454
rect 522368 57134 522688 57218
rect 522368 56898 522410 57134
rect 522646 56898 522688 57134
rect 522368 56866 522688 56898
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 7174 42134 40000
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 10894 45854 40000
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 40000
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 40000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 40000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 40000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 40000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 40000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 40000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 40000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 40000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 40000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 40000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 40000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 40000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 40000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 40000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 40000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 40000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 40000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 40000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 40000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 40000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 40000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 7174 150134 40000
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 40000
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 40000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 40000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 40000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 40000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 40000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 40000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 40000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 40000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 40000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 40000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 40000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 40000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 40000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 40000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 40000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 40000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 40000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 40000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 40000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 40000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 40000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 40000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 40000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 40000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 40000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 40000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 40000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 40000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 40000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 40000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 40000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 40000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 40000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 40000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 40000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 40000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 40000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 40000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 40000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 40000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 40000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 40000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 40000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 40000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 40000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 40000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 40000
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 40000
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 40000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 40000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 40000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 40000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 40000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 40000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 40000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 40000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 40000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 40000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 40000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 40000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 40000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 40000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 40000
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 40000
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 40000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 40000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 40000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 40000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 40000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 40000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 7174 474134 40000
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 10894 477854 40000
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 40000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 40000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 40000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 40000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 40000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 40000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 7174 510134 40000
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 10894 513854 40000
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 40000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 40000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 40000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 28894 531854 40000
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 32614 535574 40000
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 39454 542414 40000
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 7174 546134 40000
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 46250 543218 46486 543454
rect 46250 542898 46486 543134
rect 76970 543218 77206 543454
rect 76970 542898 77206 543134
rect 107690 543218 107926 543454
rect 107690 542898 107926 543134
rect 138410 543218 138646 543454
rect 138410 542898 138646 543134
rect 169130 543218 169366 543454
rect 169130 542898 169366 543134
rect 199850 543218 200086 543454
rect 199850 542898 200086 543134
rect 230570 543218 230806 543454
rect 230570 542898 230806 543134
rect 261290 543218 261526 543454
rect 261290 542898 261526 543134
rect 292010 543218 292246 543454
rect 292010 542898 292246 543134
rect 322730 543218 322966 543454
rect 322730 542898 322966 543134
rect 353450 543218 353686 543454
rect 353450 542898 353686 543134
rect 384170 543218 384406 543454
rect 384170 542898 384406 543134
rect 414890 543218 415126 543454
rect 414890 542898 415126 543134
rect 445610 543218 445846 543454
rect 445610 542898 445846 543134
rect 476330 543218 476566 543454
rect 476330 542898 476566 543134
rect 507050 543218 507286 543454
rect 507050 542898 507286 543134
rect 537770 543218 538006 543454
rect 537770 542898 538006 543134
rect 61610 525218 61846 525454
rect 61610 524898 61846 525134
rect 92330 525218 92566 525454
rect 92330 524898 92566 525134
rect 123050 525218 123286 525454
rect 123050 524898 123286 525134
rect 153770 525218 154006 525454
rect 153770 524898 154006 525134
rect 184490 525218 184726 525454
rect 184490 524898 184726 525134
rect 215210 525218 215446 525454
rect 215210 524898 215446 525134
rect 245930 525218 246166 525454
rect 245930 524898 246166 525134
rect 276650 525218 276886 525454
rect 276650 524898 276886 525134
rect 307370 525218 307606 525454
rect 307370 524898 307606 525134
rect 338090 525218 338326 525454
rect 338090 524898 338326 525134
rect 368810 525218 369046 525454
rect 368810 524898 369046 525134
rect 399530 525218 399766 525454
rect 399530 524898 399766 525134
rect 430250 525218 430486 525454
rect 430250 524898 430486 525134
rect 460970 525218 461206 525454
rect 460970 524898 461206 525134
rect 491690 525218 491926 525454
rect 491690 524898 491926 525134
rect 522410 525218 522646 525454
rect 522410 524898 522646 525134
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 46250 507218 46486 507454
rect 46250 506898 46486 507134
rect 76970 507218 77206 507454
rect 76970 506898 77206 507134
rect 107690 507218 107926 507454
rect 107690 506898 107926 507134
rect 138410 507218 138646 507454
rect 138410 506898 138646 507134
rect 169130 507218 169366 507454
rect 169130 506898 169366 507134
rect 199850 507218 200086 507454
rect 199850 506898 200086 507134
rect 230570 507218 230806 507454
rect 230570 506898 230806 507134
rect 261290 507218 261526 507454
rect 261290 506898 261526 507134
rect 292010 507218 292246 507454
rect 292010 506898 292246 507134
rect 322730 507218 322966 507454
rect 322730 506898 322966 507134
rect 353450 507218 353686 507454
rect 353450 506898 353686 507134
rect 384170 507218 384406 507454
rect 384170 506898 384406 507134
rect 414890 507218 415126 507454
rect 414890 506898 415126 507134
rect 445610 507218 445846 507454
rect 445610 506898 445846 507134
rect 476330 507218 476566 507454
rect 476330 506898 476566 507134
rect 507050 507218 507286 507454
rect 507050 506898 507286 507134
rect 537770 507218 538006 507454
rect 537770 506898 538006 507134
rect 61610 489218 61846 489454
rect 61610 488898 61846 489134
rect 92330 489218 92566 489454
rect 92330 488898 92566 489134
rect 123050 489218 123286 489454
rect 123050 488898 123286 489134
rect 153770 489218 154006 489454
rect 153770 488898 154006 489134
rect 184490 489218 184726 489454
rect 184490 488898 184726 489134
rect 215210 489218 215446 489454
rect 215210 488898 215446 489134
rect 245930 489218 246166 489454
rect 245930 488898 246166 489134
rect 276650 489218 276886 489454
rect 276650 488898 276886 489134
rect 307370 489218 307606 489454
rect 307370 488898 307606 489134
rect 338090 489218 338326 489454
rect 338090 488898 338326 489134
rect 368810 489218 369046 489454
rect 368810 488898 369046 489134
rect 399530 489218 399766 489454
rect 399530 488898 399766 489134
rect 430250 489218 430486 489454
rect 430250 488898 430486 489134
rect 460970 489218 461206 489454
rect 460970 488898 461206 489134
rect 491690 489218 491926 489454
rect 491690 488898 491926 489134
rect 522410 489218 522646 489454
rect 522410 488898 522646 489134
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 46250 471218 46486 471454
rect 46250 470898 46486 471134
rect 76970 471218 77206 471454
rect 76970 470898 77206 471134
rect 107690 471218 107926 471454
rect 107690 470898 107926 471134
rect 138410 471218 138646 471454
rect 138410 470898 138646 471134
rect 169130 471218 169366 471454
rect 169130 470898 169366 471134
rect 199850 471218 200086 471454
rect 199850 470898 200086 471134
rect 230570 471218 230806 471454
rect 230570 470898 230806 471134
rect 261290 471218 261526 471454
rect 261290 470898 261526 471134
rect 292010 471218 292246 471454
rect 292010 470898 292246 471134
rect 322730 471218 322966 471454
rect 322730 470898 322966 471134
rect 353450 471218 353686 471454
rect 353450 470898 353686 471134
rect 384170 471218 384406 471454
rect 384170 470898 384406 471134
rect 414890 471218 415126 471454
rect 414890 470898 415126 471134
rect 445610 471218 445846 471454
rect 445610 470898 445846 471134
rect 476330 471218 476566 471454
rect 476330 470898 476566 471134
rect 507050 471218 507286 471454
rect 507050 470898 507286 471134
rect 537770 471218 538006 471454
rect 537770 470898 538006 471134
rect 61610 453218 61846 453454
rect 61610 452898 61846 453134
rect 92330 453218 92566 453454
rect 92330 452898 92566 453134
rect 123050 453218 123286 453454
rect 123050 452898 123286 453134
rect 153770 453218 154006 453454
rect 153770 452898 154006 453134
rect 184490 453218 184726 453454
rect 184490 452898 184726 453134
rect 215210 453218 215446 453454
rect 215210 452898 215446 453134
rect 245930 453218 246166 453454
rect 245930 452898 246166 453134
rect 276650 453218 276886 453454
rect 276650 452898 276886 453134
rect 307370 453218 307606 453454
rect 307370 452898 307606 453134
rect 338090 453218 338326 453454
rect 338090 452898 338326 453134
rect 368810 453218 369046 453454
rect 368810 452898 369046 453134
rect 399530 453218 399766 453454
rect 399530 452898 399766 453134
rect 430250 453218 430486 453454
rect 430250 452898 430486 453134
rect 460970 453218 461206 453454
rect 460970 452898 461206 453134
rect 491690 453218 491926 453454
rect 491690 452898 491926 453134
rect 522410 453218 522646 453454
rect 522410 452898 522646 453134
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 46250 435218 46486 435454
rect 46250 434898 46486 435134
rect 76970 435218 77206 435454
rect 76970 434898 77206 435134
rect 107690 435218 107926 435454
rect 107690 434898 107926 435134
rect 138410 435218 138646 435454
rect 138410 434898 138646 435134
rect 169130 435218 169366 435454
rect 169130 434898 169366 435134
rect 199850 435218 200086 435454
rect 199850 434898 200086 435134
rect 230570 435218 230806 435454
rect 230570 434898 230806 435134
rect 261290 435218 261526 435454
rect 261290 434898 261526 435134
rect 292010 435218 292246 435454
rect 292010 434898 292246 435134
rect 322730 435218 322966 435454
rect 322730 434898 322966 435134
rect 353450 435218 353686 435454
rect 353450 434898 353686 435134
rect 384170 435218 384406 435454
rect 384170 434898 384406 435134
rect 414890 435218 415126 435454
rect 414890 434898 415126 435134
rect 445610 435218 445846 435454
rect 445610 434898 445846 435134
rect 476330 435218 476566 435454
rect 476330 434898 476566 435134
rect 507050 435218 507286 435454
rect 507050 434898 507286 435134
rect 537770 435218 538006 435454
rect 537770 434898 538006 435134
rect 61610 417218 61846 417454
rect 61610 416898 61846 417134
rect 92330 417218 92566 417454
rect 92330 416898 92566 417134
rect 123050 417218 123286 417454
rect 123050 416898 123286 417134
rect 153770 417218 154006 417454
rect 153770 416898 154006 417134
rect 184490 417218 184726 417454
rect 184490 416898 184726 417134
rect 215210 417218 215446 417454
rect 215210 416898 215446 417134
rect 245930 417218 246166 417454
rect 245930 416898 246166 417134
rect 276650 417218 276886 417454
rect 276650 416898 276886 417134
rect 307370 417218 307606 417454
rect 307370 416898 307606 417134
rect 338090 417218 338326 417454
rect 338090 416898 338326 417134
rect 368810 417218 369046 417454
rect 368810 416898 369046 417134
rect 399530 417218 399766 417454
rect 399530 416898 399766 417134
rect 430250 417218 430486 417454
rect 430250 416898 430486 417134
rect 460970 417218 461206 417454
rect 460970 416898 461206 417134
rect 491690 417218 491926 417454
rect 491690 416898 491926 417134
rect 522410 417218 522646 417454
rect 522410 416898 522646 417134
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 46250 399218 46486 399454
rect 46250 398898 46486 399134
rect 76970 399218 77206 399454
rect 76970 398898 77206 399134
rect 107690 399218 107926 399454
rect 107690 398898 107926 399134
rect 138410 399218 138646 399454
rect 138410 398898 138646 399134
rect 169130 399218 169366 399454
rect 169130 398898 169366 399134
rect 199850 399218 200086 399454
rect 199850 398898 200086 399134
rect 230570 399218 230806 399454
rect 230570 398898 230806 399134
rect 261290 399218 261526 399454
rect 261290 398898 261526 399134
rect 292010 399218 292246 399454
rect 292010 398898 292246 399134
rect 322730 399218 322966 399454
rect 322730 398898 322966 399134
rect 353450 399218 353686 399454
rect 353450 398898 353686 399134
rect 384170 399218 384406 399454
rect 384170 398898 384406 399134
rect 414890 399218 415126 399454
rect 414890 398898 415126 399134
rect 445610 399218 445846 399454
rect 445610 398898 445846 399134
rect 476330 399218 476566 399454
rect 476330 398898 476566 399134
rect 507050 399218 507286 399454
rect 507050 398898 507286 399134
rect 537770 399218 538006 399454
rect 537770 398898 538006 399134
rect 61610 381218 61846 381454
rect 61610 380898 61846 381134
rect 92330 381218 92566 381454
rect 92330 380898 92566 381134
rect 123050 381218 123286 381454
rect 123050 380898 123286 381134
rect 153770 381218 154006 381454
rect 153770 380898 154006 381134
rect 184490 381218 184726 381454
rect 184490 380898 184726 381134
rect 215210 381218 215446 381454
rect 215210 380898 215446 381134
rect 245930 381218 246166 381454
rect 245930 380898 246166 381134
rect 276650 381218 276886 381454
rect 276650 380898 276886 381134
rect 307370 381218 307606 381454
rect 307370 380898 307606 381134
rect 338090 381218 338326 381454
rect 338090 380898 338326 381134
rect 368810 381218 369046 381454
rect 368810 380898 369046 381134
rect 399530 381218 399766 381454
rect 399530 380898 399766 381134
rect 430250 381218 430486 381454
rect 430250 380898 430486 381134
rect 460970 381218 461206 381454
rect 460970 380898 461206 381134
rect 491690 381218 491926 381454
rect 491690 380898 491926 381134
rect 522410 381218 522646 381454
rect 522410 380898 522646 381134
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 46250 363218 46486 363454
rect 46250 362898 46486 363134
rect 76970 363218 77206 363454
rect 76970 362898 77206 363134
rect 107690 363218 107926 363454
rect 107690 362898 107926 363134
rect 138410 363218 138646 363454
rect 138410 362898 138646 363134
rect 169130 363218 169366 363454
rect 169130 362898 169366 363134
rect 199850 363218 200086 363454
rect 199850 362898 200086 363134
rect 230570 363218 230806 363454
rect 230570 362898 230806 363134
rect 261290 363218 261526 363454
rect 261290 362898 261526 363134
rect 292010 363218 292246 363454
rect 292010 362898 292246 363134
rect 322730 363218 322966 363454
rect 322730 362898 322966 363134
rect 353450 363218 353686 363454
rect 353450 362898 353686 363134
rect 384170 363218 384406 363454
rect 384170 362898 384406 363134
rect 414890 363218 415126 363454
rect 414890 362898 415126 363134
rect 445610 363218 445846 363454
rect 445610 362898 445846 363134
rect 476330 363218 476566 363454
rect 476330 362898 476566 363134
rect 507050 363218 507286 363454
rect 507050 362898 507286 363134
rect 537770 363218 538006 363454
rect 537770 362898 538006 363134
rect 61610 345218 61846 345454
rect 61610 344898 61846 345134
rect 92330 345218 92566 345454
rect 92330 344898 92566 345134
rect 123050 345218 123286 345454
rect 123050 344898 123286 345134
rect 153770 345218 154006 345454
rect 153770 344898 154006 345134
rect 184490 345218 184726 345454
rect 184490 344898 184726 345134
rect 215210 345218 215446 345454
rect 215210 344898 215446 345134
rect 245930 345218 246166 345454
rect 245930 344898 246166 345134
rect 276650 345218 276886 345454
rect 276650 344898 276886 345134
rect 307370 345218 307606 345454
rect 307370 344898 307606 345134
rect 338090 345218 338326 345454
rect 338090 344898 338326 345134
rect 368810 345218 369046 345454
rect 368810 344898 369046 345134
rect 399530 345218 399766 345454
rect 399530 344898 399766 345134
rect 430250 345218 430486 345454
rect 430250 344898 430486 345134
rect 460970 345218 461206 345454
rect 460970 344898 461206 345134
rect 491690 345218 491926 345454
rect 491690 344898 491926 345134
rect 522410 345218 522646 345454
rect 522410 344898 522646 345134
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 46250 327218 46486 327454
rect 46250 326898 46486 327134
rect 76970 327218 77206 327454
rect 76970 326898 77206 327134
rect 107690 327218 107926 327454
rect 107690 326898 107926 327134
rect 138410 327218 138646 327454
rect 138410 326898 138646 327134
rect 169130 327218 169366 327454
rect 169130 326898 169366 327134
rect 199850 327218 200086 327454
rect 199850 326898 200086 327134
rect 230570 327218 230806 327454
rect 230570 326898 230806 327134
rect 261290 327218 261526 327454
rect 261290 326898 261526 327134
rect 292010 327218 292246 327454
rect 292010 326898 292246 327134
rect 322730 327218 322966 327454
rect 322730 326898 322966 327134
rect 353450 327218 353686 327454
rect 353450 326898 353686 327134
rect 384170 327218 384406 327454
rect 384170 326898 384406 327134
rect 414890 327218 415126 327454
rect 414890 326898 415126 327134
rect 445610 327218 445846 327454
rect 445610 326898 445846 327134
rect 476330 327218 476566 327454
rect 476330 326898 476566 327134
rect 507050 327218 507286 327454
rect 507050 326898 507286 327134
rect 537770 327218 538006 327454
rect 537770 326898 538006 327134
rect 61610 309218 61846 309454
rect 61610 308898 61846 309134
rect 92330 309218 92566 309454
rect 92330 308898 92566 309134
rect 123050 309218 123286 309454
rect 123050 308898 123286 309134
rect 153770 309218 154006 309454
rect 153770 308898 154006 309134
rect 184490 309218 184726 309454
rect 184490 308898 184726 309134
rect 215210 309218 215446 309454
rect 215210 308898 215446 309134
rect 245930 309218 246166 309454
rect 245930 308898 246166 309134
rect 276650 309218 276886 309454
rect 276650 308898 276886 309134
rect 307370 309218 307606 309454
rect 307370 308898 307606 309134
rect 338090 309218 338326 309454
rect 338090 308898 338326 309134
rect 368810 309218 369046 309454
rect 368810 308898 369046 309134
rect 399530 309218 399766 309454
rect 399530 308898 399766 309134
rect 430250 309218 430486 309454
rect 430250 308898 430486 309134
rect 460970 309218 461206 309454
rect 460970 308898 461206 309134
rect 491690 309218 491926 309454
rect 491690 308898 491926 309134
rect 522410 309218 522646 309454
rect 522410 308898 522646 309134
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 46250 291218 46486 291454
rect 46250 290898 46486 291134
rect 76970 291218 77206 291454
rect 76970 290898 77206 291134
rect 107690 291218 107926 291454
rect 107690 290898 107926 291134
rect 138410 291218 138646 291454
rect 138410 290898 138646 291134
rect 169130 291218 169366 291454
rect 169130 290898 169366 291134
rect 199850 291218 200086 291454
rect 199850 290898 200086 291134
rect 230570 291218 230806 291454
rect 230570 290898 230806 291134
rect 261290 291218 261526 291454
rect 261290 290898 261526 291134
rect 292010 291218 292246 291454
rect 292010 290898 292246 291134
rect 322730 291218 322966 291454
rect 322730 290898 322966 291134
rect 353450 291218 353686 291454
rect 353450 290898 353686 291134
rect 384170 291218 384406 291454
rect 384170 290898 384406 291134
rect 414890 291218 415126 291454
rect 414890 290898 415126 291134
rect 445610 291218 445846 291454
rect 445610 290898 445846 291134
rect 476330 291218 476566 291454
rect 476330 290898 476566 291134
rect 507050 291218 507286 291454
rect 507050 290898 507286 291134
rect 537770 291218 538006 291454
rect 537770 290898 538006 291134
rect 61610 273218 61846 273454
rect 61610 272898 61846 273134
rect 92330 273218 92566 273454
rect 92330 272898 92566 273134
rect 123050 273218 123286 273454
rect 123050 272898 123286 273134
rect 153770 273218 154006 273454
rect 153770 272898 154006 273134
rect 184490 273218 184726 273454
rect 184490 272898 184726 273134
rect 215210 273218 215446 273454
rect 215210 272898 215446 273134
rect 245930 273218 246166 273454
rect 245930 272898 246166 273134
rect 276650 273218 276886 273454
rect 276650 272898 276886 273134
rect 307370 273218 307606 273454
rect 307370 272898 307606 273134
rect 338090 273218 338326 273454
rect 338090 272898 338326 273134
rect 368810 273218 369046 273454
rect 368810 272898 369046 273134
rect 399530 273218 399766 273454
rect 399530 272898 399766 273134
rect 430250 273218 430486 273454
rect 430250 272898 430486 273134
rect 460970 273218 461206 273454
rect 460970 272898 461206 273134
rect 491690 273218 491926 273454
rect 491690 272898 491926 273134
rect 522410 273218 522646 273454
rect 522410 272898 522646 273134
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 46250 255218 46486 255454
rect 46250 254898 46486 255134
rect 76970 255218 77206 255454
rect 76970 254898 77206 255134
rect 107690 255218 107926 255454
rect 107690 254898 107926 255134
rect 138410 255218 138646 255454
rect 138410 254898 138646 255134
rect 169130 255218 169366 255454
rect 169130 254898 169366 255134
rect 199850 255218 200086 255454
rect 199850 254898 200086 255134
rect 230570 255218 230806 255454
rect 230570 254898 230806 255134
rect 261290 255218 261526 255454
rect 261290 254898 261526 255134
rect 292010 255218 292246 255454
rect 292010 254898 292246 255134
rect 322730 255218 322966 255454
rect 322730 254898 322966 255134
rect 353450 255218 353686 255454
rect 353450 254898 353686 255134
rect 384170 255218 384406 255454
rect 384170 254898 384406 255134
rect 414890 255218 415126 255454
rect 414890 254898 415126 255134
rect 445610 255218 445846 255454
rect 445610 254898 445846 255134
rect 476330 255218 476566 255454
rect 476330 254898 476566 255134
rect 507050 255218 507286 255454
rect 507050 254898 507286 255134
rect 537770 255218 538006 255454
rect 537770 254898 538006 255134
rect 61610 237218 61846 237454
rect 61610 236898 61846 237134
rect 92330 237218 92566 237454
rect 92330 236898 92566 237134
rect 123050 237218 123286 237454
rect 123050 236898 123286 237134
rect 153770 237218 154006 237454
rect 153770 236898 154006 237134
rect 184490 237218 184726 237454
rect 184490 236898 184726 237134
rect 215210 237218 215446 237454
rect 215210 236898 215446 237134
rect 245930 237218 246166 237454
rect 245930 236898 246166 237134
rect 276650 237218 276886 237454
rect 276650 236898 276886 237134
rect 307370 237218 307606 237454
rect 307370 236898 307606 237134
rect 338090 237218 338326 237454
rect 338090 236898 338326 237134
rect 368810 237218 369046 237454
rect 368810 236898 369046 237134
rect 399530 237218 399766 237454
rect 399530 236898 399766 237134
rect 430250 237218 430486 237454
rect 430250 236898 430486 237134
rect 460970 237218 461206 237454
rect 460970 236898 461206 237134
rect 491690 237218 491926 237454
rect 491690 236898 491926 237134
rect 522410 237218 522646 237454
rect 522410 236898 522646 237134
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 46250 219218 46486 219454
rect 46250 218898 46486 219134
rect 76970 219218 77206 219454
rect 76970 218898 77206 219134
rect 107690 219218 107926 219454
rect 107690 218898 107926 219134
rect 138410 219218 138646 219454
rect 138410 218898 138646 219134
rect 169130 219218 169366 219454
rect 169130 218898 169366 219134
rect 199850 219218 200086 219454
rect 199850 218898 200086 219134
rect 230570 219218 230806 219454
rect 230570 218898 230806 219134
rect 261290 219218 261526 219454
rect 261290 218898 261526 219134
rect 292010 219218 292246 219454
rect 292010 218898 292246 219134
rect 322730 219218 322966 219454
rect 322730 218898 322966 219134
rect 353450 219218 353686 219454
rect 353450 218898 353686 219134
rect 384170 219218 384406 219454
rect 384170 218898 384406 219134
rect 414890 219218 415126 219454
rect 414890 218898 415126 219134
rect 445610 219218 445846 219454
rect 445610 218898 445846 219134
rect 476330 219218 476566 219454
rect 476330 218898 476566 219134
rect 507050 219218 507286 219454
rect 507050 218898 507286 219134
rect 537770 219218 538006 219454
rect 537770 218898 538006 219134
rect 61610 201218 61846 201454
rect 61610 200898 61846 201134
rect 92330 201218 92566 201454
rect 92330 200898 92566 201134
rect 123050 201218 123286 201454
rect 123050 200898 123286 201134
rect 153770 201218 154006 201454
rect 153770 200898 154006 201134
rect 184490 201218 184726 201454
rect 184490 200898 184726 201134
rect 215210 201218 215446 201454
rect 215210 200898 215446 201134
rect 245930 201218 246166 201454
rect 245930 200898 246166 201134
rect 276650 201218 276886 201454
rect 276650 200898 276886 201134
rect 307370 201218 307606 201454
rect 307370 200898 307606 201134
rect 338090 201218 338326 201454
rect 338090 200898 338326 201134
rect 368810 201218 369046 201454
rect 368810 200898 369046 201134
rect 399530 201218 399766 201454
rect 399530 200898 399766 201134
rect 430250 201218 430486 201454
rect 430250 200898 430486 201134
rect 460970 201218 461206 201454
rect 460970 200898 461206 201134
rect 491690 201218 491926 201454
rect 491690 200898 491926 201134
rect 522410 201218 522646 201454
rect 522410 200898 522646 201134
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 46250 183218 46486 183454
rect 46250 182898 46486 183134
rect 76970 183218 77206 183454
rect 76970 182898 77206 183134
rect 107690 183218 107926 183454
rect 107690 182898 107926 183134
rect 138410 183218 138646 183454
rect 138410 182898 138646 183134
rect 169130 183218 169366 183454
rect 169130 182898 169366 183134
rect 199850 183218 200086 183454
rect 199850 182898 200086 183134
rect 230570 183218 230806 183454
rect 230570 182898 230806 183134
rect 261290 183218 261526 183454
rect 261290 182898 261526 183134
rect 292010 183218 292246 183454
rect 292010 182898 292246 183134
rect 322730 183218 322966 183454
rect 322730 182898 322966 183134
rect 353450 183218 353686 183454
rect 353450 182898 353686 183134
rect 384170 183218 384406 183454
rect 384170 182898 384406 183134
rect 414890 183218 415126 183454
rect 414890 182898 415126 183134
rect 445610 183218 445846 183454
rect 445610 182898 445846 183134
rect 476330 183218 476566 183454
rect 476330 182898 476566 183134
rect 507050 183218 507286 183454
rect 507050 182898 507286 183134
rect 537770 183218 538006 183454
rect 537770 182898 538006 183134
rect 61610 165218 61846 165454
rect 61610 164898 61846 165134
rect 92330 165218 92566 165454
rect 92330 164898 92566 165134
rect 123050 165218 123286 165454
rect 123050 164898 123286 165134
rect 153770 165218 154006 165454
rect 153770 164898 154006 165134
rect 184490 165218 184726 165454
rect 184490 164898 184726 165134
rect 215210 165218 215446 165454
rect 215210 164898 215446 165134
rect 245930 165218 246166 165454
rect 245930 164898 246166 165134
rect 276650 165218 276886 165454
rect 276650 164898 276886 165134
rect 307370 165218 307606 165454
rect 307370 164898 307606 165134
rect 338090 165218 338326 165454
rect 338090 164898 338326 165134
rect 368810 165218 369046 165454
rect 368810 164898 369046 165134
rect 399530 165218 399766 165454
rect 399530 164898 399766 165134
rect 430250 165218 430486 165454
rect 430250 164898 430486 165134
rect 460970 165218 461206 165454
rect 460970 164898 461206 165134
rect 491690 165218 491926 165454
rect 491690 164898 491926 165134
rect 522410 165218 522646 165454
rect 522410 164898 522646 165134
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 46250 147218 46486 147454
rect 46250 146898 46486 147134
rect 76970 147218 77206 147454
rect 76970 146898 77206 147134
rect 107690 147218 107926 147454
rect 107690 146898 107926 147134
rect 138410 147218 138646 147454
rect 138410 146898 138646 147134
rect 169130 147218 169366 147454
rect 169130 146898 169366 147134
rect 199850 147218 200086 147454
rect 199850 146898 200086 147134
rect 230570 147218 230806 147454
rect 230570 146898 230806 147134
rect 261290 147218 261526 147454
rect 261290 146898 261526 147134
rect 292010 147218 292246 147454
rect 292010 146898 292246 147134
rect 322730 147218 322966 147454
rect 322730 146898 322966 147134
rect 353450 147218 353686 147454
rect 353450 146898 353686 147134
rect 384170 147218 384406 147454
rect 384170 146898 384406 147134
rect 414890 147218 415126 147454
rect 414890 146898 415126 147134
rect 445610 147218 445846 147454
rect 445610 146898 445846 147134
rect 476330 147218 476566 147454
rect 476330 146898 476566 147134
rect 507050 147218 507286 147454
rect 507050 146898 507286 147134
rect 537770 147218 538006 147454
rect 537770 146898 538006 147134
rect 61610 129218 61846 129454
rect 61610 128898 61846 129134
rect 92330 129218 92566 129454
rect 92330 128898 92566 129134
rect 123050 129218 123286 129454
rect 123050 128898 123286 129134
rect 153770 129218 154006 129454
rect 153770 128898 154006 129134
rect 184490 129218 184726 129454
rect 184490 128898 184726 129134
rect 215210 129218 215446 129454
rect 215210 128898 215446 129134
rect 245930 129218 246166 129454
rect 245930 128898 246166 129134
rect 276650 129218 276886 129454
rect 276650 128898 276886 129134
rect 307370 129218 307606 129454
rect 307370 128898 307606 129134
rect 338090 129218 338326 129454
rect 338090 128898 338326 129134
rect 368810 129218 369046 129454
rect 368810 128898 369046 129134
rect 399530 129218 399766 129454
rect 399530 128898 399766 129134
rect 430250 129218 430486 129454
rect 430250 128898 430486 129134
rect 460970 129218 461206 129454
rect 460970 128898 461206 129134
rect 491690 129218 491926 129454
rect 491690 128898 491926 129134
rect 522410 129218 522646 129454
rect 522410 128898 522646 129134
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 46250 111218 46486 111454
rect 46250 110898 46486 111134
rect 76970 111218 77206 111454
rect 76970 110898 77206 111134
rect 107690 111218 107926 111454
rect 107690 110898 107926 111134
rect 138410 111218 138646 111454
rect 138410 110898 138646 111134
rect 169130 111218 169366 111454
rect 169130 110898 169366 111134
rect 199850 111218 200086 111454
rect 199850 110898 200086 111134
rect 230570 111218 230806 111454
rect 230570 110898 230806 111134
rect 261290 111218 261526 111454
rect 261290 110898 261526 111134
rect 292010 111218 292246 111454
rect 292010 110898 292246 111134
rect 322730 111218 322966 111454
rect 322730 110898 322966 111134
rect 353450 111218 353686 111454
rect 353450 110898 353686 111134
rect 384170 111218 384406 111454
rect 384170 110898 384406 111134
rect 414890 111218 415126 111454
rect 414890 110898 415126 111134
rect 445610 111218 445846 111454
rect 445610 110898 445846 111134
rect 476330 111218 476566 111454
rect 476330 110898 476566 111134
rect 507050 111218 507286 111454
rect 507050 110898 507286 111134
rect 537770 111218 538006 111454
rect 537770 110898 538006 111134
rect 61610 93218 61846 93454
rect 61610 92898 61846 93134
rect 92330 93218 92566 93454
rect 92330 92898 92566 93134
rect 123050 93218 123286 93454
rect 123050 92898 123286 93134
rect 153770 93218 154006 93454
rect 153770 92898 154006 93134
rect 184490 93218 184726 93454
rect 184490 92898 184726 93134
rect 215210 93218 215446 93454
rect 215210 92898 215446 93134
rect 245930 93218 246166 93454
rect 245930 92898 246166 93134
rect 276650 93218 276886 93454
rect 276650 92898 276886 93134
rect 307370 93218 307606 93454
rect 307370 92898 307606 93134
rect 338090 93218 338326 93454
rect 338090 92898 338326 93134
rect 368810 93218 369046 93454
rect 368810 92898 369046 93134
rect 399530 93218 399766 93454
rect 399530 92898 399766 93134
rect 430250 93218 430486 93454
rect 430250 92898 430486 93134
rect 460970 93218 461206 93454
rect 460970 92898 461206 93134
rect 491690 93218 491926 93454
rect 491690 92898 491926 93134
rect 522410 93218 522646 93454
rect 522410 92898 522646 93134
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 46250 75218 46486 75454
rect 46250 74898 46486 75134
rect 76970 75218 77206 75454
rect 76970 74898 77206 75134
rect 107690 75218 107926 75454
rect 107690 74898 107926 75134
rect 138410 75218 138646 75454
rect 138410 74898 138646 75134
rect 169130 75218 169366 75454
rect 169130 74898 169366 75134
rect 199850 75218 200086 75454
rect 199850 74898 200086 75134
rect 230570 75218 230806 75454
rect 230570 74898 230806 75134
rect 261290 75218 261526 75454
rect 261290 74898 261526 75134
rect 292010 75218 292246 75454
rect 292010 74898 292246 75134
rect 322730 75218 322966 75454
rect 322730 74898 322966 75134
rect 353450 75218 353686 75454
rect 353450 74898 353686 75134
rect 384170 75218 384406 75454
rect 384170 74898 384406 75134
rect 414890 75218 415126 75454
rect 414890 74898 415126 75134
rect 445610 75218 445846 75454
rect 445610 74898 445846 75134
rect 476330 75218 476566 75454
rect 476330 74898 476566 75134
rect 507050 75218 507286 75454
rect 507050 74898 507286 75134
rect 537770 75218 538006 75454
rect 537770 74898 538006 75134
rect 61610 57218 61846 57454
rect 61610 56898 61846 57134
rect 92330 57218 92566 57454
rect 92330 56898 92566 57134
rect 123050 57218 123286 57454
rect 123050 56898 123286 57134
rect 153770 57218 154006 57454
rect 153770 56898 154006 57134
rect 184490 57218 184726 57454
rect 184490 56898 184726 57134
rect 215210 57218 215446 57454
rect 215210 56898 215446 57134
rect 245930 57218 246166 57454
rect 245930 56898 246166 57134
rect 276650 57218 276886 57454
rect 276650 56898 276886 57134
rect 307370 57218 307606 57454
rect 307370 56898 307606 57134
rect 338090 57218 338326 57454
rect 338090 56898 338326 57134
rect 368810 57218 369046 57454
rect 368810 56898 369046 57134
rect 399530 57218 399766 57454
rect 399530 56898 399766 57134
rect 430250 57218 430486 57454
rect 430250 56898 430486 57134
rect 460970 57218 461206 57454
rect 460970 56898 461206 57134
rect 491690 57218 491926 57454
rect 491690 56898 491926 57134
rect 522410 57218 522646 57454
rect 522410 56898 522646 57134
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 46250 543454
rect 46486 543218 76970 543454
rect 77206 543218 107690 543454
rect 107926 543218 138410 543454
rect 138646 543218 169130 543454
rect 169366 543218 199850 543454
rect 200086 543218 230570 543454
rect 230806 543218 261290 543454
rect 261526 543218 292010 543454
rect 292246 543218 322730 543454
rect 322966 543218 353450 543454
rect 353686 543218 384170 543454
rect 384406 543218 414890 543454
rect 415126 543218 445610 543454
rect 445846 543218 476330 543454
rect 476566 543218 507050 543454
rect 507286 543218 537770 543454
rect 538006 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 46250 543134
rect 46486 542898 76970 543134
rect 77206 542898 107690 543134
rect 107926 542898 138410 543134
rect 138646 542898 169130 543134
rect 169366 542898 199850 543134
rect 200086 542898 230570 543134
rect 230806 542898 261290 543134
rect 261526 542898 292010 543134
rect 292246 542898 322730 543134
rect 322966 542898 353450 543134
rect 353686 542898 384170 543134
rect 384406 542898 414890 543134
rect 415126 542898 445610 543134
rect 445846 542898 476330 543134
rect 476566 542898 507050 543134
rect 507286 542898 537770 543134
rect 538006 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 61610 525454
rect 61846 525218 92330 525454
rect 92566 525218 123050 525454
rect 123286 525218 153770 525454
rect 154006 525218 184490 525454
rect 184726 525218 215210 525454
rect 215446 525218 245930 525454
rect 246166 525218 276650 525454
rect 276886 525218 307370 525454
rect 307606 525218 338090 525454
rect 338326 525218 368810 525454
rect 369046 525218 399530 525454
rect 399766 525218 430250 525454
rect 430486 525218 460970 525454
rect 461206 525218 491690 525454
rect 491926 525218 522410 525454
rect 522646 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 61610 525134
rect 61846 524898 92330 525134
rect 92566 524898 123050 525134
rect 123286 524898 153770 525134
rect 154006 524898 184490 525134
rect 184726 524898 215210 525134
rect 215446 524898 245930 525134
rect 246166 524898 276650 525134
rect 276886 524898 307370 525134
rect 307606 524898 338090 525134
rect 338326 524898 368810 525134
rect 369046 524898 399530 525134
rect 399766 524898 430250 525134
rect 430486 524898 460970 525134
rect 461206 524898 491690 525134
rect 491926 524898 522410 525134
rect 522646 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 46250 507454
rect 46486 507218 76970 507454
rect 77206 507218 107690 507454
rect 107926 507218 138410 507454
rect 138646 507218 169130 507454
rect 169366 507218 199850 507454
rect 200086 507218 230570 507454
rect 230806 507218 261290 507454
rect 261526 507218 292010 507454
rect 292246 507218 322730 507454
rect 322966 507218 353450 507454
rect 353686 507218 384170 507454
rect 384406 507218 414890 507454
rect 415126 507218 445610 507454
rect 445846 507218 476330 507454
rect 476566 507218 507050 507454
rect 507286 507218 537770 507454
rect 538006 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 46250 507134
rect 46486 506898 76970 507134
rect 77206 506898 107690 507134
rect 107926 506898 138410 507134
rect 138646 506898 169130 507134
rect 169366 506898 199850 507134
rect 200086 506898 230570 507134
rect 230806 506898 261290 507134
rect 261526 506898 292010 507134
rect 292246 506898 322730 507134
rect 322966 506898 353450 507134
rect 353686 506898 384170 507134
rect 384406 506898 414890 507134
rect 415126 506898 445610 507134
rect 445846 506898 476330 507134
rect 476566 506898 507050 507134
rect 507286 506898 537770 507134
rect 538006 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 61610 489454
rect 61846 489218 92330 489454
rect 92566 489218 123050 489454
rect 123286 489218 153770 489454
rect 154006 489218 184490 489454
rect 184726 489218 215210 489454
rect 215446 489218 245930 489454
rect 246166 489218 276650 489454
rect 276886 489218 307370 489454
rect 307606 489218 338090 489454
rect 338326 489218 368810 489454
rect 369046 489218 399530 489454
rect 399766 489218 430250 489454
rect 430486 489218 460970 489454
rect 461206 489218 491690 489454
rect 491926 489218 522410 489454
rect 522646 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 61610 489134
rect 61846 488898 92330 489134
rect 92566 488898 123050 489134
rect 123286 488898 153770 489134
rect 154006 488898 184490 489134
rect 184726 488898 215210 489134
rect 215446 488898 245930 489134
rect 246166 488898 276650 489134
rect 276886 488898 307370 489134
rect 307606 488898 338090 489134
rect 338326 488898 368810 489134
rect 369046 488898 399530 489134
rect 399766 488898 430250 489134
rect 430486 488898 460970 489134
rect 461206 488898 491690 489134
rect 491926 488898 522410 489134
rect 522646 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 46250 471454
rect 46486 471218 76970 471454
rect 77206 471218 107690 471454
rect 107926 471218 138410 471454
rect 138646 471218 169130 471454
rect 169366 471218 199850 471454
rect 200086 471218 230570 471454
rect 230806 471218 261290 471454
rect 261526 471218 292010 471454
rect 292246 471218 322730 471454
rect 322966 471218 353450 471454
rect 353686 471218 384170 471454
rect 384406 471218 414890 471454
rect 415126 471218 445610 471454
rect 445846 471218 476330 471454
rect 476566 471218 507050 471454
rect 507286 471218 537770 471454
rect 538006 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 46250 471134
rect 46486 470898 76970 471134
rect 77206 470898 107690 471134
rect 107926 470898 138410 471134
rect 138646 470898 169130 471134
rect 169366 470898 199850 471134
rect 200086 470898 230570 471134
rect 230806 470898 261290 471134
rect 261526 470898 292010 471134
rect 292246 470898 322730 471134
rect 322966 470898 353450 471134
rect 353686 470898 384170 471134
rect 384406 470898 414890 471134
rect 415126 470898 445610 471134
rect 445846 470898 476330 471134
rect 476566 470898 507050 471134
rect 507286 470898 537770 471134
rect 538006 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 61610 453454
rect 61846 453218 92330 453454
rect 92566 453218 123050 453454
rect 123286 453218 153770 453454
rect 154006 453218 184490 453454
rect 184726 453218 215210 453454
rect 215446 453218 245930 453454
rect 246166 453218 276650 453454
rect 276886 453218 307370 453454
rect 307606 453218 338090 453454
rect 338326 453218 368810 453454
rect 369046 453218 399530 453454
rect 399766 453218 430250 453454
rect 430486 453218 460970 453454
rect 461206 453218 491690 453454
rect 491926 453218 522410 453454
rect 522646 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 61610 453134
rect 61846 452898 92330 453134
rect 92566 452898 123050 453134
rect 123286 452898 153770 453134
rect 154006 452898 184490 453134
rect 184726 452898 215210 453134
rect 215446 452898 245930 453134
rect 246166 452898 276650 453134
rect 276886 452898 307370 453134
rect 307606 452898 338090 453134
rect 338326 452898 368810 453134
rect 369046 452898 399530 453134
rect 399766 452898 430250 453134
rect 430486 452898 460970 453134
rect 461206 452898 491690 453134
rect 491926 452898 522410 453134
rect 522646 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 46250 435454
rect 46486 435218 76970 435454
rect 77206 435218 107690 435454
rect 107926 435218 138410 435454
rect 138646 435218 169130 435454
rect 169366 435218 199850 435454
rect 200086 435218 230570 435454
rect 230806 435218 261290 435454
rect 261526 435218 292010 435454
rect 292246 435218 322730 435454
rect 322966 435218 353450 435454
rect 353686 435218 384170 435454
rect 384406 435218 414890 435454
rect 415126 435218 445610 435454
rect 445846 435218 476330 435454
rect 476566 435218 507050 435454
rect 507286 435218 537770 435454
rect 538006 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 46250 435134
rect 46486 434898 76970 435134
rect 77206 434898 107690 435134
rect 107926 434898 138410 435134
rect 138646 434898 169130 435134
rect 169366 434898 199850 435134
rect 200086 434898 230570 435134
rect 230806 434898 261290 435134
rect 261526 434898 292010 435134
rect 292246 434898 322730 435134
rect 322966 434898 353450 435134
rect 353686 434898 384170 435134
rect 384406 434898 414890 435134
rect 415126 434898 445610 435134
rect 445846 434898 476330 435134
rect 476566 434898 507050 435134
rect 507286 434898 537770 435134
rect 538006 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 61610 417454
rect 61846 417218 92330 417454
rect 92566 417218 123050 417454
rect 123286 417218 153770 417454
rect 154006 417218 184490 417454
rect 184726 417218 215210 417454
rect 215446 417218 245930 417454
rect 246166 417218 276650 417454
rect 276886 417218 307370 417454
rect 307606 417218 338090 417454
rect 338326 417218 368810 417454
rect 369046 417218 399530 417454
rect 399766 417218 430250 417454
rect 430486 417218 460970 417454
rect 461206 417218 491690 417454
rect 491926 417218 522410 417454
rect 522646 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 61610 417134
rect 61846 416898 92330 417134
rect 92566 416898 123050 417134
rect 123286 416898 153770 417134
rect 154006 416898 184490 417134
rect 184726 416898 215210 417134
rect 215446 416898 245930 417134
rect 246166 416898 276650 417134
rect 276886 416898 307370 417134
rect 307606 416898 338090 417134
rect 338326 416898 368810 417134
rect 369046 416898 399530 417134
rect 399766 416898 430250 417134
rect 430486 416898 460970 417134
rect 461206 416898 491690 417134
rect 491926 416898 522410 417134
rect 522646 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 46250 399454
rect 46486 399218 76970 399454
rect 77206 399218 107690 399454
rect 107926 399218 138410 399454
rect 138646 399218 169130 399454
rect 169366 399218 199850 399454
rect 200086 399218 230570 399454
rect 230806 399218 261290 399454
rect 261526 399218 292010 399454
rect 292246 399218 322730 399454
rect 322966 399218 353450 399454
rect 353686 399218 384170 399454
rect 384406 399218 414890 399454
rect 415126 399218 445610 399454
rect 445846 399218 476330 399454
rect 476566 399218 507050 399454
rect 507286 399218 537770 399454
rect 538006 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 46250 399134
rect 46486 398898 76970 399134
rect 77206 398898 107690 399134
rect 107926 398898 138410 399134
rect 138646 398898 169130 399134
rect 169366 398898 199850 399134
rect 200086 398898 230570 399134
rect 230806 398898 261290 399134
rect 261526 398898 292010 399134
rect 292246 398898 322730 399134
rect 322966 398898 353450 399134
rect 353686 398898 384170 399134
rect 384406 398898 414890 399134
rect 415126 398898 445610 399134
rect 445846 398898 476330 399134
rect 476566 398898 507050 399134
rect 507286 398898 537770 399134
rect 538006 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 61610 381454
rect 61846 381218 92330 381454
rect 92566 381218 123050 381454
rect 123286 381218 153770 381454
rect 154006 381218 184490 381454
rect 184726 381218 215210 381454
rect 215446 381218 245930 381454
rect 246166 381218 276650 381454
rect 276886 381218 307370 381454
rect 307606 381218 338090 381454
rect 338326 381218 368810 381454
rect 369046 381218 399530 381454
rect 399766 381218 430250 381454
rect 430486 381218 460970 381454
rect 461206 381218 491690 381454
rect 491926 381218 522410 381454
rect 522646 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 61610 381134
rect 61846 380898 92330 381134
rect 92566 380898 123050 381134
rect 123286 380898 153770 381134
rect 154006 380898 184490 381134
rect 184726 380898 215210 381134
rect 215446 380898 245930 381134
rect 246166 380898 276650 381134
rect 276886 380898 307370 381134
rect 307606 380898 338090 381134
rect 338326 380898 368810 381134
rect 369046 380898 399530 381134
rect 399766 380898 430250 381134
rect 430486 380898 460970 381134
rect 461206 380898 491690 381134
rect 491926 380898 522410 381134
rect 522646 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 46250 363454
rect 46486 363218 76970 363454
rect 77206 363218 107690 363454
rect 107926 363218 138410 363454
rect 138646 363218 169130 363454
rect 169366 363218 199850 363454
rect 200086 363218 230570 363454
rect 230806 363218 261290 363454
rect 261526 363218 292010 363454
rect 292246 363218 322730 363454
rect 322966 363218 353450 363454
rect 353686 363218 384170 363454
rect 384406 363218 414890 363454
rect 415126 363218 445610 363454
rect 445846 363218 476330 363454
rect 476566 363218 507050 363454
rect 507286 363218 537770 363454
rect 538006 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 46250 363134
rect 46486 362898 76970 363134
rect 77206 362898 107690 363134
rect 107926 362898 138410 363134
rect 138646 362898 169130 363134
rect 169366 362898 199850 363134
rect 200086 362898 230570 363134
rect 230806 362898 261290 363134
rect 261526 362898 292010 363134
rect 292246 362898 322730 363134
rect 322966 362898 353450 363134
rect 353686 362898 384170 363134
rect 384406 362898 414890 363134
rect 415126 362898 445610 363134
rect 445846 362898 476330 363134
rect 476566 362898 507050 363134
rect 507286 362898 537770 363134
rect 538006 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 61610 345454
rect 61846 345218 92330 345454
rect 92566 345218 123050 345454
rect 123286 345218 153770 345454
rect 154006 345218 184490 345454
rect 184726 345218 215210 345454
rect 215446 345218 245930 345454
rect 246166 345218 276650 345454
rect 276886 345218 307370 345454
rect 307606 345218 338090 345454
rect 338326 345218 368810 345454
rect 369046 345218 399530 345454
rect 399766 345218 430250 345454
rect 430486 345218 460970 345454
rect 461206 345218 491690 345454
rect 491926 345218 522410 345454
rect 522646 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 61610 345134
rect 61846 344898 92330 345134
rect 92566 344898 123050 345134
rect 123286 344898 153770 345134
rect 154006 344898 184490 345134
rect 184726 344898 215210 345134
rect 215446 344898 245930 345134
rect 246166 344898 276650 345134
rect 276886 344898 307370 345134
rect 307606 344898 338090 345134
rect 338326 344898 368810 345134
rect 369046 344898 399530 345134
rect 399766 344898 430250 345134
rect 430486 344898 460970 345134
rect 461206 344898 491690 345134
rect 491926 344898 522410 345134
rect 522646 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 46250 327454
rect 46486 327218 76970 327454
rect 77206 327218 107690 327454
rect 107926 327218 138410 327454
rect 138646 327218 169130 327454
rect 169366 327218 199850 327454
rect 200086 327218 230570 327454
rect 230806 327218 261290 327454
rect 261526 327218 292010 327454
rect 292246 327218 322730 327454
rect 322966 327218 353450 327454
rect 353686 327218 384170 327454
rect 384406 327218 414890 327454
rect 415126 327218 445610 327454
rect 445846 327218 476330 327454
rect 476566 327218 507050 327454
rect 507286 327218 537770 327454
rect 538006 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 46250 327134
rect 46486 326898 76970 327134
rect 77206 326898 107690 327134
rect 107926 326898 138410 327134
rect 138646 326898 169130 327134
rect 169366 326898 199850 327134
rect 200086 326898 230570 327134
rect 230806 326898 261290 327134
rect 261526 326898 292010 327134
rect 292246 326898 322730 327134
rect 322966 326898 353450 327134
rect 353686 326898 384170 327134
rect 384406 326898 414890 327134
rect 415126 326898 445610 327134
rect 445846 326898 476330 327134
rect 476566 326898 507050 327134
rect 507286 326898 537770 327134
rect 538006 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 61610 309454
rect 61846 309218 92330 309454
rect 92566 309218 123050 309454
rect 123286 309218 153770 309454
rect 154006 309218 184490 309454
rect 184726 309218 215210 309454
rect 215446 309218 245930 309454
rect 246166 309218 276650 309454
rect 276886 309218 307370 309454
rect 307606 309218 338090 309454
rect 338326 309218 368810 309454
rect 369046 309218 399530 309454
rect 399766 309218 430250 309454
rect 430486 309218 460970 309454
rect 461206 309218 491690 309454
rect 491926 309218 522410 309454
rect 522646 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 61610 309134
rect 61846 308898 92330 309134
rect 92566 308898 123050 309134
rect 123286 308898 153770 309134
rect 154006 308898 184490 309134
rect 184726 308898 215210 309134
rect 215446 308898 245930 309134
rect 246166 308898 276650 309134
rect 276886 308898 307370 309134
rect 307606 308898 338090 309134
rect 338326 308898 368810 309134
rect 369046 308898 399530 309134
rect 399766 308898 430250 309134
rect 430486 308898 460970 309134
rect 461206 308898 491690 309134
rect 491926 308898 522410 309134
rect 522646 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 46250 291454
rect 46486 291218 76970 291454
rect 77206 291218 107690 291454
rect 107926 291218 138410 291454
rect 138646 291218 169130 291454
rect 169366 291218 199850 291454
rect 200086 291218 230570 291454
rect 230806 291218 261290 291454
rect 261526 291218 292010 291454
rect 292246 291218 322730 291454
rect 322966 291218 353450 291454
rect 353686 291218 384170 291454
rect 384406 291218 414890 291454
rect 415126 291218 445610 291454
rect 445846 291218 476330 291454
rect 476566 291218 507050 291454
rect 507286 291218 537770 291454
rect 538006 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 46250 291134
rect 46486 290898 76970 291134
rect 77206 290898 107690 291134
rect 107926 290898 138410 291134
rect 138646 290898 169130 291134
rect 169366 290898 199850 291134
rect 200086 290898 230570 291134
rect 230806 290898 261290 291134
rect 261526 290898 292010 291134
rect 292246 290898 322730 291134
rect 322966 290898 353450 291134
rect 353686 290898 384170 291134
rect 384406 290898 414890 291134
rect 415126 290898 445610 291134
rect 445846 290898 476330 291134
rect 476566 290898 507050 291134
rect 507286 290898 537770 291134
rect 538006 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 61610 273454
rect 61846 273218 92330 273454
rect 92566 273218 123050 273454
rect 123286 273218 153770 273454
rect 154006 273218 184490 273454
rect 184726 273218 215210 273454
rect 215446 273218 245930 273454
rect 246166 273218 276650 273454
rect 276886 273218 307370 273454
rect 307606 273218 338090 273454
rect 338326 273218 368810 273454
rect 369046 273218 399530 273454
rect 399766 273218 430250 273454
rect 430486 273218 460970 273454
rect 461206 273218 491690 273454
rect 491926 273218 522410 273454
rect 522646 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 61610 273134
rect 61846 272898 92330 273134
rect 92566 272898 123050 273134
rect 123286 272898 153770 273134
rect 154006 272898 184490 273134
rect 184726 272898 215210 273134
rect 215446 272898 245930 273134
rect 246166 272898 276650 273134
rect 276886 272898 307370 273134
rect 307606 272898 338090 273134
rect 338326 272898 368810 273134
rect 369046 272898 399530 273134
rect 399766 272898 430250 273134
rect 430486 272898 460970 273134
rect 461206 272898 491690 273134
rect 491926 272898 522410 273134
rect 522646 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 46250 255454
rect 46486 255218 76970 255454
rect 77206 255218 107690 255454
rect 107926 255218 138410 255454
rect 138646 255218 169130 255454
rect 169366 255218 199850 255454
rect 200086 255218 230570 255454
rect 230806 255218 261290 255454
rect 261526 255218 292010 255454
rect 292246 255218 322730 255454
rect 322966 255218 353450 255454
rect 353686 255218 384170 255454
rect 384406 255218 414890 255454
rect 415126 255218 445610 255454
rect 445846 255218 476330 255454
rect 476566 255218 507050 255454
rect 507286 255218 537770 255454
rect 538006 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 46250 255134
rect 46486 254898 76970 255134
rect 77206 254898 107690 255134
rect 107926 254898 138410 255134
rect 138646 254898 169130 255134
rect 169366 254898 199850 255134
rect 200086 254898 230570 255134
rect 230806 254898 261290 255134
rect 261526 254898 292010 255134
rect 292246 254898 322730 255134
rect 322966 254898 353450 255134
rect 353686 254898 384170 255134
rect 384406 254898 414890 255134
rect 415126 254898 445610 255134
rect 445846 254898 476330 255134
rect 476566 254898 507050 255134
rect 507286 254898 537770 255134
rect 538006 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 61610 237454
rect 61846 237218 92330 237454
rect 92566 237218 123050 237454
rect 123286 237218 153770 237454
rect 154006 237218 184490 237454
rect 184726 237218 215210 237454
rect 215446 237218 245930 237454
rect 246166 237218 276650 237454
rect 276886 237218 307370 237454
rect 307606 237218 338090 237454
rect 338326 237218 368810 237454
rect 369046 237218 399530 237454
rect 399766 237218 430250 237454
rect 430486 237218 460970 237454
rect 461206 237218 491690 237454
rect 491926 237218 522410 237454
rect 522646 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 61610 237134
rect 61846 236898 92330 237134
rect 92566 236898 123050 237134
rect 123286 236898 153770 237134
rect 154006 236898 184490 237134
rect 184726 236898 215210 237134
rect 215446 236898 245930 237134
rect 246166 236898 276650 237134
rect 276886 236898 307370 237134
rect 307606 236898 338090 237134
rect 338326 236898 368810 237134
rect 369046 236898 399530 237134
rect 399766 236898 430250 237134
rect 430486 236898 460970 237134
rect 461206 236898 491690 237134
rect 491926 236898 522410 237134
rect 522646 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 46250 219454
rect 46486 219218 76970 219454
rect 77206 219218 107690 219454
rect 107926 219218 138410 219454
rect 138646 219218 169130 219454
rect 169366 219218 199850 219454
rect 200086 219218 230570 219454
rect 230806 219218 261290 219454
rect 261526 219218 292010 219454
rect 292246 219218 322730 219454
rect 322966 219218 353450 219454
rect 353686 219218 384170 219454
rect 384406 219218 414890 219454
rect 415126 219218 445610 219454
rect 445846 219218 476330 219454
rect 476566 219218 507050 219454
rect 507286 219218 537770 219454
rect 538006 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 46250 219134
rect 46486 218898 76970 219134
rect 77206 218898 107690 219134
rect 107926 218898 138410 219134
rect 138646 218898 169130 219134
rect 169366 218898 199850 219134
rect 200086 218898 230570 219134
rect 230806 218898 261290 219134
rect 261526 218898 292010 219134
rect 292246 218898 322730 219134
rect 322966 218898 353450 219134
rect 353686 218898 384170 219134
rect 384406 218898 414890 219134
rect 415126 218898 445610 219134
rect 445846 218898 476330 219134
rect 476566 218898 507050 219134
rect 507286 218898 537770 219134
rect 538006 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 61610 201454
rect 61846 201218 92330 201454
rect 92566 201218 123050 201454
rect 123286 201218 153770 201454
rect 154006 201218 184490 201454
rect 184726 201218 215210 201454
rect 215446 201218 245930 201454
rect 246166 201218 276650 201454
rect 276886 201218 307370 201454
rect 307606 201218 338090 201454
rect 338326 201218 368810 201454
rect 369046 201218 399530 201454
rect 399766 201218 430250 201454
rect 430486 201218 460970 201454
rect 461206 201218 491690 201454
rect 491926 201218 522410 201454
rect 522646 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 61610 201134
rect 61846 200898 92330 201134
rect 92566 200898 123050 201134
rect 123286 200898 153770 201134
rect 154006 200898 184490 201134
rect 184726 200898 215210 201134
rect 215446 200898 245930 201134
rect 246166 200898 276650 201134
rect 276886 200898 307370 201134
rect 307606 200898 338090 201134
rect 338326 200898 368810 201134
rect 369046 200898 399530 201134
rect 399766 200898 430250 201134
rect 430486 200898 460970 201134
rect 461206 200898 491690 201134
rect 491926 200898 522410 201134
rect 522646 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 46250 183454
rect 46486 183218 76970 183454
rect 77206 183218 107690 183454
rect 107926 183218 138410 183454
rect 138646 183218 169130 183454
rect 169366 183218 199850 183454
rect 200086 183218 230570 183454
rect 230806 183218 261290 183454
rect 261526 183218 292010 183454
rect 292246 183218 322730 183454
rect 322966 183218 353450 183454
rect 353686 183218 384170 183454
rect 384406 183218 414890 183454
rect 415126 183218 445610 183454
rect 445846 183218 476330 183454
rect 476566 183218 507050 183454
rect 507286 183218 537770 183454
rect 538006 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 46250 183134
rect 46486 182898 76970 183134
rect 77206 182898 107690 183134
rect 107926 182898 138410 183134
rect 138646 182898 169130 183134
rect 169366 182898 199850 183134
rect 200086 182898 230570 183134
rect 230806 182898 261290 183134
rect 261526 182898 292010 183134
rect 292246 182898 322730 183134
rect 322966 182898 353450 183134
rect 353686 182898 384170 183134
rect 384406 182898 414890 183134
rect 415126 182898 445610 183134
rect 445846 182898 476330 183134
rect 476566 182898 507050 183134
rect 507286 182898 537770 183134
rect 538006 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 61610 165454
rect 61846 165218 92330 165454
rect 92566 165218 123050 165454
rect 123286 165218 153770 165454
rect 154006 165218 184490 165454
rect 184726 165218 215210 165454
rect 215446 165218 245930 165454
rect 246166 165218 276650 165454
rect 276886 165218 307370 165454
rect 307606 165218 338090 165454
rect 338326 165218 368810 165454
rect 369046 165218 399530 165454
rect 399766 165218 430250 165454
rect 430486 165218 460970 165454
rect 461206 165218 491690 165454
rect 491926 165218 522410 165454
rect 522646 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 61610 165134
rect 61846 164898 92330 165134
rect 92566 164898 123050 165134
rect 123286 164898 153770 165134
rect 154006 164898 184490 165134
rect 184726 164898 215210 165134
rect 215446 164898 245930 165134
rect 246166 164898 276650 165134
rect 276886 164898 307370 165134
rect 307606 164898 338090 165134
rect 338326 164898 368810 165134
rect 369046 164898 399530 165134
rect 399766 164898 430250 165134
rect 430486 164898 460970 165134
rect 461206 164898 491690 165134
rect 491926 164898 522410 165134
rect 522646 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 46250 147454
rect 46486 147218 76970 147454
rect 77206 147218 107690 147454
rect 107926 147218 138410 147454
rect 138646 147218 169130 147454
rect 169366 147218 199850 147454
rect 200086 147218 230570 147454
rect 230806 147218 261290 147454
rect 261526 147218 292010 147454
rect 292246 147218 322730 147454
rect 322966 147218 353450 147454
rect 353686 147218 384170 147454
rect 384406 147218 414890 147454
rect 415126 147218 445610 147454
rect 445846 147218 476330 147454
rect 476566 147218 507050 147454
rect 507286 147218 537770 147454
rect 538006 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 46250 147134
rect 46486 146898 76970 147134
rect 77206 146898 107690 147134
rect 107926 146898 138410 147134
rect 138646 146898 169130 147134
rect 169366 146898 199850 147134
rect 200086 146898 230570 147134
rect 230806 146898 261290 147134
rect 261526 146898 292010 147134
rect 292246 146898 322730 147134
rect 322966 146898 353450 147134
rect 353686 146898 384170 147134
rect 384406 146898 414890 147134
rect 415126 146898 445610 147134
rect 445846 146898 476330 147134
rect 476566 146898 507050 147134
rect 507286 146898 537770 147134
rect 538006 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 61610 129454
rect 61846 129218 92330 129454
rect 92566 129218 123050 129454
rect 123286 129218 153770 129454
rect 154006 129218 184490 129454
rect 184726 129218 215210 129454
rect 215446 129218 245930 129454
rect 246166 129218 276650 129454
rect 276886 129218 307370 129454
rect 307606 129218 338090 129454
rect 338326 129218 368810 129454
rect 369046 129218 399530 129454
rect 399766 129218 430250 129454
rect 430486 129218 460970 129454
rect 461206 129218 491690 129454
rect 491926 129218 522410 129454
rect 522646 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 61610 129134
rect 61846 128898 92330 129134
rect 92566 128898 123050 129134
rect 123286 128898 153770 129134
rect 154006 128898 184490 129134
rect 184726 128898 215210 129134
rect 215446 128898 245930 129134
rect 246166 128898 276650 129134
rect 276886 128898 307370 129134
rect 307606 128898 338090 129134
rect 338326 128898 368810 129134
rect 369046 128898 399530 129134
rect 399766 128898 430250 129134
rect 430486 128898 460970 129134
rect 461206 128898 491690 129134
rect 491926 128898 522410 129134
rect 522646 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 46250 111454
rect 46486 111218 76970 111454
rect 77206 111218 107690 111454
rect 107926 111218 138410 111454
rect 138646 111218 169130 111454
rect 169366 111218 199850 111454
rect 200086 111218 230570 111454
rect 230806 111218 261290 111454
rect 261526 111218 292010 111454
rect 292246 111218 322730 111454
rect 322966 111218 353450 111454
rect 353686 111218 384170 111454
rect 384406 111218 414890 111454
rect 415126 111218 445610 111454
rect 445846 111218 476330 111454
rect 476566 111218 507050 111454
rect 507286 111218 537770 111454
rect 538006 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 46250 111134
rect 46486 110898 76970 111134
rect 77206 110898 107690 111134
rect 107926 110898 138410 111134
rect 138646 110898 169130 111134
rect 169366 110898 199850 111134
rect 200086 110898 230570 111134
rect 230806 110898 261290 111134
rect 261526 110898 292010 111134
rect 292246 110898 322730 111134
rect 322966 110898 353450 111134
rect 353686 110898 384170 111134
rect 384406 110898 414890 111134
rect 415126 110898 445610 111134
rect 445846 110898 476330 111134
rect 476566 110898 507050 111134
rect 507286 110898 537770 111134
rect 538006 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 61610 93454
rect 61846 93218 92330 93454
rect 92566 93218 123050 93454
rect 123286 93218 153770 93454
rect 154006 93218 184490 93454
rect 184726 93218 215210 93454
rect 215446 93218 245930 93454
rect 246166 93218 276650 93454
rect 276886 93218 307370 93454
rect 307606 93218 338090 93454
rect 338326 93218 368810 93454
rect 369046 93218 399530 93454
rect 399766 93218 430250 93454
rect 430486 93218 460970 93454
rect 461206 93218 491690 93454
rect 491926 93218 522410 93454
rect 522646 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 61610 93134
rect 61846 92898 92330 93134
rect 92566 92898 123050 93134
rect 123286 92898 153770 93134
rect 154006 92898 184490 93134
rect 184726 92898 215210 93134
rect 215446 92898 245930 93134
rect 246166 92898 276650 93134
rect 276886 92898 307370 93134
rect 307606 92898 338090 93134
rect 338326 92898 368810 93134
rect 369046 92898 399530 93134
rect 399766 92898 430250 93134
rect 430486 92898 460970 93134
rect 461206 92898 491690 93134
rect 491926 92898 522410 93134
rect 522646 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 46250 75454
rect 46486 75218 76970 75454
rect 77206 75218 107690 75454
rect 107926 75218 138410 75454
rect 138646 75218 169130 75454
rect 169366 75218 199850 75454
rect 200086 75218 230570 75454
rect 230806 75218 261290 75454
rect 261526 75218 292010 75454
rect 292246 75218 322730 75454
rect 322966 75218 353450 75454
rect 353686 75218 384170 75454
rect 384406 75218 414890 75454
rect 415126 75218 445610 75454
rect 445846 75218 476330 75454
rect 476566 75218 507050 75454
rect 507286 75218 537770 75454
rect 538006 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 46250 75134
rect 46486 74898 76970 75134
rect 77206 74898 107690 75134
rect 107926 74898 138410 75134
rect 138646 74898 169130 75134
rect 169366 74898 199850 75134
rect 200086 74898 230570 75134
rect 230806 74898 261290 75134
rect 261526 74898 292010 75134
rect 292246 74898 322730 75134
rect 322966 74898 353450 75134
rect 353686 74898 384170 75134
rect 384406 74898 414890 75134
rect 415126 74898 445610 75134
rect 445846 74898 476330 75134
rect 476566 74898 507050 75134
rect 507286 74898 537770 75134
rect 538006 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 61610 57454
rect 61846 57218 92330 57454
rect 92566 57218 123050 57454
rect 123286 57218 153770 57454
rect 154006 57218 184490 57454
rect 184726 57218 215210 57454
rect 215446 57218 245930 57454
rect 246166 57218 276650 57454
rect 276886 57218 307370 57454
rect 307606 57218 338090 57454
rect 338326 57218 368810 57454
rect 369046 57218 399530 57454
rect 399766 57218 430250 57454
rect 430486 57218 460970 57454
rect 461206 57218 491690 57454
rect 491926 57218 522410 57454
rect 522646 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 61610 57134
rect 61846 56898 92330 57134
rect 92566 56898 123050 57134
rect 123286 56898 153770 57134
rect 154006 56898 184490 57134
rect 184726 56898 215210 57134
rect 215446 56898 245930 57134
rect 246166 56898 276650 57134
rect 276886 56898 307370 57134
rect 307606 56898 338090 57134
rect 338326 56898 368810 57134
rect 369046 56898 399530 57134
rect 399766 56898 430250 57134
rect 430486 56898 460970 57134
rect 461206 56898 491690 57134
rect 491926 56898 522410 57134
rect 522646 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1636060364
transform 1 0 42000 0 1 42000
box 474 0 501386 504086
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 548086 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 548086 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 548086 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 548086 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 548086 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 548086 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 548086 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 548086 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 548086 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 548086 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 548086 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 548086 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 548086 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 548086 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 548086 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 548086 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 548086 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 548086 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 548086 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 548086 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 548086 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 548086 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 548086 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 548086 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 548086 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 548086 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 548086 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 548086 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 548086 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 548086 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 548086 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 548086 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 548086 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 548086 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 548086 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 548086 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 548086 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 548086 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 548086 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 548086 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 548086 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 548086 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 548086 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 548086 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 548086 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 548086 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 548086 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 548086 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 548086 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 548086 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 548086 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 548086 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 548086 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 548086 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 548086 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 548086 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 548086 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 548086 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 548086 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 548086 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 548086 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 548086 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 548086 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 548086 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 548086 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 548086 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 548086 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 548086 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 548086 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 548086 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 548086 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 548086 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 548086 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 548086 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 548086 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 548086 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 548086 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 548086 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 548086 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 548086 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 548086 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 548086 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 548086 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 548086 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 548086 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 548086 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 548086 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 548086 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 548086 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 548086 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 548086 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 548086 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 548086 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 548086 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 548086 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 548086 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 548086 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 548086 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 548086 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 548086 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 548086 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 548086 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 548086 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 548086 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 548086 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 548086 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 548086 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 548086 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 548086 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 548086 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 548086 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 548086 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 548086 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
