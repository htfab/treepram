magic
tech sky130A
magscale 1 2
timestamp 1636029682
<< obsli1 >>
rect 1104 85 500756 501585
<< obsm1 >>
rect 474 8 501386 501616
<< metal2 >>
rect 2134 503286 2190 504086
rect 6458 503286 6514 504086
rect 10874 503286 10930 504086
rect 15290 503286 15346 504086
rect 19706 503286 19762 504086
rect 24122 503286 24178 504086
rect 28538 503286 28594 504086
rect 32954 503286 33010 504086
rect 37278 503286 37334 504086
rect 41694 503286 41750 504086
rect 46110 503286 46166 504086
rect 50526 503286 50582 504086
rect 54942 503286 54998 504086
rect 59358 503286 59414 504086
rect 63774 503286 63830 504086
rect 68098 503286 68154 504086
rect 72514 503286 72570 504086
rect 76930 503286 76986 504086
rect 81346 503286 81402 504086
rect 85762 503286 85818 504086
rect 90178 503286 90234 504086
rect 94594 503286 94650 504086
rect 98918 503286 98974 504086
rect 103334 503286 103390 504086
rect 107750 503286 107806 504086
rect 112166 503286 112222 504086
rect 116582 503286 116638 504086
rect 120998 503286 121054 504086
rect 125414 503286 125470 504086
rect 129738 503286 129794 504086
rect 134154 503286 134210 504086
rect 138570 503286 138626 504086
rect 142986 503286 143042 504086
rect 147402 503286 147458 504086
rect 151818 503286 151874 504086
rect 156234 503286 156290 504086
rect 160558 503286 160614 504086
rect 164974 503286 165030 504086
rect 169390 503286 169446 504086
rect 173806 503286 173862 504086
rect 178222 503286 178278 504086
rect 182638 503286 182694 504086
rect 187054 503286 187110 504086
rect 191378 503286 191434 504086
rect 195794 503286 195850 504086
rect 200210 503286 200266 504086
rect 204626 503286 204682 504086
rect 209042 503286 209098 504086
rect 213458 503286 213514 504086
rect 217874 503286 217930 504086
rect 222198 503286 222254 504086
rect 226614 503286 226670 504086
rect 231030 503286 231086 504086
rect 235446 503286 235502 504086
rect 239862 503286 239918 504086
rect 244278 503286 244334 504086
rect 248694 503286 248750 504086
rect 253110 503286 253166 504086
rect 257434 503286 257490 504086
rect 261850 503286 261906 504086
rect 266266 503286 266322 504086
rect 270682 503286 270738 504086
rect 275098 503286 275154 504086
rect 279514 503286 279570 504086
rect 283930 503286 283986 504086
rect 288254 503286 288310 504086
rect 292670 503286 292726 504086
rect 297086 503286 297142 504086
rect 301502 503286 301558 504086
rect 305918 503286 305974 504086
rect 310334 503286 310390 504086
rect 314750 503286 314806 504086
rect 319074 503286 319130 504086
rect 323490 503286 323546 504086
rect 327906 503286 327962 504086
rect 332322 503286 332378 504086
rect 336738 503286 336794 504086
rect 341154 503286 341210 504086
rect 345570 503286 345626 504086
rect 349894 503286 349950 504086
rect 354310 503286 354366 504086
rect 358726 503286 358782 504086
rect 363142 503286 363198 504086
rect 367558 503286 367614 504086
rect 371974 503286 372030 504086
rect 376390 503286 376446 504086
rect 380714 503286 380770 504086
rect 385130 503286 385186 504086
rect 389546 503286 389602 504086
rect 393962 503286 394018 504086
rect 398378 503286 398434 504086
rect 402794 503286 402850 504086
rect 407210 503286 407266 504086
rect 411534 503286 411590 504086
rect 415950 503286 416006 504086
rect 420366 503286 420422 504086
rect 424782 503286 424838 504086
rect 429198 503286 429254 504086
rect 433614 503286 433670 504086
rect 438030 503286 438086 504086
rect 442354 503286 442410 504086
rect 446770 503286 446826 504086
rect 451186 503286 451242 504086
rect 455602 503286 455658 504086
rect 460018 503286 460074 504086
rect 464434 503286 464490 504086
rect 468850 503286 468906 504086
rect 473174 503286 473230 504086
rect 477590 503286 477646 504086
rect 482006 503286 482062 504086
rect 486422 503286 486478 504086
rect 490838 503286 490894 504086
rect 495254 503286 495310 504086
rect 499670 503286 499726 504086
rect 478 0 534 800
rect 1490 0 1546 800
rect 2502 0 2558 800
rect 3514 0 3570 800
rect 4526 0 4582 800
rect 5538 0 5594 800
rect 6550 0 6606 800
rect 7562 0 7618 800
rect 8574 0 8630 800
rect 9586 0 9642 800
rect 10598 0 10654 800
rect 11610 0 11666 800
rect 12622 0 12678 800
rect 13634 0 13690 800
rect 14646 0 14702 800
rect 15750 0 15806 800
rect 16762 0 16818 800
rect 17774 0 17830 800
rect 18786 0 18842 800
rect 19798 0 19854 800
rect 20810 0 20866 800
rect 21822 0 21878 800
rect 22834 0 22890 800
rect 23846 0 23902 800
rect 24858 0 24914 800
rect 25870 0 25926 800
rect 26882 0 26938 800
rect 27894 0 27950 800
rect 28906 0 28962 800
rect 29918 0 29974 800
rect 31022 0 31078 800
rect 32034 0 32090 800
rect 33046 0 33102 800
rect 34058 0 34114 800
rect 35070 0 35126 800
rect 36082 0 36138 800
rect 37094 0 37150 800
rect 38106 0 38162 800
rect 39118 0 39174 800
rect 40130 0 40186 800
rect 41142 0 41198 800
rect 42154 0 42210 800
rect 43166 0 43222 800
rect 44178 0 44234 800
rect 45190 0 45246 800
rect 46294 0 46350 800
rect 47306 0 47362 800
rect 48318 0 48374 800
rect 49330 0 49386 800
rect 50342 0 50398 800
rect 51354 0 51410 800
rect 52366 0 52422 800
rect 53378 0 53434 800
rect 54390 0 54446 800
rect 55402 0 55458 800
rect 56414 0 56470 800
rect 57426 0 57482 800
rect 58438 0 58494 800
rect 59450 0 59506 800
rect 60462 0 60518 800
rect 61566 0 61622 800
rect 62578 0 62634 800
rect 63590 0 63646 800
rect 64602 0 64658 800
rect 65614 0 65670 800
rect 66626 0 66682 800
rect 67638 0 67694 800
rect 68650 0 68706 800
rect 69662 0 69718 800
rect 70674 0 70730 800
rect 71686 0 71742 800
rect 72698 0 72754 800
rect 73710 0 73766 800
rect 74722 0 74778 800
rect 75734 0 75790 800
rect 76838 0 76894 800
rect 77850 0 77906 800
rect 78862 0 78918 800
rect 79874 0 79930 800
rect 80886 0 80942 800
rect 81898 0 81954 800
rect 82910 0 82966 800
rect 83922 0 83978 800
rect 84934 0 84990 800
rect 85946 0 86002 800
rect 86958 0 87014 800
rect 87970 0 88026 800
rect 88982 0 89038 800
rect 89994 0 90050 800
rect 91006 0 91062 800
rect 92110 0 92166 800
rect 93122 0 93178 800
rect 94134 0 94190 800
rect 95146 0 95202 800
rect 96158 0 96214 800
rect 97170 0 97226 800
rect 98182 0 98238 800
rect 99194 0 99250 800
rect 100206 0 100262 800
rect 101218 0 101274 800
rect 102230 0 102286 800
rect 103242 0 103298 800
rect 104254 0 104310 800
rect 105266 0 105322 800
rect 106278 0 106334 800
rect 107382 0 107438 800
rect 108394 0 108450 800
rect 109406 0 109462 800
rect 110418 0 110474 800
rect 111430 0 111486 800
rect 112442 0 112498 800
rect 113454 0 113510 800
rect 114466 0 114522 800
rect 115478 0 115534 800
rect 116490 0 116546 800
rect 117502 0 117558 800
rect 118514 0 118570 800
rect 119526 0 119582 800
rect 120538 0 120594 800
rect 121550 0 121606 800
rect 122654 0 122710 800
rect 123666 0 123722 800
rect 124678 0 124734 800
rect 125690 0 125746 800
rect 126702 0 126758 800
rect 127714 0 127770 800
rect 128726 0 128782 800
rect 129738 0 129794 800
rect 130750 0 130806 800
rect 131762 0 131818 800
rect 132774 0 132830 800
rect 133786 0 133842 800
rect 134798 0 134854 800
rect 135810 0 135866 800
rect 136822 0 136878 800
rect 137926 0 137982 800
rect 138938 0 138994 800
rect 139950 0 140006 800
rect 140962 0 141018 800
rect 141974 0 142030 800
rect 142986 0 143042 800
rect 143998 0 144054 800
rect 145010 0 145066 800
rect 146022 0 146078 800
rect 147034 0 147090 800
rect 148046 0 148102 800
rect 149058 0 149114 800
rect 150070 0 150126 800
rect 151082 0 151138 800
rect 152094 0 152150 800
rect 153198 0 153254 800
rect 154210 0 154266 800
rect 155222 0 155278 800
rect 156234 0 156290 800
rect 157246 0 157302 800
rect 158258 0 158314 800
rect 159270 0 159326 800
rect 160282 0 160338 800
rect 161294 0 161350 800
rect 162306 0 162362 800
rect 163318 0 163374 800
rect 164330 0 164386 800
rect 165342 0 165398 800
rect 166354 0 166410 800
rect 167366 0 167422 800
rect 168470 0 168526 800
rect 169482 0 169538 800
rect 170494 0 170550 800
rect 171506 0 171562 800
rect 172518 0 172574 800
rect 173530 0 173586 800
rect 174542 0 174598 800
rect 175554 0 175610 800
rect 176566 0 176622 800
rect 177578 0 177634 800
rect 178590 0 178646 800
rect 179602 0 179658 800
rect 180614 0 180670 800
rect 181626 0 181682 800
rect 182638 0 182694 800
rect 183742 0 183798 800
rect 184754 0 184810 800
rect 185766 0 185822 800
rect 186778 0 186834 800
rect 187790 0 187846 800
rect 188802 0 188858 800
rect 189814 0 189870 800
rect 190826 0 190882 800
rect 191838 0 191894 800
rect 192850 0 192906 800
rect 193862 0 193918 800
rect 194874 0 194930 800
rect 195886 0 195942 800
rect 196898 0 196954 800
rect 197910 0 197966 800
rect 199014 0 199070 800
rect 200026 0 200082 800
rect 201038 0 201094 800
rect 202050 0 202106 800
rect 203062 0 203118 800
rect 204074 0 204130 800
rect 205086 0 205142 800
rect 206098 0 206154 800
rect 207110 0 207166 800
rect 208122 0 208178 800
rect 209134 0 209190 800
rect 210146 0 210202 800
rect 211158 0 211214 800
rect 212170 0 212226 800
rect 213182 0 213238 800
rect 214286 0 214342 800
rect 215298 0 215354 800
rect 216310 0 216366 800
rect 217322 0 217378 800
rect 218334 0 218390 800
rect 219346 0 219402 800
rect 220358 0 220414 800
rect 221370 0 221426 800
rect 222382 0 222438 800
rect 223394 0 223450 800
rect 224406 0 224462 800
rect 225418 0 225474 800
rect 226430 0 226486 800
rect 227442 0 227498 800
rect 228454 0 228510 800
rect 229558 0 229614 800
rect 230570 0 230626 800
rect 231582 0 231638 800
rect 232594 0 232650 800
rect 233606 0 233662 800
rect 234618 0 234674 800
rect 235630 0 235686 800
rect 236642 0 236698 800
rect 237654 0 237710 800
rect 238666 0 238722 800
rect 239678 0 239734 800
rect 240690 0 240746 800
rect 241702 0 241758 800
rect 242714 0 242770 800
rect 243726 0 243782 800
rect 244830 0 244886 800
rect 245842 0 245898 800
rect 246854 0 246910 800
rect 247866 0 247922 800
rect 248878 0 248934 800
rect 249890 0 249946 800
rect 250902 0 250958 800
rect 251914 0 251970 800
rect 252926 0 252982 800
rect 253938 0 253994 800
rect 254950 0 255006 800
rect 255962 0 256018 800
rect 256974 0 257030 800
rect 257986 0 258042 800
rect 259090 0 259146 800
rect 260102 0 260158 800
rect 261114 0 261170 800
rect 262126 0 262182 800
rect 263138 0 263194 800
rect 264150 0 264206 800
rect 265162 0 265218 800
rect 266174 0 266230 800
rect 267186 0 267242 800
rect 268198 0 268254 800
rect 269210 0 269266 800
rect 270222 0 270278 800
rect 271234 0 271290 800
rect 272246 0 272302 800
rect 273258 0 273314 800
rect 274362 0 274418 800
rect 275374 0 275430 800
rect 276386 0 276442 800
rect 277398 0 277454 800
rect 278410 0 278466 800
rect 279422 0 279478 800
rect 280434 0 280490 800
rect 281446 0 281502 800
rect 282458 0 282514 800
rect 283470 0 283526 800
rect 284482 0 284538 800
rect 285494 0 285550 800
rect 286506 0 286562 800
rect 287518 0 287574 800
rect 288530 0 288586 800
rect 289634 0 289690 800
rect 290646 0 290702 800
rect 291658 0 291714 800
rect 292670 0 292726 800
rect 293682 0 293738 800
rect 294694 0 294750 800
rect 295706 0 295762 800
rect 296718 0 296774 800
rect 297730 0 297786 800
rect 298742 0 298798 800
rect 299754 0 299810 800
rect 300766 0 300822 800
rect 301778 0 301834 800
rect 302790 0 302846 800
rect 303802 0 303858 800
rect 304906 0 304962 800
rect 305918 0 305974 800
rect 306930 0 306986 800
rect 307942 0 307998 800
rect 308954 0 309010 800
rect 309966 0 310022 800
rect 310978 0 311034 800
rect 311990 0 312046 800
rect 313002 0 313058 800
rect 314014 0 314070 800
rect 315026 0 315082 800
rect 316038 0 316094 800
rect 317050 0 317106 800
rect 318062 0 318118 800
rect 319074 0 319130 800
rect 320178 0 320234 800
rect 321190 0 321246 800
rect 322202 0 322258 800
rect 323214 0 323270 800
rect 324226 0 324282 800
rect 325238 0 325294 800
rect 326250 0 326306 800
rect 327262 0 327318 800
rect 328274 0 328330 800
rect 329286 0 329342 800
rect 330298 0 330354 800
rect 331310 0 331366 800
rect 332322 0 332378 800
rect 333334 0 333390 800
rect 334346 0 334402 800
rect 335450 0 335506 800
rect 336462 0 336518 800
rect 337474 0 337530 800
rect 338486 0 338542 800
rect 339498 0 339554 800
rect 340510 0 340566 800
rect 341522 0 341578 800
rect 342534 0 342590 800
rect 343546 0 343602 800
rect 344558 0 344614 800
rect 345570 0 345626 800
rect 346582 0 346638 800
rect 347594 0 347650 800
rect 348606 0 348662 800
rect 349618 0 349674 800
rect 350722 0 350778 800
rect 351734 0 351790 800
rect 352746 0 352802 800
rect 353758 0 353814 800
rect 354770 0 354826 800
rect 355782 0 355838 800
rect 356794 0 356850 800
rect 357806 0 357862 800
rect 358818 0 358874 800
rect 359830 0 359886 800
rect 360842 0 360898 800
rect 361854 0 361910 800
rect 362866 0 362922 800
rect 363878 0 363934 800
rect 364890 0 364946 800
rect 365994 0 366050 800
rect 367006 0 367062 800
rect 368018 0 368074 800
rect 369030 0 369086 800
rect 370042 0 370098 800
rect 371054 0 371110 800
rect 372066 0 372122 800
rect 373078 0 373134 800
rect 374090 0 374146 800
rect 375102 0 375158 800
rect 376114 0 376170 800
rect 377126 0 377182 800
rect 378138 0 378194 800
rect 379150 0 379206 800
rect 380162 0 380218 800
rect 381266 0 381322 800
rect 382278 0 382334 800
rect 383290 0 383346 800
rect 384302 0 384358 800
rect 385314 0 385370 800
rect 386326 0 386382 800
rect 387338 0 387394 800
rect 388350 0 388406 800
rect 389362 0 389418 800
rect 390374 0 390430 800
rect 391386 0 391442 800
rect 392398 0 392454 800
rect 393410 0 393466 800
rect 394422 0 394478 800
rect 395434 0 395490 800
rect 396538 0 396594 800
rect 397550 0 397606 800
rect 398562 0 398618 800
rect 399574 0 399630 800
rect 400586 0 400642 800
rect 401598 0 401654 800
rect 402610 0 402666 800
rect 403622 0 403678 800
rect 404634 0 404690 800
rect 405646 0 405702 800
rect 406658 0 406714 800
rect 407670 0 407726 800
rect 408682 0 408738 800
rect 409694 0 409750 800
rect 410706 0 410762 800
rect 411810 0 411866 800
rect 412822 0 412878 800
rect 413834 0 413890 800
rect 414846 0 414902 800
rect 415858 0 415914 800
rect 416870 0 416926 800
rect 417882 0 417938 800
rect 418894 0 418950 800
rect 419906 0 419962 800
rect 420918 0 420974 800
rect 421930 0 421986 800
rect 422942 0 422998 800
rect 423954 0 424010 800
rect 424966 0 425022 800
rect 425978 0 426034 800
rect 427082 0 427138 800
rect 428094 0 428150 800
rect 429106 0 429162 800
rect 430118 0 430174 800
rect 431130 0 431186 800
rect 432142 0 432198 800
rect 433154 0 433210 800
rect 434166 0 434222 800
rect 435178 0 435234 800
rect 436190 0 436246 800
rect 437202 0 437258 800
rect 438214 0 438270 800
rect 439226 0 439282 800
rect 440238 0 440294 800
rect 441250 0 441306 800
rect 442354 0 442410 800
rect 443366 0 443422 800
rect 444378 0 444434 800
rect 445390 0 445446 800
rect 446402 0 446458 800
rect 447414 0 447470 800
rect 448426 0 448482 800
rect 449438 0 449494 800
rect 450450 0 450506 800
rect 451462 0 451518 800
rect 452474 0 452530 800
rect 453486 0 453542 800
rect 454498 0 454554 800
rect 455510 0 455566 800
rect 456522 0 456578 800
rect 457626 0 457682 800
rect 458638 0 458694 800
rect 459650 0 459706 800
rect 460662 0 460718 800
rect 461674 0 461730 800
rect 462686 0 462742 800
rect 463698 0 463754 800
rect 464710 0 464766 800
rect 465722 0 465778 800
rect 466734 0 466790 800
rect 467746 0 467802 800
rect 468758 0 468814 800
rect 469770 0 469826 800
rect 470782 0 470838 800
rect 471794 0 471850 800
rect 472898 0 472954 800
rect 473910 0 473966 800
rect 474922 0 474978 800
rect 475934 0 475990 800
rect 476946 0 477002 800
rect 477958 0 478014 800
rect 478970 0 479026 800
rect 479982 0 480038 800
rect 480994 0 481050 800
rect 482006 0 482062 800
rect 483018 0 483074 800
rect 484030 0 484086 800
rect 485042 0 485098 800
rect 486054 0 486110 800
rect 487066 0 487122 800
rect 488170 0 488226 800
rect 489182 0 489238 800
rect 490194 0 490250 800
rect 491206 0 491262 800
rect 492218 0 492274 800
rect 493230 0 493286 800
rect 494242 0 494298 800
rect 495254 0 495310 800
rect 496266 0 496322 800
rect 497278 0 497334 800
rect 498290 0 498346 800
rect 499302 0 499358 800
rect 500314 0 500370 800
rect 501326 0 501382 800
<< obsm2 >>
rect 480 503230 2078 503286
rect 2246 503230 6402 503286
rect 6570 503230 10818 503286
rect 10986 503230 15234 503286
rect 15402 503230 19650 503286
rect 19818 503230 24066 503286
rect 24234 503230 28482 503286
rect 28650 503230 32898 503286
rect 33066 503230 37222 503286
rect 37390 503230 41638 503286
rect 41806 503230 46054 503286
rect 46222 503230 50470 503286
rect 50638 503230 54886 503286
rect 55054 503230 59302 503286
rect 59470 503230 63718 503286
rect 63886 503230 68042 503286
rect 68210 503230 72458 503286
rect 72626 503230 76874 503286
rect 77042 503230 81290 503286
rect 81458 503230 85706 503286
rect 85874 503230 90122 503286
rect 90290 503230 94538 503286
rect 94706 503230 98862 503286
rect 99030 503230 103278 503286
rect 103446 503230 107694 503286
rect 107862 503230 112110 503286
rect 112278 503230 116526 503286
rect 116694 503230 120942 503286
rect 121110 503230 125358 503286
rect 125526 503230 129682 503286
rect 129850 503230 134098 503286
rect 134266 503230 138514 503286
rect 138682 503230 142930 503286
rect 143098 503230 147346 503286
rect 147514 503230 151762 503286
rect 151930 503230 156178 503286
rect 156346 503230 160502 503286
rect 160670 503230 164918 503286
rect 165086 503230 169334 503286
rect 169502 503230 173750 503286
rect 173918 503230 178166 503286
rect 178334 503230 182582 503286
rect 182750 503230 186998 503286
rect 187166 503230 191322 503286
rect 191490 503230 195738 503286
rect 195906 503230 200154 503286
rect 200322 503230 204570 503286
rect 204738 503230 208986 503286
rect 209154 503230 213402 503286
rect 213570 503230 217818 503286
rect 217986 503230 222142 503286
rect 222310 503230 226558 503286
rect 226726 503230 230974 503286
rect 231142 503230 235390 503286
rect 235558 503230 239806 503286
rect 239974 503230 244222 503286
rect 244390 503230 248638 503286
rect 248806 503230 253054 503286
rect 253222 503230 257378 503286
rect 257546 503230 261794 503286
rect 261962 503230 266210 503286
rect 266378 503230 270626 503286
rect 270794 503230 275042 503286
rect 275210 503230 279458 503286
rect 279626 503230 283874 503286
rect 284042 503230 288198 503286
rect 288366 503230 292614 503286
rect 292782 503230 297030 503286
rect 297198 503230 301446 503286
rect 301614 503230 305862 503286
rect 306030 503230 310278 503286
rect 310446 503230 314694 503286
rect 314862 503230 319018 503286
rect 319186 503230 323434 503286
rect 323602 503230 327850 503286
rect 328018 503230 332266 503286
rect 332434 503230 336682 503286
rect 336850 503230 341098 503286
rect 341266 503230 345514 503286
rect 345682 503230 349838 503286
rect 350006 503230 354254 503286
rect 354422 503230 358670 503286
rect 358838 503230 363086 503286
rect 363254 503230 367502 503286
rect 367670 503230 371918 503286
rect 372086 503230 376334 503286
rect 376502 503230 380658 503286
rect 380826 503230 385074 503286
rect 385242 503230 389490 503286
rect 389658 503230 393906 503286
rect 394074 503230 398322 503286
rect 398490 503230 402738 503286
rect 402906 503230 407154 503286
rect 407322 503230 411478 503286
rect 411646 503230 415894 503286
rect 416062 503230 420310 503286
rect 420478 503230 424726 503286
rect 424894 503230 429142 503286
rect 429310 503230 433558 503286
rect 433726 503230 437974 503286
rect 438142 503230 442298 503286
rect 442466 503230 446714 503286
rect 446882 503230 451130 503286
rect 451298 503230 455546 503286
rect 455714 503230 459962 503286
rect 460130 503230 464378 503286
rect 464546 503230 468794 503286
rect 468962 503230 473118 503286
rect 473286 503230 477534 503286
rect 477702 503230 481950 503286
rect 482118 503230 486366 503286
rect 486534 503230 490782 503286
rect 490950 503230 495198 503286
rect 495366 503230 499614 503286
rect 499782 503230 501380 503286
rect 480 856 501380 503230
rect 590 2 1434 856
rect 1602 2 2446 856
rect 2614 2 3458 856
rect 3626 2 4470 856
rect 4638 2 5482 856
rect 5650 2 6494 856
rect 6662 2 7506 856
rect 7674 2 8518 856
rect 8686 2 9530 856
rect 9698 2 10542 856
rect 10710 2 11554 856
rect 11722 2 12566 856
rect 12734 2 13578 856
rect 13746 2 14590 856
rect 14758 2 15694 856
rect 15862 2 16706 856
rect 16874 2 17718 856
rect 17886 2 18730 856
rect 18898 2 19742 856
rect 19910 2 20754 856
rect 20922 2 21766 856
rect 21934 2 22778 856
rect 22946 2 23790 856
rect 23958 2 24802 856
rect 24970 2 25814 856
rect 25982 2 26826 856
rect 26994 2 27838 856
rect 28006 2 28850 856
rect 29018 2 29862 856
rect 30030 2 30966 856
rect 31134 2 31978 856
rect 32146 2 32990 856
rect 33158 2 34002 856
rect 34170 2 35014 856
rect 35182 2 36026 856
rect 36194 2 37038 856
rect 37206 2 38050 856
rect 38218 2 39062 856
rect 39230 2 40074 856
rect 40242 2 41086 856
rect 41254 2 42098 856
rect 42266 2 43110 856
rect 43278 2 44122 856
rect 44290 2 45134 856
rect 45302 2 46238 856
rect 46406 2 47250 856
rect 47418 2 48262 856
rect 48430 2 49274 856
rect 49442 2 50286 856
rect 50454 2 51298 856
rect 51466 2 52310 856
rect 52478 2 53322 856
rect 53490 2 54334 856
rect 54502 2 55346 856
rect 55514 2 56358 856
rect 56526 2 57370 856
rect 57538 2 58382 856
rect 58550 2 59394 856
rect 59562 2 60406 856
rect 60574 2 61510 856
rect 61678 2 62522 856
rect 62690 2 63534 856
rect 63702 2 64546 856
rect 64714 2 65558 856
rect 65726 2 66570 856
rect 66738 2 67582 856
rect 67750 2 68594 856
rect 68762 2 69606 856
rect 69774 2 70618 856
rect 70786 2 71630 856
rect 71798 2 72642 856
rect 72810 2 73654 856
rect 73822 2 74666 856
rect 74834 2 75678 856
rect 75846 2 76782 856
rect 76950 2 77794 856
rect 77962 2 78806 856
rect 78974 2 79818 856
rect 79986 2 80830 856
rect 80998 2 81842 856
rect 82010 2 82854 856
rect 83022 2 83866 856
rect 84034 2 84878 856
rect 85046 2 85890 856
rect 86058 2 86902 856
rect 87070 2 87914 856
rect 88082 2 88926 856
rect 89094 2 89938 856
rect 90106 2 90950 856
rect 91118 2 92054 856
rect 92222 2 93066 856
rect 93234 2 94078 856
rect 94246 2 95090 856
rect 95258 2 96102 856
rect 96270 2 97114 856
rect 97282 2 98126 856
rect 98294 2 99138 856
rect 99306 2 100150 856
rect 100318 2 101162 856
rect 101330 2 102174 856
rect 102342 2 103186 856
rect 103354 2 104198 856
rect 104366 2 105210 856
rect 105378 2 106222 856
rect 106390 2 107326 856
rect 107494 2 108338 856
rect 108506 2 109350 856
rect 109518 2 110362 856
rect 110530 2 111374 856
rect 111542 2 112386 856
rect 112554 2 113398 856
rect 113566 2 114410 856
rect 114578 2 115422 856
rect 115590 2 116434 856
rect 116602 2 117446 856
rect 117614 2 118458 856
rect 118626 2 119470 856
rect 119638 2 120482 856
rect 120650 2 121494 856
rect 121662 2 122598 856
rect 122766 2 123610 856
rect 123778 2 124622 856
rect 124790 2 125634 856
rect 125802 2 126646 856
rect 126814 2 127658 856
rect 127826 2 128670 856
rect 128838 2 129682 856
rect 129850 2 130694 856
rect 130862 2 131706 856
rect 131874 2 132718 856
rect 132886 2 133730 856
rect 133898 2 134742 856
rect 134910 2 135754 856
rect 135922 2 136766 856
rect 136934 2 137870 856
rect 138038 2 138882 856
rect 139050 2 139894 856
rect 140062 2 140906 856
rect 141074 2 141918 856
rect 142086 2 142930 856
rect 143098 2 143942 856
rect 144110 2 144954 856
rect 145122 2 145966 856
rect 146134 2 146978 856
rect 147146 2 147990 856
rect 148158 2 149002 856
rect 149170 2 150014 856
rect 150182 2 151026 856
rect 151194 2 152038 856
rect 152206 2 153142 856
rect 153310 2 154154 856
rect 154322 2 155166 856
rect 155334 2 156178 856
rect 156346 2 157190 856
rect 157358 2 158202 856
rect 158370 2 159214 856
rect 159382 2 160226 856
rect 160394 2 161238 856
rect 161406 2 162250 856
rect 162418 2 163262 856
rect 163430 2 164274 856
rect 164442 2 165286 856
rect 165454 2 166298 856
rect 166466 2 167310 856
rect 167478 2 168414 856
rect 168582 2 169426 856
rect 169594 2 170438 856
rect 170606 2 171450 856
rect 171618 2 172462 856
rect 172630 2 173474 856
rect 173642 2 174486 856
rect 174654 2 175498 856
rect 175666 2 176510 856
rect 176678 2 177522 856
rect 177690 2 178534 856
rect 178702 2 179546 856
rect 179714 2 180558 856
rect 180726 2 181570 856
rect 181738 2 182582 856
rect 182750 2 183686 856
rect 183854 2 184698 856
rect 184866 2 185710 856
rect 185878 2 186722 856
rect 186890 2 187734 856
rect 187902 2 188746 856
rect 188914 2 189758 856
rect 189926 2 190770 856
rect 190938 2 191782 856
rect 191950 2 192794 856
rect 192962 2 193806 856
rect 193974 2 194818 856
rect 194986 2 195830 856
rect 195998 2 196842 856
rect 197010 2 197854 856
rect 198022 2 198958 856
rect 199126 2 199970 856
rect 200138 2 200982 856
rect 201150 2 201994 856
rect 202162 2 203006 856
rect 203174 2 204018 856
rect 204186 2 205030 856
rect 205198 2 206042 856
rect 206210 2 207054 856
rect 207222 2 208066 856
rect 208234 2 209078 856
rect 209246 2 210090 856
rect 210258 2 211102 856
rect 211270 2 212114 856
rect 212282 2 213126 856
rect 213294 2 214230 856
rect 214398 2 215242 856
rect 215410 2 216254 856
rect 216422 2 217266 856
rect 217434 2 218278 856
rect 218446 2 219290 856
rect 219458 2 220302 856
rect 220470 2 221314 856
rect 221482 2 222326 856
rect 222494 2 223338 856
rect 223506 2 224350 856
rect 224518 2 225362 856
rect 225530 2 226374 856
rect 226542 2 227386 856
rect 227554 2 228398 856
rect 228566 2 229502 856
rect 229670 2 230514 856
rect 230682 2 231526 856
rect 231694 2 232538 856
rect 232706 2 233550 856
rect 233718 2 234562 856
rect 234730 2 235574 856
rect 235742 2 236586 856
rect 236754 2 237598 856
rect 237766 2 238610 856
rect 238778 2 239622 856
rect 239790 2 240634 856
rect 240802 2 241646 856
rect 241814 2 242658 856
rect 242826 2 243670 856
rect 243838 2 244774 856
rect 244942 2 245786 856
rect 245954 2 246798 856
rect 246966 2 247810 856
rect 247978 2 248822 856
rect 248990 2 249834 856
rect 250002 2 250846 856
rect 251014 2 251858 856
rect 252026 2 252870 856
rect 253038 2 253882 856
rect 254050 2 254894 856
rect 255062 2 255906 856
rect 256074 2 256918 856
rect 257086 2 257930 856
rect 258098 2 259034 856
rect 259202 2 260046 856
rect 260214 2 261058 856
rect 261226 2 262070 856
rect 262238 2 263082 856
rect 263250 2 264094 856
rect 264262 2 265106 856
rect 265274 2 266118 856
rect 266286 2 267130 856
rect 267298 2 268142 856
rect 268310 2 269154 856
rect 269322 2 270166 856
rect 270334 2 271178 856
rect 271346 2 272190 856
rect 272358 2 273202 856
rect 273370 2 274306 856
rect 274474 2 275318 856
rect 275486 2 276330 856
rect 276498 2 277342 856
rect 277510 2 278354 856
rect 278522 2 279366 856
rect 279534 2 280378 856
rect 280546 2 281390 856
rect 281558 2 282402 856
rect 282570 2 283414 856
rect 283582 2 284426 856
rect 284594 2 285438 856
rect 285606 2 286450 856
rect 286618 2 287462 856
rect 287630 2 288474 856
rect 288642 2 289578 856
rect 289746 2 290590 856
rect 290758 2 291602 856
rect 291770 2 292614 856
rect 292782 2 293626 856
rect 293794 2 294638 856
rect 294806 2 295650 856
rect 295818 2 296662 856
rect 296830 2 297674 856
rect 297842 2 298686 856
rect 298854 2 299698 856
rect 299866 2 300710 856
rect 300878 2 301722 856
rect 301890 2 302734 856
rect 302902 2 303746 856
rect 303914 2 304850 856
rect 305018 2 305862 856
rect 306030 2 306874 856
rect 307042 2 307886 856
rect 308054 2 308898 856
rect 309066 2 309910 856
rect 310078 2 310922 856
rect 311090 2 311934 856
rect 312102 2 312946 856
rect 313114 2 313958 856
rect 314126 2 314970 856
rect 315138 2 315982 856
rect 316150 2 316994 856
rect 317162 2 318006 856
rect 318174 2 319018 856
rect 319186 2 320122 856
rect 320290 2 321134 856
rect 321302 2 322146 856
rect 322314 2 323158 856
rect 323326 2 324170 856
rect 324338 2 325182 856
rect 325350 2 326194 856
rect 326362 2 327206 856
rect 327374 2 328218 856
rect 328386 2 329230 856
rect 329398 2 330242 856
rect 330410 2 331254 856
rect 331422 2 332266 856
rect 332434 2 333278 856
rect 333446 2 334290 856
rect 334458 2 335394 856
rect 335562 2 336406 856
rect 336574 2 337418 856
rect 337586 2 338430 856
rect 338598 2 339442 856
rect 339610 2 340454 856
rect 340622 2 341466 856
rect 341634 2 342478 856
rect 342646 2 343490 856
rect 343658 2 344502 856
rect 344670 2 345514 856
rect 345682 2 346526 856
rect 346694 2 347538 856
rect 347706 2 348550 856
rect 348718 2 349562 856
rect 349730 2 350666 856
rect 350834 2 351678 856
rect 351846 2 352690 856
rect 352858 2 353702 856
rect 353870 2 354714 856
rect 354882 2 355726 856
rect 355894 2 356738 856
rect 356906 2 357750 856
rect 357918 2 358762 856
rect 358930 2 359774 856
rect 359942 2 360786 856
rect 360954 2 361798 856
rect 361966 2 362810 856
rect 362978 2 363822 856
rect 363990 2 364834 856
rect 365002 2 365938 856
rect 366106 2 366950 856
rect 367118 2 367962 856
rect 368130 2 368974 856
rect 369142 2 369986 856
rect 370154 2 370998 856
rect 371166 2 372010 856
rect 372178 2 373022 856
rect 373190 2 374034 856
rect 374202 2 375046 856
rect 375214 2 376058 856
rect 376226 2 377070 856
rect 377238 2 378082 856
rect 378250 2 379094 856
rect 379262 2 380106 856
rect 380274 2 381210 856
rect 381378 2 382222 856
rect 382390 2 383234 856
rect 383402 2 384246 856
rect 384414 2 385258 856
rect 385426 2 386270 856
rect 386438 2 387282 856
rect 387450 2 388294 856
rect 388462 2 389306 856
rect 389474 2 390318 856
rect 390486 2 391330 856
rect 391498 2 392342 856
rect 392510 2 393354 856
rect 393522 2 394366 856
rect 394534 2 395378 856
rect 395546 2 396482 856
rect 396650 2 397494 856
rect 397662 2 398506 856
rect 398674 2 399518 856
rect 399686 2 400530 856
rect 400698 2 401542 856
rect 401710 2 402554 856
rect 402722 2 403566 856
rect 403734 2 404578 856
rect 404746 2 405590 856
rect 405758 2 406602 856
rect 406770 2 407614 856
rect 407782 2 408626 856
rect 408794 2 409638 856
rect 409806 2 410650 856
rect 410818 2 411754 856
rect 411922 2 412766 856
rect 412934 2 413778 856
rect 413946 2 414790 856
rect 414958 2 415802 856
rect 415970 2 416814 856
rect 416982 2 417826 856
rect 417994 2 418838 856
rect 419006 2 419850 856
rect 420018 2 420862 856
rect 421030 2 421874 856
rect 422042 2 422886 856
rect 423054 2 423898 856
rect 424066 2 424910 856
rect 425078 2 425922 856
rect 426090 2 427026 856
rect 427194 2 428038 856
rect 428206 2 429050 856
rect 429218 2 430062 856
rect 430230 2 431074 856
rect 431242 2 432086 856
rect 432254 2 433098 856
rect 433266 2 434110 856
rect 434278 2 435122 856
rect 435290 2 436134 856
rect 436302 2 437146 856
rect 437314 2 438158 856
rect 438326 2 439170 856
rect 439338 2 440182 856
rect 440350 2 441194 856
rect 441362 2 442298 856
rect 442466 2 443310 856
rect 443478 2 444322 856
rect 444490 2 445334 856
rect 445502 2 446346 856
rect 446514 2 447358 856
rect 447526 2 448370 856
rect 448538 2 449382 856
rect 449550 2 450394 856
rect 450562 2 451406 856
rect 451574 2 452418 856
rect 452586 2 453430 856
rect 453598 2 454442 856
rect 454610 2 455454 856
rect 455622 2 456466 856
rect 456634 2 457570 856
rect 457738 2 458582 856
rect 458750 2 459594 856
rect 459762 2 460606 856
rect 460774 2 461618 856
rect 461786 2 462630 856
rect 462798 2 463642 856
rect 463810 2 464654 856
rect 464822 2 465666 856
rect 465834 2 466678 856
rect 466846 2 467690 856
rect 467858 2 468702 856
rect 468870 2 469714 856
rect 469882 2 470726 856
rect 470894 2 471738 856
rect 471906 2 472842 856
rect 473010 2 473854 856
rect 474022 2 474866 856
rect 475034 2 475878 856
rect 476046 2 476890 856
rect 477058 2 477902 856
rect 478070 2 478914 856
rect 479082 2 479926 856
rect 480094 2 480938 856
rect 481106 2 481950 856
rect 482118 2 482962 856
rect 483130 2 483974 856
rect 484142 2 484986 856
rect 485154 2 485998 856
rect 486166 2 487010 856
rect 487178 2 488114 856
rect 488282 2 489126 856
rect 489294 2 490138 856
rect 490306 2 491150 856
rect 491318 2 492162 856
rect 492330 2 493174 856
rect 493342 2 494186 856
rect 494354 2 495198 856
rect 495366 2 496210 856
rect 496378 2 497222 856
rect 497390 2 498234 856
rect 498402 2 499246 856
rect 499414 2 500258 856
rect 500426 2 501270 856
<< obsm3 >>
rect 3969 171 496048 501601
<< metal4 >>
rect 4208 2128 4528 501616
rect 19568 2128 19888 501616
rect 34928 2128 35248 501616
rect 50288 2128 50608 501616
rect 65648 2128 65968 501616
rect 81008 2128 81328 501616
rect 96368 2128 96688 501616
rect 111728 2128 112048 501616
rect 127088 2128 127408 501616
rect 142448 2128 142768 501616
rect 157808 2128 158128 501616
rect 173168 2128 173488 501616
rect 188528 2128 188848 501616
rect 203888 2128 204208 501616
rect 219248 2128 219568 501616
rect 234608 2128 234928 501616
rect 249968 2128 250288 501616
rect 265328 2128 265648 501616
rect 280688 2128 281008 501616
rect 296048 2128 296368 501616
rect 311408 2128 311728 501616
rect 326768 2128 327088 501616
rect 342128 2128 342448 501616
rect 357488 2128 357808 501616
rect 372848 2128 373168 501616
rect 388208 2128 388528 501616
rect 403568 2128 403888 501616
rect 418928 2128 419248 501616
rect 434288 2128 434608 501616
rect 449648 2128 449968 501616
rect 465008 2128 465328 501616
rect 480368 2128 480688 501616
rect 495728 2128 496048 501616
<< obsm4 >>
rect 19379 2048 19488 501397
rect 19968 2048 34848 501397
rect 35328 2048 50208 501397
rect 50688 2048 65568 501397
rect 66048 2048 80928 501397
rect 81408 2048 96288 501397
rect 96768 2048 111648 501397
rect 112128 2048 127008 501397
rect 127488 2048 142368 501397
rect 142848 2048 157728 501397
rect 158208 2048 173088 501397
rect 173568 2048 188448 501397
rect 188928 2048 203808 501397
rect 204288 2048 219168 501397
rect 219648 2048 234528 501397
rect 235008 2048 249888 501397
rect 250368 2048 265248 501397
rect 265728 2048 280608 501397
rect 281088 2048 295968 501397
rect 296448 2048 311328 501397
rect 311808 2048 326688 501397
rect 327168 2048 342048 501397
rect 342528 2048 357408 501397
rect 357888 2048 372768 501397
rect 373248 2048 388128 501397
rect 388608 2048 403488 501397
rect 403968 2048 418848 501397
rect 419328 2048 434208 501397
rect 434688 2048 449568 501397
rect 450048 2048 464928 501397
rect 465408 2048 475949 501397
rect 19379 1395 475949 2048
<< labels >>
rlabel metal2 s 2134 503286 2190 504086 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 134154 503286 134210 504086 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 147402 503286 147458 504086 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 160558 503286 160614 504086 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 173806 503286 173862 504086 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 187054 503286 187110 504086 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 200210 503286 200266 504086 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 213458 503286 213514 504086 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 226614 503286 226670 504086 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 239862 503286 239918 504086 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 253110 503286 253166 504086 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 15290 503286 15346 504086 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 266266 503286 266322 504086 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 279514 503286 279570 504086 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 292670 503286 292726 504086 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 305918 503286 305974 504086 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 319074 503286 319130 504086 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 332322 503286 332378 504086 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 345570 503286 345626 504086 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 358726 503286 358782 504086 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 371974 503286 372030 504086 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 385130 503286 385186 504086 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 28538 503286 28594 504086 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 398378 503286 398434 504086 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 411534 503286 411590 504086 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 424782 503286 424838 504086 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 438030 503286 438086 504086 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 451186 503286 451242 504086 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 464434 503286 464490 504086 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 477590 503286 477646 504086 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 490838 503286 490894 504086 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 41694 503286 41750 504086 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 54942 503286 54998 504086 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 68098 503286 68154 504086 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 81346 503286 81402 504086 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 94594 503286 94650 504086 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 107750 503286 107806 504086 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 120998 503286 121054 504086 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6458 503286 6514 504086 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 138570 503286 138626 504086 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 151818 503286 151874 504086 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 164974 503286 165030 504086 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 178222 503286 178278 504086 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 191378 503286 191434 504086 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 204626 503286 204682 504086 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 217874 503286 217930 504086 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 231030 503286 231086 504086 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 244278 503286 244334 504086 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 257434 503286 257490 504086 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 19706 503286 19762 504086 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 270682 503286 270738 504086 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 283930 503286 283986 504086 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 297086 503286 297142 504086 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 310334 503286 310390 504086 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 323490 503286 323546 504086 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 336738 503286 336794 504086 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 349894 503286 349950 504086 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 363142 503286 363198 504086 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 376390 503286 376446 504086 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 389546 503286 389602 504086 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 32954 503286 33010 504086 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 402794 503286 402850 504086 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 415950 503286 416006 504086 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 429198 503286 429254 504086 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 442354 503286 442410 504086 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 455602 503286 455658 504086 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 468850 503286 468906 504086 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 482006 503286 482062 504086 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 495254 503286 495310 504086 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 46110 503286 46166 504086 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 59358 503286 59414 504086 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 72514 503286 72570 504086 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 85762 503286 85818 504086 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 98918 503286 98974 504086 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 112166 503286 112222 504086 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 125414 503286 125470 504086 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 10874 503286 10930 504086 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 142986 503286 143042 504086 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 156234 503286 156290 504086 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 169390 503286 169446 504086 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 182638 503286 182694 504086 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 195794 503286 195850 504086 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 209042 503286 209098 504086 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 222198 503286 222254 504086 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 235446 503286 235502 504086 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 248694 503286 248750 504086 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 261850 503286 261906 504086 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 24122 503286 24178 504086 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 275098 503286 275154 504086 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 288254 503286 288310 504086 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 301502 503286 301558 504086 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 314750 503286 314806 504086 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 327906 503286 327962 504086 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 341154 503286 341210 504086 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 354310 503286 354366 504086 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 367558 503286 367614 504086 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 380714 503286 380770 504086 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 393962 503286 394018 504086 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 37278 503286 37334 504086 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 407210 503286 407266 504086 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 420366 503286 420422 504086 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 433614 503286 433670 504086 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 446770 503286 446826 504086 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 460018 503286 460074 504086 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 473174 503286 473230 504086 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 486422 503286 486478 504086 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 499670 503286 499726 504086 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 50526 503286 50582 504086 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 63774 503286 63830 504086 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 76930 503286 76986 504086 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 90178 503286 90234 504086 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 103334 503286 103390 504086 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 116582 503286 116638 504086 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 129738 503286 129794 504086 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 499302 0 499358 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 500314 0 500370 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 501326 0 501382 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 413834 0 413890 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 416870 0 416926 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 419906 0 419962 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 422942 0 422998 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 425978 0 426034 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 429106 0 429162 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 432142 0 432198 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 435178 0 435234 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 438214 0 438270 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 441250 0 441306 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 444378 0 444434 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 447414 0 447470 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 450450 0 450506 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 453486 0 453542 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 456522 0 456578 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 459650 0 459706 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 462686 0 462742 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 465722 0 465778 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 468758 0 468814 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 471794 0 471850 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 474922 0 474978 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 477958 0 478014 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 480994 0 481050 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 484030 0 484086 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 487066 0 487122 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 490194 0 490250 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 493230 0 493286 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 496266 0 496322 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 184754 0 184810 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 200026 0 200082 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 209134 0 209190 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 212170 0 212226 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 215298 0 215354 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 221370 0 221426 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 224406 0 224462 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 230570 0 230626 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 233606 0 233662 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 242714 0 242770 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 245842 0 245898 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 248878 0 248934 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 251914 0 251970 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 254950 0 255006 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 257986 0 258042 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 264150 0 264206 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 267186 0 267242 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 270222 0 270278 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 273258 0 273314 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 276386 0 276442 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 279422 0 279478 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 282458 0 282514 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 285494 0 285550 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 288530 0 288586 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 291658 0 291714 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 294694 0 294750 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 297730 0 297786 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 300766 0 300822 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 303802 0 303858 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 306930 0 306986 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 309966 0 310022 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 313002 0 313058 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 316038 0 316094 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 319074 0 319130 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 322202 0 322258 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 325238 0 325294 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 328274 0 328330 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 331310 0 331366 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 334346 0 334402 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 337474 0 337530 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 340510 0 340566 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 343546 0 343602 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 346582 0 346638 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 349618 0 349674 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 352746 0 352802 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 355782 0 355838 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 358818 0 358874 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 361854 0 361910 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 364890 0 364946 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 368018 0 368074 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 371054 0 371110 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 374090 0 374146 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 377126 0 377182 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 380162 0 380218 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 383290 0 383346 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 386326 0 386382 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 389362 0 389418 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 392398 0 392454 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 395434 0 395490 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 398562 0 398618 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 401598 0 401654 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 404634 0 404690 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 407670 0 407726 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 410706 0 410762 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 414846 0 414902 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 417882 0 417938 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 420918 0 420974 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 423954 0 424010 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 427082 0 427138 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 430118 0 430174 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 433154 0 433210 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 436190 0 436246 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 439226 0 439282 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 442354 0 442410 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 445390 0 445446 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 448426 0 448482 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 451462 0 451518 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 454498 0 454554 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 457626 0 457682 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 460662 0 460718 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 463698 0 463754 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 466734 0 466790 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 469770 0 469826 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 472898 0 472954 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 475934 0 475990 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 478970 0 479026 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 482006 0 482062 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 485042 0 485098 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 488170 0 488226 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 491206 0 491262 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 494242 0 494298 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 497278 0 497334 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 149058 0 149114 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 152094 0 152150 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 158258 0 158314 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 161294 0 161350 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 167366 0 167422 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 112442 0 112498 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 170494 0 170550 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 179602 0 179658 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 182638 0 182694 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 185766 0 185822 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 188802 0 188858 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 191838 0 191894 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 197910 0 197966 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 207110 0 207166 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 210146 0 210202 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 213182 0 213238 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 216310 0 216366 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 219346 0 219402 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 222382 0 222438 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 225418 0 225474 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 228454 0 228510 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 231582 0 231638 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 234618 0 234674 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 237654 0 237710 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 240690 0 240746 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 243726 0 243782 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 246854 0 246910 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 249890 0 249946 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 252926 0 252982 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 255962 0 256018 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 259090 0 259146 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 121550 0 121606 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 262126 0 262182 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 265162 0 265218 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 268198 0 268254 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 271234 0 271290 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 274362 0 274418 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 277398 0 277454 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 280434 0 280490 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 283470 0 283526 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 286506 0 286562 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 289634 0 289690 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 292670 0 292726 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 295706 0 295762 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 298742 0 298798 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 301778 0 301834 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 304906 0 304962 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 307942 0 307998 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 310978 0 311034 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 314014 0 314070 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 317050 0 317106 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 320178 0 320234 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 323214 0 323270 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 326250 0 326306 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 329286 0 329342 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 332322 0 332378 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 335450 0 335506 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 338486 0 338542 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 341522 0 341578 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 344558 0 344614 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 347594 0 347650 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 350722 0 350778 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 353758 0 353814 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 356794 0 356850 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 359830 0 359886 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 362866 0 362922 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 365994 0 366050 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 369030 0 369086 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 372066 0 372122 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 375102 0 375158 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 378138 0 378194 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 381266 0 381322 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 133786 0 133842 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 384302 0 384358 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 387338 0 387394 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 390374 0 390430 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 393410 0 393466 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 396538 0 396594 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 399574 0 399630 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 402610 0 402666 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 405646 0 405702 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 408682 0 408738 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 411810 0 411866 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 415858 0 415914 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 418894 0 418950 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 421930 0 421986 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 424966 0 425022 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 428094 0 428150 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 431130 0 431186 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 434166 0 434222 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 437202 0 437258 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 440238 0 440294 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 443366 0 443422 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 446402 0 446458 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 449438 0 449494 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 452474 0 452530 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 455510 0 455566 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 458638 0 458694 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 461674 0 461730 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 464710 0 464766 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 467746 0 467802 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 470782 0 470838 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 473910 0 473966 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 476946 0 477002 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 479982 0 480038 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 483018 0 483074 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 486054 0 486110 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 489182 0 489238 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 492218 0 492274 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 495254 0 495310 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 498290 0 498346 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 165342 0 165398 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 192850 0 192906 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 199014 0 199070 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 202050 0 202106 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 205086 0 205142 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 208122 0 208178 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 211158 0 211214 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 214286 0 214342 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 217322 0 217378 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 223394 0 223450 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 226430 0 226486 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 229558 0 229614 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 232594 0 232650 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 238666 0 238722 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 247866 0 247922 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 250902 0 250958 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 253938 0 253994 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 256974 0 257030 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 263138 0 263194 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 266174 0 266230 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 272246 0 272302 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 275374 0 275430 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 278410 0 278466 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 281446 0 281502 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 284482 0 284538 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 287518 0 287574 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 290646 0 290702 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 293682 0 293738 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 296718 0 296774 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 299754 0 299810 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 305918 0 305974 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 308954 0 309010 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 311990 0 312046 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 315026 0 315082 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 318062 0 318118 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 321190 0 321246 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 324226 0 324282 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 327262 0 327318 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 330298 0 330354 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 333334 0 333390 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 336462 0 336518 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 339498 0 339554 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 342534 0 342590 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 345570 0 345626 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 348606 0 348662 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 351734 0 351790 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 354770 0 354826 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 357806 0 357862 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 360842 0 360898 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 363878 0 363934 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 367006 0 367062 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 370042 0 370098 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 373078 0 373134 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 376114 0 376170 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 379150 0 379206 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 382278 0 382334 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 385314 0 385370 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 388350 0 388406 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 391386 0 391442 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 394422 0 394478 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 397550 0 397606 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 400586 0 400642 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 403622 0 403678 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 406658 0 406714 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 409694 0 409750 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 412822 0 412878 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 434288 2128 434608 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 465008 2128 465328 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 495728 2128 496048 501616 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 418928 2128 419248 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 449648 2128 449968 501616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 480368 2128 480688 501616 6 vssd1
port 503 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 501942 504086
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 482293310
string GDS_START 1802832
<< end >>

