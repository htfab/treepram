magic
tech sky130A
magscale 1 2
timestamp 1635542372
<< obsli1 >>
rect 1104 17 574603 692529
<< obsm1 >>
rect 566 8 574618 692560
<< metal2 >>
rect 2502 694400 2558 695200
rect 7470 694400 7526 695200
rect 12530 694400 12586 695200
rect 17590 694400 17646 695200
rect 22650 694400 22706 695200
rect 27710 694400 27766 695200
rect 32770 694400 32826 695200
rect 37738 694400 37794 695200
rect 42798 694400 42854 695200
rect 47858 694400 47914 695200
rect 52918 694400 52974 695200
rect 57978 694400 58034 695200
rect 63038 694400 63094 695200
rect 68006 694400 68062 695200
rect 73066 694400 73122 695200
rect 78126 694400 78182 695200
rect 83186 694400 83242 695200
rect 88246 694400 88302 695200
rect 93306 694400 93362 695200
rect 98366 694400 98422 695200
rect 103334 694400 103390 695200
rect 108394 694400 108450 695200
rect 113454 694400 113510 695200
rect 118514 694400 118570 695200
rect 123574 694400 123630 695200
rect 128634 694400 128690 695200
rect 133602 694400 133658 695200
rect 138662 694400 138718 695200
rect 143722 694400 143778 695200
rect 148782 694400 148838 695200
rect 153842 694400 153898 695200
rect 158902 694400 158958 695200
rect 163870 694400 163926 695200
rect 168930 694400 168986 695200
rect 173990 694400 174046 695200
rect 179050 694400 179106 695200
rect 184110 694400 184166 695200
rect 189170 694400 189226 695200
rect 194230 694400 194286 695200
rect 199198 694400 199254 695200
rect 204258 694400 204314 695200
rect 209318 694400 209374 695200
rect 214378 694400 214434 695200
rect 219438 694400 219494 695200
rect 224498 694400 224554 695200
rect 229466 694400 229522 695200
rect 234526 694400 234582 695200
rect 239586 694400 239642 695200
rect 244646 694400 244702 695200
rect 249706 694400 249762 695200
rect 254766 694400 254822 695200
rect 259734 694400 259790 695200
rect 264794 694400 264850 695200
rect 269854 694400 269910 695200
rect 274914 694400 274970 695200
rect 279974 694400 280030 695200
rect 285034 694400 285090 695200
rect 290094 694400 290150 695200
rect 295062 694400 295118 695200
rect 300122 694400 300178 695200
rect 305182 694400 305238 695200
rect 310242 694400 310298 695200
rect 315302 694400 315358 695200
rect 320362 694400 320418 695200
rect 325330 694400 325386 695200
rect 330390 694400 330446 695200
rect 335450 694400 335506 695200
rect 340510 694400 340566 695200
rect 345570 694400 345626 695200
rect 350630 694400 350686 695200
rect 355598 694400 355654 695200
rect 360658 694400 360714 695200
rect 365718 694400 365774 695200
rect 370778 694400 370834 695200
rect 375838 694400 375894 695200
rect 380898 694400 380954 695200
rect 385958 694400 386014 695200
rect 390926 694400 390982 695200
rect 395986 694400 396042 695200
rect 401046 694400 401102 695200
rect 406106 694400 406162 695200
rect 411166 694400 411222 695200
rect 416226 694400 416282 695200
rect 421194 694400 421250 695200
rect 426254 694400 426310 695200
rect 431314 694400 431370 695200
rect 436374 694400 436430 695200
rect 441434 694400 441490 695200
rect 446494 694400 446550 695200
rect 451462 694400 451518 695200
rect 456522 694400 456578 695200
rect 461582 694400 461638 695200
rect 466642 694400 466698 695200
rect 471702 694400 471758 695200
rect 476762 694400 476818 695200
rect 481822 694400 481878 695200
rect 486790 694400 486846 695200
rect 491850 694400 491906 695200
rect 496910 694400 496966 695200
rect 501970 694400 502026 695200
rect 507030 694400 507086 695200
rect 512090 694400 512146 695200
rect 517058 694400 517114 695200
rect 522118 694400 522174 695200
rect 527178 694400 527234 695200
rect 532238 694400 532294 695200
rect 537298 694400 537354 695200
rect 542358 694400 542414 695200
rect 547326 694400 547382 695200
rect 552386 694400 552442 695200
rect 557446 694400 557502 695200
rect 562506 694400 562562 695200
rect 567566 694400 567622 695200
rect 572626 694400 572682 695200
rect 570 0 626 800
rect 1674 0 1730 800
rect 2870 0 2926 800
rect 4066 0 4122 800
rect 5170 0 5226 800
rect 6366 0 6422 800
rect 7562 0 7618 800
rect 8666 0 8722 800
rect 9862 0 9918 800
rect 11058 0 11114 800
rect 12162 0 12218 800
rect 13358 0 13414 800
rect 14554 0 14610 800
rect 15658 0 15714 800
rect 16854 0 16910 800
rect 18050 0 18106 800
rect 19154 0 19210 800
rect 20350 0 20406 800
rect 21546 0 21602 800
rect 22650 0 22706 800
rect 23846 0 23902 800
rect 25042 0 25098 800
rect 26146 0 26202 800
rect 27342 0 27398 800
rect 28538 0 28594 800
rect 29734 0 29790 800
rect 30838 0 30894 800
rect 32034 0 32090 800
rect 33230 0 33286 800
rect 34334 0 34390 800
rect 35530 0 35586 800
rect 36726 0 36782 800
rect 37830 0 37886 800
rect 39026 0 39082 800
rect 40222 0 40278 800
rect 41326 0 41382 800
rect 42522 0 42578 800
rect 43718 0 43774 800
rect 44822 0 44878 800
rect 46018 0 46074 800
rect 47214 0 47270 800
rect 48318 0 48374 800
rect 49514 0 49570 800
rect 50710 0 50766 800
rect 51814 0 51870 800
rect 53010 0 53066 800
rect 54206 0 54262 800
rect 55402 0 55458 800
rect 56506 0 56562 800
rect 57702 0 57758 800
rect 58898 0 58954 800
rect 60002 0 60058 800
rect 61198 0 61254 800
rect 62394 0 62450 800
rect 63498 0 63554 800
rect 64694 0 64750 800
rect 65890 0 65946 800
rect 66994 0 67050 800
rect 68190 0 68246 800
rect 69386 0 69442 800
rect 70490 0 70546 800
rect 71686 0 71742 800
rect 72882 0 72938 800
rect 73986 0 74042 800
rect 75182 0 75238 800
rect 76378 0 76434 800
rect 77482 0 77538 800
rect 78678 0 78734 800
rect 79874 0 79930 800
rect 81070 0 81126 800
rect 82174 0 82230 800
rect 83370 0 83426 800
rect 84566 0 84622 800
rect 85670 0 85726 800
rect 86866 0 86922 800
rect 88062 0 88118 800
rect 89166 0 89222 800
rect 90362 0 90418 800
rect 91558 0 91614 800
rect 92662 0 92718 800
rect 93858 0 93914 800
rect 95054 0 95110 800
rect 96158 0 96214 800
rect 97354 0 97410 800
rect 98550 0 98606 800
rect 99654 0 99710 800
rect 100850 0 100906 800
rect 102046 0 102102 800
rect 103150 0 103206 800
rect 104346 0 104402 800
rect 105542 0 105598 800
rect 106738 0 106794 800
rect 107842 0 107898 800
rect 109038 0 109094 800
rect 110234 0 110290 800
rect 111338 0 111394 800
rect 112534 0 112590 800
rect 113730 0 113786 800
rect 114834 0 114890 800
rect 116030 0 116086 800
rect 117226 0 117282 800
rect 118330 0 118386 800
rect 119526 0 119582 800
rect 120722 0 120778 800
rect 121826 0 121882 800
rect 123022 0 123078 800
rect 124218 0 124274 800
rect 125322 0 125378 800
rect 126518 0 126574 800
rect 127714 0 127770 800
rect 128818 0 128874 800
rect 130014 0 130070 800
rect 131210 0 131266 800
rect 132406 0 132462 800
rect 133510 0 133566 800
rect 134706 0 134762 800
rect 135902 0 135958 800
rect 137006 0 137062 800
rect 138202 0 138258 800
rect 139398 0 139454 800
rect 140502 0 140558 800
rect 141698 0 141754 800
rect 142894 0 142950 800
rect 143998 0 144054 800
rect 145194 0 145250 800
rect 146390 0 146446 800
rect 147494 0 147550 800
rect 148690 0 148746 800
rect 149886 0 149942 800
rect 150990 0 151046 800
rect 152186 0 152242 800
rect 153382 0 153438 800
rect 154486 0 154542 800
rect 155682 0 155738 800
rect 156878 0 156934 800
rect 158074 0 158130 800
rect 159178 0 159234 800
rect 160374 0 160430 800
rect 161570 0 161626 800
rect 162674 0 162730 800
rect 163870 0 163926 800
rect 165066 0 165122 800
rect 166170 0 166226 800
rect 167366 0 167422 800
rect 168562 0 168618 800
rect 169666 0 169722 800
rect 170862 0 170918 800
rect 172058 0 172114 800
rect 173162 0 173218 800
rect 174358 0 174414 800
rect 175554 0 175610 800
rect 176658 0 176714 800
rect 177854 0 177910 800
rect 179050 0 179106 800
rect 180154 0 180210 800
rect 181350 0 181406 800
rect 182546 0 182602 800
rect 183742 0 183798 800
rect 184846 0 184902 800
rect 186042 0 186098 800
rect 187238 0 187294 800
rect 188342 0 188398 800
rect 189538 0 189594 800
rect 190734 0 190790 800
rect 191838 0 191894 800
rect 193034 0 193090 800
rect 194230 0 194286 800
rect 195334 0 195390 800
rect 196530 0 196586 800
rect 197726 0 197782 800
rect 198830 0 198886 800
rect 200026 0 200082 800
rect 201222 0 201278 800
rect 202326 0 202382 800
rect 203522 0 203578 800
rect 204718 0 204774 800
rect 205822 0 205878 800
rect 207018 0 207074 800
rect 208214 0 208270 800
rect 209318 0 209374 800
rect 210514 0 210570 800
rect 211710 0 211766 800
rect 212906 0 212962 800
rect 214010 0 214066 800
rect 215206 0 215262 800
rect 216402 0 216458 800
rect 217506 0 217562 800
rect 218702 0 218758 800
rect 219898 0 219954 800
rect 221002 0 221058 800
rect 222198 0 222254 800
rect 223394 0 223450 800
rect 224498 0 224554 800
rect 225694 0 225750 800
rect 226890 0 226946 800
rect 227994 0 228050 800
rect 229190 0 229246 800
rect 230386 0 230442 800
rect 231490 0 231546 800
rect 232686 0 232742 800
rect 233882 0 233938 800
rect 234986 0 235042 800
rect 236182 0 236238 800
rect 237378 0 237434 800
rect 238574 0 238630 800
rect 239678 0 239734 800
rect 240874 0 240930 800
rect 242070 0 242126 800
rect 243174 0 243230 800
rect 244370 0 244426 800
rect 245566 0 245622 800
rect 246670 0 246726 800
rect 247866 0 247922 800
rect 249062 0 249118 800
rect 250166 0 250222 800
rect 251362 0 251418 800
rect 252558 0 252614 800
rect 253662 0 253718 800
rect 254858 0 254914 800
rect 256054 0 256110 800
rect 257158 0 257214 800
rect 258354 0 258410 800
rect 259550 0 259606 800
rect 260654 0 260710 800
rect 261850 0 261906 800
rect 263046 0 263102 800
rect 264242 0 264298 800
rect 265346 0 265402 800
rect 266542 0 266598 800
rect 267738 0 267794 800
rect 268842 0 268898 800
rect 270038 0 270094 800
rect 271234 0 271290 800
rect 272338 0 272394 800
rect 273534 0 273590 800
rect 274730 0 274786 800
rect 275834 0 275890 800
rect 277030 0 277086 800
rect 278226 0 278282 800
rect 279330 0 279386 800
rect 280526 0 280582 800
rect 281722 0 281778 800
rect 282826 0 282882 800
rect 284022 0 284078 800
rect 285218 0 285274 800
rect 286322 0 286378 800
rect 287518 0 287574 800
rect 288714 0 288770 800
rect 289910 0 289966 800
rect 291014 0 291070 800
rect 292210 0 292266 800
rect 293406 0 293462 800
rect 294510 0 294566 800
rect 295706 0 295762 800
rect 296902 0 296958 800
rect 298006 0 298062 800
rect 299202 0 299258 800
rect 300398 0 300454 800
rect 301502 0 301558 800
rect 302698 0 302754 800
rect 303894 0 303950 800
rect 304998 0 305054 800
rect 306194 0 306250 800
rect 307390 0 307446 800
rect 308494 0 308550 800
rect 309690 0 309746 800
rect 310886 0 310942 800
rect 311990 0 312046 800
rect 313186 0 313242 800
rect 314382 0 314438 800
rect 315578 0 315634 800
rect 316682 0 316738 800
rect 317878 0 317934 800
rect 319074 0 319130 800
rect 320178 0 320234 800
rect 321374 0 321430 800
rect 322570 0 322626 800
rect 323674 0 323730 800
rect 324870 0 324926 800
rect 326066 0 326122 800
rect 327170 0 327226 800
rect 328366 0 328422 800
rect 329562 0 329618 800
rect 330666 0 330722 800
rect 331862 0 331918 800
rect 333058 0 333114 800
rect 334162 0 334218 800
rect 335358 0 335414 800
rect 336554 0 336610 800
rect 337658 0 337714 800
rect 338854 0 338910 800
rect 340050 0 340106 800
rect 341246 0 341302 800
rect 342350 0 342406 800
rect 343546 0 343602 800
rect 344742 0 344798 800
rect 345846 0 345902 800
rect 347042 0 347098 800
rect 348238 0 348294 800
rect 349342 0 349398 800
rect 350538 0 350594 800
rect 351734 0 351790 800
rect 352838 0 352894 800
rect 354034 0 354090 800
rect 355230 0 355286 800
rect 356334 0 356390 800
rect 357530 0 357586 800
rect 358726 0 358782 800
rect 359830 0 359886 800
rect 361026 0 361082 800
rect 362222 0 362278 800
rect 363326 0 363382 800
rect 364522 0 364578 800
rect 365718 0 365774 800
rect 366914 0 366970 800
rect 368018 0 368074 800
rect 369214 0 369270 800
rect 370410 0 370466 800
rect 371514 0 371570 800
rect 372710 0 372766 800
rect 373906 0 373962 800
rect 375010 0 375066 800
rect 376206 0 376262 800
rect 377402 0 377458 800
rect 378506 0 378562 800
rect 379702 0 379758 800
rect 380898 0 380954 800
rect 382002 0 382058 800
rect 383198 0 383254 800
rect 384394 0 384450 800
rect 385498 0 385554 800
rect 386694 0 386750 800
rect 387890 0 387946 800
rect 388994 0 389050 800
rect 390190 0 390246 800
rect 391386 0 391442 800
rect 392490 0 392546 800
rect 393686 0 393742 800
rect 394882 0 394938 800
rect 396078 0 396134 800
rect 397182 0 397238 800
rect 398378 0 398434 800
rect 399574 0 399630 800
rect 400678 0 400734 800
rect 401874 0 401930 800
rect 403070 0 403126 800
rect 404174 0 404230 800
rect 405370 0 405426 800
rect 406566 0 406622 800
rect 407670 0 407726 800
rect 408866 0 408922 800
rect 410062 0 410118 800
rect 411166 0 411222 800
rect 412362 0 412418 800
rect 413558 0 413614 800
rect 414662 0 414718 800
rect 415858 0 415914 800
rect 417054 0 417110 800
rect 418158 0 418214 800
rect 419354 0 419410 800
rect 420550 0 420606 800
rect 421746 0 421802 800
rect 422850 0 422906 800
rect 424046 0 424102 800
rect 425242 0 425298 800
rect 426346 0 426402 800
rect 427542 0 427598 800
rect 428738 0 428794 800
rect 429842 0 429898 800
rect 431038 0 431094 800
rect 432234 0 432290 800
rect 433338 0 433394 800
rect 434534 0 434590 800
rect 435730 0 435786 800
rect 436834 0 436890 800
rect 438030 0 438086 800
rect 439226 0 439282 800
rect 440330 0 440386 800
rect 441526 0 441582 800
rect 442722 0 442778 800
rect 443826 0 443882 800
rect 445022 0 445078 800
rect 446218 0 446274 800
rect 447414 0 447470 800
rect 448518 0 448574 800
rect 449714 0 449770 800
rect 450910 0 450966 800
rect 452014 0 452070 800
rect 453210 0 453266 800
rect 454406 0 454462 800
rect 455510 0 455566 800
rect 456706 0 456762 800
rect 457902 0 457958 800
rect 459006 0 459062 800
rect 460202 0 460258 800
rect 461398 0 461454 800
rect 462502 0 462558 800
rect 463698 0 463754 800
rect 464894 0 464950 800
rect 465998 0 466054 800
rect 467194 0 467250 800
rect 468390 0 468446 800
rect 469494 0 469550 800
rect 470690 0 470746 800
rect 471886 0 471942 800
rect 473082 0 473138 800
rect 474186 0 474242 800
rect 475382 0 475438 800
rect 476578 0 476634 800
rect 477682 0 477738 800
rect 478878 0 478934 800
rect 480074 0 480130 800
rect 481178 0 481234 800
rect 482374 0 482430 800
rect 483570 0 483626 800
rect 484674 0 484730 800
rect 485870 0 485926 800
rect 487066 0 487122 800
rect 488170 0 488226 800
rect 489366 0 489422 800
rect 490562 0 490618 800
rect 491666 0 491722 800
rect 492862 0 492918 800
rect 494058 0 494114 800
rect 495162 0 495218 800
rect 496358 0 496414 800
rect 497554 0 497610 800
rect 498750 0 498806 800
rect 499854 0 499910 800
rect 501050 0 501106 800
rect 502246 0 502302 800
rect 503350 0 503406 800
rect 504546 0 504602 800
rect 505742 0 505798 800
rect 506846 0 506902 800
rect 508042 0 508098 800
rect 509238 0 509294 800
rect 510342 0 510398 800
rect 511538 0 511594 800
rect 512734 0 512790 800
rect 513838 0 513894 800
rect 515034 0 515090 800
rect 516230 0 516286 800
rect 517334 0 517390 800
rect 518530 0 518586 800
rect 519726 0 519782 800
rect 520830 0 520886 800
rect 522026 0 522082 800
rect 523222 0 523278 800
rect 524418 0 524474 800
rect 525522 0 525578 800
rect 526718 0 526774 800
rect 527914 0 527970 800
rect 529018 0 529074 800
rect 530214 0 530270 800
rect 531410 0 531466 800
rect 532514 0 532570 800
rect 533710 0 533766 800
rect 534906 0 534962 800
rect 536010 0 536066 800
rect 537206 0 537262 800
rect 538402 0 538458 800
rect 539506 0 539562 800
rect 540702 0 540758 800
rect 541898 0 541954 800
rect 543002 0 543058 800
rect 544198 0 544254 800
rect 545394 0 545450 800
rect 546498 0 546554 800
rect 547694 0 547750 800
rect 548890 0 548946 800
rect 550086 0 550142 800
rect 551190 0 551246 800
rect 552386 0 552442 800
rect 553582 0 553638 800
rect 554686 0 554742 800
rect 555882 0 555938 800
rect 557078 0 557134 800
rect 558182 0 558238 800
rect 559378 0 559434 800
rect 560574 0 560630 800
rect 561678 0 561734 800
rect 562874 0 562930 800
rect 564070 0 564126 800
rect 565174 0 565230 800
rect 566370 0 566426 800
rect 567566 0 567622 800
rect 568670 0 568726 800
rect 569866 0 569922 800
rect 571062 0 571118 800
rect 572166 0 572222 800
rect 573362 0 573418 800
rect 574558 0 574614 800
<< obsm2 >>
rect 572 694344 2446 694498
rect 2614 694344 7414 694498
rect 7582 694344 12474 694498
rect 12642 694344 17534 694498
rect 17702 694344 22594 694498
rect 22762 694344 27654 694498
rect 27822 694344 32714 694498
rect 32882 694344 37682 694498
rect 37850 694344 42742 694498
rect 42910 694344 47802 694498
rect 47970 694344 52862 694498
rect 53030 694344 57922 694498
rect 58090 694344 62982 694498
rect 63150 694344 67950 694498
rect 68118 694344 73010 694498
rect 73178 694344 78070 694498
rect 78238 694344 83130 694498
rect 83298 694344 88190 694498
rect 88358 694344 93250 694498
rect 93418 694344 98310 694498
rect 98478 694344 103278 694498
rect 103446 694344 108338 694498
rect 108506 694344 113398 694498
rect 113566 694344 118458 694498
rect 118626 694344 123518 694498
rect 123686 694344 128578 694498
rect 128746 694344 133546 694498
rect 133714 694344 138606 694498
rect 138774 694344 143666 694498
rect 143834 694344 148726 694498
rect 148894 694344 153786 694498
rect 153954 694344 158846 694498
rect 159014 694344 163814 694498
rect 163982 694344 168874 694498
rect 169042 694344 173934 694498
rect 174102 694344 178994 694498
rect 179162 694344 184054 694498
rect 184222 694344 189114 694498
rect 189282 694344 194174 694498
rect 194342 694344 199142 694498
rect 199310 694344 204202 694498
rect 204370 694344 209262 694498
rect 209430 694344 214322 694498
rect 214490 694344 219382 694498
rect 219550 694344 224442 694498
rect 224610 694344 229410 694498
rect 229578 694344 234470 694498
rect 234638 694344 239530 694498
rect 239698 694344 244590 694498
rect 244758 694344 249650 694498
rect 249818 694344 254710 694498
rect 254878 694344 259678 694498
rect 259846 694344 264738 694498
rect 264906 694344 269798 694498
rect 269966 694344 274858 694498
rect 275026 694344 279918 694498
rect 280086 694344 284978 694498
rect 285146 694344 290038 694498
rect 290206 694344 295006 694498
rect 295174 694344 300066 694498
rect 300234 694344 305126 694498
rect 305294 694344 310186 694498
rect 310354 694344 315246 694498
rect 315414 694344 320306 694498
rect 320474 694344 325274 694498
rect 325442 694344 330334 694498
rect 330502 694344 335394 694498
rect 335562 694344 340454 694498
rect 340622 694344 345514 694498
rect 345682 694344 350574 694498
rect 350742 694344 355542 694498
rect 355710 694344 360602 694498
rect 360770 694344 365662 694498
rect 365830 694344 370722 694498
rect 370890 694344 375782 694498
rect 375950 694344 380842 694498
rect 381010 694344 385902 694498
rect 386070 694344 390870 694498
rect 391038 694344 395930 694498
rect 396098 694344 400990 694498
rect 401158 694344 406050 694498
rect 406218 694344 411110 694498
rect 411278 694344 416170 694498
rect 416338 694344 421138 694498
rect 421306 694344 426198 694498
rect 426366 694344 431258 694498
rect 431426 694344 436318 694498
rect 436486 694344 441378 694498
rect 441546 694344 446438 694498
rect 446606 694344 451406 694498
rect 451574 694344 456466 694498
rect 456634 694344 461526 694498
rect 461694 694344 466586 694498
rect 466754 694344 471646 694498
rect 471814 694344 476706 694498
rect 476874 694344 481766 694498
rect 481934 694344 486734 694498
rect 486902 694344 491794 694498
rect 491962 694344 496854 694498
rect 497022 694344 501914 694498
rect 502082 694344 506974 694498
rect 507142 694344 512034 694498
rect 512202 694344 517002 694498
rect 517170 694344 522062 694498
rect 522230 694344 527122 694498
rect 527290 694344 532182 694498
rect 532350 694344 537242 694498
rect 537410 694344 542302 694498
rect 542470 694344 547270 694498
rect 547438 694344 552330 694498
rect 552498 694344 557390 694498
rect 557558 694344 562450 694498
rect 562618 694344 567510 694498
rect 567678 694344 572570 694498
rect 572738 694344 574612 694498
rect 572 856 574612 694344
rect 682 2 1618 856
rect 1786 2 2814 856
rect 2982 2 4010 856
rect 4178 2 5114 856
rect 5282 2 6310 856
rect 6478 2 7506 856
rect 7674 2 8610 856
rect 8778 2 9806 856
rect 9974 2 11002 856
rect 11170 2 12106 856
rect 12274 2 13302 856
rect 13470 2 14498 856
rect 14666 2 15602 856
rect 15770 2 16798 856
rect 16966 2 17994 856
rect 18162 2 19098 856
rect 19266 2 20294 856
rect 20462 2 21490 856
rect 21658 2 22594 856
rect 22762 2 23790 856
rect 23958 2 24986 856
rect 25154 2 26090 856
rect 26258 2 27286 856
rect 27454 2 28482 856
rect 28650 2 29678 856
rect 29846 2 30782 856
rect 30950 2 31978 856
rect 32146 2 33174 856
rect 33342 2 34278 856
rect 34446 2 35474 856
rect 35642 2 36670 856
rect 36838 2 37774 856
rect 37942 2 38970 856
rect 39138 2 40166 856
rect 40334 2 41270 856
rect 41438 2 42466 856
rect 42634 2 43662 856
rect 43830 2 44766 856
rect 44934 2 45962 856
rect 46130 2 47158 856
rect 47326 2 48262 856
rect 48430 2 49458 856
rect 49626 2 50654 856
rect 50822 2 51758 856
rect 51926 2 52954 856
rect 53122 2 54150 856
rect 54318 2 55346 856
rect 55514 2 56450 856
rect 56618 2 57646 856
rect 57814 2 58842 856
rect 59010 2 59946 856
rect 60114 2 61142 856
rect 61310 2 62338 856
rect 62506 2 63442 856
rect 63610 2 64638 856
rect 64806 2 65834 856
rect 66002 2 66938 856
rect 67106 2 68134 856
rect 68302 2 69330 856
rect 69498 2 70434 856
rect 70602 2 71630 856
rect 71798 2 72826 856
rect 72994 2 73930 856
rect 74098 2 75126 856
rect 75294 2 76322 856
rect 76490 2 77426 856
rect 77594 2 78622 856
rect 78790 2 79818 856
rect 79986 2 81014 856
rect 81182 2 82118 856
rect 82286 2 83314 856
rect 83482 2 84510 856
rect 84678 2 85614 856
rect 85782 2 86810 856
rect 86978 2 88006 856
rect 88174 2 89110 856
rect 89278 2 90306 856
rect 90474 2 91502 856
rect 91670 2 92606 856
rect 92774 2 93802 856
rect 93970 2 94998 856
rect 95166 2 96102 856
rect 96270 2 97298 856
rect 97466 2 98494 856
rect 98662 2 99598 856
rect 99766 2 100794 856
rect 100962 2 101990 856
rect 102158 2 103094 856
rect 103262 2 104290 856
rect 104458 2 105486 856
rect 105654 2 106682 856
rect 106850 2 107786 856
rect 107954 2 108982 856
rect 109150 2 110178 856
rect 110346 2 111282 856
rect 111450 2 112478 856
rect 112646 2 113674 856
rect 113842 2 114778 856
rect 114946 2 115974 856
rect 116142 2 117170 856
rect 117338 2 118274 856
rect 118442 2 119470 856
rect 119638 2 120666 856
rect 120834 2 121770 856
rect 121938 2 122966 856
rect 123134 2 124162 856
rect 124330 2 125266 856
rect 125434 2 126462 856
rect 126630 2 127658 856
rect 127826 2 128762 856
rect 128930 2 129958 856
rect 130126 2 131154 856
rect 131322 2 132350 856
rect 132518 2 133454 856
rect 133622 2 134650 856
rect 134818 2 135846 856
rect 136014 2 136950 856
rect 137118 2 138146 856
rect 138314 2 139342 856
rect 139510 2 140446 856
rect 140614 2 141642 856
rect 141810 2 142838 856
rect 143006 2 143942 856
rect 144110 2 145138 856
rect 145306 2 146334 856
rect 146502 2 147438 856
rect 147606 2 148634 856
rect 148802 2 149830 856
rect 149998 2 150934 856
rect 151102 2 152130 856
rect 152298 2 153326 856
rect 153494 2 154430 856
rect 154598 2 155626 856
rect 155794 2 156822 856
rect 156990 2 158018 856
rect 158186 2 159122 856
rect 159290 2 160318 856
rect 160486 2 161514 856
rect 161682 2 162618 856
rect 162786 2 163814 856
rect 163982 2 165010 856
rect 165178 2 166114 856
rect 166282 2 167310 856
rect 167478 2 168506 856
rect 168674 2 169610 856
rect 169778 2 170806 856
rect 170974 2 172002 856
rect 172170 2 173106 856
rect 173274 2 174302 856
rect 174470 2 175498 856
rect 175666 2 176602 856
rect 176770 2 177798 856
rect 177966 2 178994 856
rect 179162 2 180098 856
rect 180266 2 181294 856
rect 181462 2 182490 856
rect 182658 2 183686 856
rect 183854 2 184790 856
rect 184958 2 185986 856
rect 186154 2 187182 856
rect 187350 2 188286 856
rect 188454 2 189482 856
rect 189650 2 190678 856
rect 190846 2 191782 856
rect 191950 2 192978 856
rect 193146 2 194174 856
rect 194342 2 195278 856
rect 195446 2 196474 856
rect 196642 2 197670 856
rect 197838 2 198774 856
rect 198942 2 199970 856
rect 200138 2 201166 856
rect 201334 2 202270 856
rect 202438 2 203466 856
rect 203634 2 204662 856
rect 204830 2 205766 856
rect 205934 2 206962 856
rect 207130 2 208158 856
rect 208326 2 209262 856
rect 209430 2 210458 856
rect 210626 2 211654 856
rect 211822 2 212850 856
rect 213018 2 213954 856
rect 214122 2 215150 856
rect 215318 2 216346 856
rect 216514 2 217450 856
rect 217618 2 218646 856
rect 218814 2 219842 856
rect 220010 2 220946 856
rect 221114 2 222142 856
rect 222310 2 223338 856
rect 223506 2 224442 856
rect 224610 2 225638 856
rect 225806 2 226834 856
rect 227002 2 227938 856
rect 228106 2 229134 856
rect 229302 2 230330 856
rect 230498 2 231434 856
rect 231602 2 232630 856
rect 232798 2 233826 856
rect 233994 2 234930 856
rect 235098 2 236126 856
rect 236294 2 237322 856
rect 237490 2 238518 856
rect 238686 2 239622 856
rect 239790 2 240818 856
rect 240986 2 242014 856
rect 242182 2 243118 856
rect 243286 2 244314 856
rect 244482 2 245510 856
rect 245678 2 246614 856
rect 246782 2 247810 856
rect 247978 2 249006 856
rect 249174 2 250110 856
rect 250278 2 251306 856
rect 251474 2 252502 856
rect 252670 2 253606 856
rect 253774 2 254802 856
rect 254970 2 255998 856
rect 256166 2 257102 856
rect 257270 2 258298 856
rect 258466 2 259494 856
rect 259662 2 260598 856
rect 260766 2 261794 856
rect 261962 2 262990 856
rect 263158 2 264186 856
rect 264354 2 265290 856
rect 265458 2 266486 856
rect 266654 2 267682 856
rect 267850 2 268786 856
rect 268954 2 269982 856
rect 270150 2 271178 856
rect 271346 2 272282 856
rect 272450 2 273478 856
rect 273646 2 274674 856
rect 274842 2 275778 856
rect 275946 2 276974 856
rect 277142 2 278170 856
rect 278338 2 279274 856
rect 279442 2 280470 856
rect 280638 2 281666 856
rect 281834 2 282770 856
rect 282938 2 283966 856
rect 284134 2 285162 856
rect 285330 2 286266 856
rect 286434 2 287462 856
rect 287630 2 288658 856
rect 288826 2 289854 856
rect 290022 2 290958 856
rect 291126 2 292154 856
rect 292322 2 293350 856
rect 293518 2 294454 856
rect 294622 2 295650 856
rect 295818 2 296846 856
rect 297014 2 297950 856
rect 298118 2 299146 856
rect 299314 2 300342 856
rect 300510 2 301446 856
rect 301614 2 302642 856
rect 302810 2 303838 856
rect 304006 2 304942 856
rect 305110 2 306138 856
rect 306306 2 307334 856
rect 307502 2 308438 856
rect 308606 2 309634 856
rect 309802 2 310830 856
rect 310998 2 311934 856
rect 312102 2 313130 856
rect 313298 2 314326 856
rect 314494 2 315522 856
rect 315690 2 316626 856
rect 316794 2 317822 856
rect 317990 2 319018 856
rect 319186 2 320122 856
rect 320290 2 321318 856
rect 321486 2 322514 856
rect 322682 2 323618 856
rect 323786 2 324814 856
rect 324982 2 326010 856
rect 326178 2 327114 856
rect 327282 2 328310 856
rect 328478 2 329506 856
rect 329674 2 330610 856
rect 330778 2 331806 856
rect 331974 2 333002 856
rect 333170 2 334106 856
rect 334274 2 335302 856
rect 335470 2 336498 856
rect 336666 2 337602 856
rect 337770 2 338798 856
rect 338966 2 339994 856
rect 340162 2 341190 856
rect 341358 2 342294 856
rect 342462 2 343490 856
rect 343658 2 344686 856
rect 344854 2 345790 856
rect 345958 2 346986 856
rect 347154 2 348182 856
rect 348350 2 349286 856
rect 349454 2 350482 856
rect 350650 2 351678 856
rect 351846 2 352782 856
rect 352950 2 353978 856
rect 354146 2 355174 856
rect 355342 2 356278 856
rect 356446 2 357474 856
rect 357642 2 358670 856
rect 358838 2 359774 856
rect 359942 2 360970 856
rect 361138 2 362166 856
rect 362334 2 363270 856
rect 363438 2 364466 856
rect 364634 2 365662 856
rect 365830 2 366858 856
rect 367026 2 367962 856
rect 368130 2 369158 856
rect 369326 2 370354 856
rect 370522 2 371458 856
rect 371626 2 372654 856
rect 372822 2 373850 856
rect 374018 2 374954 856
rect 375122 2 376150 856
rect 376318 2 377346 856
rect 377514 2 378450 856
rect 378618 2 379646 856
rect 379814 2 380842 856
rect 381010 2 381946 856
rect 382114 2 383142 856
rect 383310 2 384338 856
rect 384506 2 385442 856
rect 385610 2 386638 856
rect 386806 2 387834 856
rect 388002 2 388938 856
rect 389106 2 390134 856
rect 390302 2 391330 856
rect 391498 2 392434 856
rect 392602 2 393630 856
rect 393798 2 394826 856
rect 394994 2 396022 856
rect 396190 2 397126 856
rect 397294 2 398322 856
rect 398490 2 399518 856
rect 399686 2 400622 856
rect 400790 2 401818 856
rect 401986 2 403014 856
rect 403182 2 404118 856
rect 404286 2 405314 856
rect 405482 2 406510 856
rect 406678 2 407614 856
rect 407782 2 408810 856
rect 408978 2 410006 856
rect 410174 2 411110 856
rect 411278 2 412306 856
rect 412474 2 413502 856
rect 413670 2 414606 856
rect 414774 2 415802 856
rect 415970 2 416998 856
rect 417166 2 418102 856
rect 418270 2 419298 856
rect 419466 2 420494 856
rect 420662 2 421690 856
rect 421858 2 422794 856
rect 422962 2 423990 856
rect 424158 2 425186 856
rect 425354 2 426290 856
rect 426458 2 427486 856
rect 427654 2 428682 856
rect 428850 2 429786 856
rect 429954 2 430982 856
rect 431150 2 432178 856
rect 432346 2 433282 856
rect 433450 2 434478 856
rect 434646 2 435674 856
rect 435842 2 436778 856
rect 436946 2 437974 856
rect 438142 2 439170 856
rect 439338 2 440274 856
rect 440442 2 441470 856
rect 441638 2 442666 856
rect 442834 2 443770 856
rect 443938 2 444966 856
rect 445134 2 446162 856
rect 446330 2 447358 856
rect 447526 2 448462 856
rect 448630 2 449658 856
rect 449826 2 450854 856
rect 451022 2 451958 856
rect 452126 2 453154 856
rect 453322 2 454350 856
rect 454518 2 455454 856
rect 455622 2 456650 856
rect 456818 2 457846 856
rect 458014 2 458950 856
rect 459118 2 460146 856
rect 460314 2 461342 856
rect 461510 2 462446 856
rect 462614 2 463642 856
rect 463810 2 464838 856
rect 465006 2 465942 856
rect 466110 2 467138 856
rect 467306 2 468334 856
rect 468502 2 469438 856
rect 469606 2 470634 856
rect 470802 2 471830 856
rect 471998 2 473026 856
rect 473194 2 474130 856
rect 474298 2 475326 856
rect 475494 2 476522 856
rect 476690 2 477626 856
rect 477794 2 478822 856
rect 478990 2 480018 856
rect 480186 2 481122 856
rect 481290 2 482318 856
rect 482486 2 483514 856
rect 483682 2 484618 856
rect 484786 2 485814 856
rect 485982 2 487010 856
rect 487178 2 488114 856
rect 488282 2 489310 856
rect 489478 2 490506 856
rect 490674 2 491610 856
rect 491778 2 492806 856
rect 492974 2 494002 856
rect 494170 2 495106 856
rect 495274 2 496302 856
rect 496470 2 497498 856
rect 497666 2 498694 856
rect 498862 2 499798 856
rect 499966 2 500994 856
rect 501162 2 502190 856
rect 502358 2 503294 856
rect 503462 2 504490 856
rect 504658 2 505686 856
rect 505854 2 506790 856
rect 506958 2 507986 856
rect 508154 2 509182 856
rect 509350 2 510286 856
rect 510454 2 511482 856
rect 511650 2 512678 856
rect 512846 2 513782 856
rect 513950 2 514978 856
rect 515146 2 516174 856
rect 516342 2 517278 856
rect 517446 2 518474 856
rect 518642 2 519670 856
rect 519838 2 520774 856
rect 520942 2 521970 856
rect 522138 2 523166 856
rect 523334 2 524362 856
rect 524530 2 525466 856
rect 525634 2 526662 856
rect 526830 2 527858 856
rect 528026 2 528962 856
rect 529130 2 530158 856
rect 530326 2 531354 856
rect 531522 2 532458 856
rect 532626 2 533654 856
rect 533822 2 534850 856
rect 535018 2 535954 856
rect 536122 2 537150 856
rect 537318 2 538346 856
rect 538514 2 539450 856
rect 539618 2 540646 856
rect 540814 2 541842 856
rect 542010 2 542946 856
rect 543114 2 544142 856
rect 544310 2 545338 856
rect 545506 2 546442 856
rect 546610 2 547638 856
rect 547806 2 548834 856
rect 549002 2 550030 856
rect 550198 2 551134 856
rect 551302 2 552330 856
rect 552498 2 553526 856
rect 553694 2 554630 856
rect 554798 2 555826 856
rect 555994 2 557022 856
rect 557190 2 558126 856
rect 558294 2 559322 856
rect 559490 2 560518 856
rect 560686 2 561622 856
rect 561790 2 562818 856
rect 562986 2 564014 856
rect 564182 2 565118 856
rect 565286 2 566314 856
rect 566482 2 567510 856
rect 567678 2 568614 856
rect 568782 2 569810 856
rect 569978 2 571006 856
rect 571174 2 572110 856
rect 572278 2 573306 856
rect 573474 2 574502 856
<< obsm3 >>
rect 2865 35 573699 692545
<< metal4 >>
rect 4208 2128 4528 692560
rect 19568 2128 19888 692560
rect 34928 2128 35248 692560
rect 50288 2128 50608 692560
rect 65648 2128 65968 692560
rect 81008 2128 81328 692560
rect 96368 2128 96688 692560
rect 111728 2128 112048 692560
rect 127088 2128 127408 692560
rect 142448 2128 142768 692560
rect 157808 2128 158128 692560
rect 173168 2128 173488 692560
rect 188528 2128 188848 692560
rect 203888 2128 204208 692560
rect 219248 2128 219568 692560
rect 234608 2128 234928 692560
rect 249968 2128 250288 692560
rect 265328 2128 265648 692560
rect 280688 2128 281008 692560
rect 296048 2128 296368 692560
rect 311408 2128 311728 692560
rect 326768 2128 327088 692560
rect 342128 2128 342448 692560
rect 357488 2128 357808 692560
rect 372848 2128 373168 692560
rect 388208 2128 388528 692560
rect 403568 2128 403888 692560
rect 418928 2128 419248 692560
rect 434288 2128 434608 692560
rect 449648 2128 449968 692560
rect 465008 2128 465328 692560
rect 480368 2128 480688 692560
rect 495728 2128 496048 692560
rect 511088 2128 511408 692560
rect 526448 2128 526768 692560
rect 541808 2128 542128 692560
rect 557168 2128 557488 692560
rect 572528 2128 572848 692560
<< obsm4 >>
rect 9811 2483 19488 692069
rect 19968 2483 34848 692069
rect 35328 2483 50208 692069
rect 50688 2483 65568 692069
rect 66048 2483 80928 692069
rect 81408 2483 96288 692069
rect 96768 2483 111648 692069
rect 112128 2483 127008 692069
rect 127488 2483 142368 692069
rect 142848 2483 157728 692069
rect 158208 2483 173088 692069
rect 173568 2483 188448 692069
rect 188928 2483 203808 692069
rect 204288 2483 219168 692069
rect 219648 2483 234528 692069
rect 235008 2483 249888 692069
rect 250368 2483 265248 692069
rect 265728 2483 280608 692069
rect 281088 2483 295968 692069
rect 296448 2483 311328 692069
rect 311808 2483 326688 692069
rect 327168 2483 342048 692069
rect 342528 2483 357408 692069
rect 357888 2483 372768 692069
rect 373248 2483 388128 692069
rect 388608 2483 403488 692069
rect 403968 2483 418848 692069
rect 419328 2483 434208 692069
rect 434688 2483 449568 692069
rect 450048 2483 464928 692069
rect 465408 2483 480288 692069
rect 480768 2483 495648 692069
rect 496128 2483 511008 692069
rect 511488 2483 526368 692069
rect 526848 2483 541728 692069
rect 542208 2483 557088 692069
rect 557568 2483 572365 692069
<< labels >>
rlabel metal2 s 2502 694400 2558 695200 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 153842 694400 153898 695200 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 168930 694400 168986 695200 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 184110 694400 184166 695200 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 199198 694400 199254 695200 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 214378 694400 214434 695200 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 229466 694400 229522 695200 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 244646 694400 244702 695200 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 259734 694400 259790 695200 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 274914 694400 274970 695200 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 290094 694400 290150 695200 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 17590 694400 17646 695200 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 305182 694400 305238 695200 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 320362 694400 320418 695200 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 335450 694400 335506 695200 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 350630 694400 350686 695200 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 365718 694400 365774 695200 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 380898 694400 380954 695200 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 395986 694400 396042 695200 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 411166 694400 411222 695200 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 426254 694400 426310 695200 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 441434 694400 441490 695200 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 32770 694400 32826 695200 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 456522 694400 456578 695200 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 471702 694400 471758 695200 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 486790 694400 486846 695200 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 501970 694400 502026 695200 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 517058 694400 517114 695200 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 532238 694400 532294 695200 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 547326 694400 547382 695200 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 562506 694400 562562 695200 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 47858 694400 47914 695200 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 63038 694400 63094 695200 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 78126 694400 78182 695200 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 93306 694400 93362 695200 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 108394 694400 108450 695200 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 123574 694400 123630 695200 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 138662 694400 138718 695200 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 7470 694400 7526 695200 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 158902 694400 158958 695200 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 173990 694400 174046 695200 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 189170 694400 189226 695200 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 204258 694400 204314 695200 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 219438 694400 219494 695200 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 234526 694400 234582 695200 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 249706 694400 249762 695200 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 264794 694400 264850 695200 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 279974 694400 280030 695200 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 295062 694400 295118 695200 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 22650 694400 22706 695200 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 310242 694400 310298 695200 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 325330 694400 325386 695200 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 340510 694400 340566 695200 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 355598 694400 355654 695200 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 370778 694400 370834 695200 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 385958 694400 386014 695200 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 401046 694400 401102 695200 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 416226 694400 416282 695200 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 431314 694400 431370 695200 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 446494 694400 446550 695200 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 37738 694400 37794 695200 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 461582 694400 461638 695200 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 476762 694400 476818 695200 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 491850 694400 491906 695200 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 507030 694400 507086 695200 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 522118 694400 522174 695200 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 537298 694400 537354 695200 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 552386 694400 552442 695200 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 567566 694400 567622 695200 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 52918 694400 52974 695200 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 68006 694400 68062 695200 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 83186 694400 83242 695200 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 98366 694400 98422 695200 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 113454 694400 113510 695200 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 128634 694400 128690 695200 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 143722 694400 143778 695200 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 12530 694400 12586 695200 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 163870 694400 163926 695200 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 179050 694400 179106 695200 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 194230 694400 194286 695200 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 209318 694400 209374 695200 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 224498 694400 224554 695200 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 239586 694400 239642 695200 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 254766 694400 254822 695200 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 269854 694400 269910 695200 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 285034 694400 285090 695200 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 300122 694400 300178 695200 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 27710 694400 27766 695200 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 315302 694400 315358 695200 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 330390 694400 330446 695200 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 345570 694400 345626 695200 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 360658 694400 360714 695200 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 375838 694400 375894 695200 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 390926 694400 390982 695200 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 406106 694400 406162 695200 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 421194 694400 421250 695200 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 436374 694400 436430 695200 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 451462 694400 451518 695200 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 42798 694400 42854 695200 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 466642 694400 466698 695200 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 481822 694400 481878 695200 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 496910 694400 496966 695200 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 512090 694400 512146 695200 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 527178 694400 527234 695200 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 542358 694400 542414 695200 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 557446 694400 557502 695200 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 572626 694400 572682 695200 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 57978 694400 58034 695200 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 73066 694400 73122 695200 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 88246 694400 88302 695200 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 103334 694400 103390 695200 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 118514 694400 118570 695200 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 133602 694400 133658 695200 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 148782 694400 148838 695200 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 572166 0 572222 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 573362 0 573418 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 574558 0 574614 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 474186 0 474242 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 477682 0 477738 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 481178 0 481234 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 484674 0 484730 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 488170 0 488226 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 491666 0 491722 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 495162 0 495218 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 498750 0 498806 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 502246 0 502302 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 505742 0 505798 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 509238 0 509294 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 512734 0 512790 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 516230 0 516286 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 519726 0 519782 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 523222 0 523278 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 526718 0 526774 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 530214 0 530270 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 533710 0 533766 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 537206 0 537262 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 540702 0 540758 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 544198 0 544254 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 547694 0 547750 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 551190 0 551246 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 554686 0 554742 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 558182 0 558238 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 561678 0 561734 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 565174 0 565230 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 568670 0 568726 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 190734 0 190790 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 194230 0 194286 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 215206 0 215262 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 229190 0 229246 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 232686 0 232742 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 236182 0 236238 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 243174 0 243230 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 253662 0 253718 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 257158 0 257214 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 260654 0 260710 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 264242 0 264298 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 267738 0 267794 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 271234 0 271290 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 274730 0 274786 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 278226 0 278282 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 281722 0 281778 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 285218 0 285274 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 288714 0 288770 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 292210 0 292266 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 295706 0 295762 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 299202 0 299258 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 302698 0 302754 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 306194 0 306250 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 309690 0 309746 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 313186 0 313242 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 316682 0 316738 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 320178 0 320234 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 323674 0 323730 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 327170 0 327226 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 330666 0 330722 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 334162 0 334218 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 337658 0 337714 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 341246 0 341302 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 344742 0 344798 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 348238 0 348294 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 351734 0 351790 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 355230 0 355286 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 358726 0 358782 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 362222 0 362278 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 365718 0 365774 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 369214 0 369270 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 372710 0 372766 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 376206 0 376262 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 379702 0 379758 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 383198 0 383254 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 386694 0 386750 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 390190 0 390246 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 393686 0 393742 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 397182 0 397238 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 400678 0 400734 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 404174 0 404230 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 407670 0 407726 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 411166 0 411222 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 414662 0 414718 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 418158 0 418214 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 421746 0 421802 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 425242 0 425298 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 428738 0 428794 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 432234 0 432290 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 435730 0 435786 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 439226 0 439282 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 442722 0 442778 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 446218 0 446274 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 449714 0 449770 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 453210 0 453266 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 456706 0 456762 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 460202 0 460258 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 463698 0 463754 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 467194 0 467250 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 470690 0 470746 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 475382 0 475438 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 478878 0 478934 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 482374 0 482430 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 485870 0 485926 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 489366 0 489422 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 492862 0 492918 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 496358 0 496414 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 499854 0 499910 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 503350 0 503406 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 506846 0 506902 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 510342 0 510398 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 513838 0 513894 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 517334 0 517390 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 520830 0 520886 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 524418 0 524474 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 527914 0 527970 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 531410 0 531466 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 534906 0 534962 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 538402 0 538458 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 541898 0 541954 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 545394 0 545450 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 548890 0 548946 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 552386 0 552442 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 555882 0 555938 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 559378 0 559434 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 562874 0 562930 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 566370 0 566426 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 569866 0 569922 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 167366 0 167422 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 177854 0 177910 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 181350 0 181406 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 184846 0 184902 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 188342 0 188398 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 191838 0 191894 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 195334 0 195390 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 198830 0 198886 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 202326 0 202382 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 205822 0 205878 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 209318 0 209374 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 216402 0 216458 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 223394 0 223450 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 226890 0 226946 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 230386 0 230442 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 233882 0 233938 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 237378 0 237434 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 240874 0 240930 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 244370 0 244426 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 247866 0 247922 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 251362 0 251418 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 254858 0 254914 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 258354 0 258410 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 261850 0 261906 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 265346 0 265402 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 268842 0 268898 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 272338 0 272394 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 275834 0 275890 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 279330 0 279386 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 282826 0 282882 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 286322 0 286378 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 289910 0 289966 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 293406 0 293462 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 296902 0 296958 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 300398 0 300454 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 303894 0 303950 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 307390 0 307446 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 310886 0 310942 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 314382 0 314438 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 317878 0 317934 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 321374 0 321430 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 324870 0 324926 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 328366 0 328422 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 331862 0 331918 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 335358 0 335414 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 338854 0 338910 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 342350 0 342406 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 345846 0 345902 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 349342 0 349398 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 352838 0 352894 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 356334 0 356390 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 359830 0 359886 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 363326 0 363382 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 366914 0 366970 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 146390 0 146446 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 370410 0 370466 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 373906 0 373962 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 377402 0 377458 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 380898 0 380954 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 384394 0 384450 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 387890 0 387946 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 391386 0 391442 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 394882 0 394938 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 398378 0 398434 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 401874 0 401930 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 405370 0 405426 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 408866 0 408922 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 412362 0 412418 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 415858 0 415914 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 419354 0 419410 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 422850 0 422906 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 426346 0 426402 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 429842 0 429898 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 433338 0 433394 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 436834 0 436890 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 440330 0 440386 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 443826 0 443882 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 447414 0 447470 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 450910 0 450966 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 454406 0 454462 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 457902 0 457958 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 461398 0 461454 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 464894 0 464950 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 468390 0 468446 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 471886 0 471942 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 156878 0 156934 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 476578 0 476634 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 480074 0 480130 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 483570 0 483626 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 487066 0 487122 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 490562 0 490618 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 494058 0 494114 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 497554 0 497610 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 501050 0 501106 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 504546 0 504602 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 508042 0 508098 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 511538 0 511594 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 515034 0 515090 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 518530 0 518586 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 522026 0 522082 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 525522 0 525578 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 529018 0 529074 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 532514 0 532570 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 536010 0 536066 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 539506 0 539562 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 543002 0 543058 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 546498 0 546554 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 550086 0 550142 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 553582 0 553638 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 557078 0 557134 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 560574 0 560630 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 564070 0 564126 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 567566 0 567622 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 571062 0 571118 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 182546 0 182602 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 186042 0 186098 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 200026 0 200082 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 203522 0 203578 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 221002 0 221058 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 224498 0 224554 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 227994 0 228050 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 231490 0 231546 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 234986 0 235042 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 238574 0 238630 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 242070 0 242126 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 249062 0 249118 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 252558 0 252614 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 256054 0 256110 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 266542 0 266598 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 270038 0 270094 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 273534 0 273590 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 277030 0 277086 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 280526 0 280582 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 284022 0 284078 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 287518 0 287574 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 291014 0 291070 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 294510 0 294566 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 298006 0 298062 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 301502 0 301558 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 304998 0 305054 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 308494 0 308550 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 311990 0 312046 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 315578 0 315634 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 319074 0 319130 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 322570 0 322626 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 326066 0 326122 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 329562 0 329618 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 333058 0 333114 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 336554 0 336610 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 343546 0 343602 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 347042 0 347098 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 350538 0 350594 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 354034 0 354090 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 357530 0 357586 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 361026 0 361082 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 364522 0 364578 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 368018 0 368074 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 371514 0 371570 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 375010 0 375066 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 378506 0 378562 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 382002 0 382058 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 385498 0 385554 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 388994 0 389050 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 392490 0 392546 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 396078 0 396134 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 399574 0 399630 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 403070 0 403126 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 406566 0 406622 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 410062 0 410118 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 413558 0 413614 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 417054 0 417110 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 420550 0 420606 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 424046 0 424102 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 427542 0 427598 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 431038 0 431094 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 434534 0 434590 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 438030 0 438086 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 441526 0 441582 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 445022 0 445078 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 448518 0 448574 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 452014 0 452070 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 455510 0 455566 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 459006 0 459062 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 462502 0 462558 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 465998 0 466054 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 469494 0 469550 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 473082 0 473138 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 434288 2128 434608 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 465008 2128 465328 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 495728 2128 496048 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 526448 2128 526768 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 557168 2128 557488 692560 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 418928 2128 419248 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 449648 2128 449968 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 480368 2128 480688 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 511088 2128 511408 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 541808 2128 542128 692560 6 vssd1
port 503 nsew ground input
rlabel metal4 s 572528 2128 572848 692560 6 vssd1
port 503 nsew ground input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 575200 695200
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 901659320
string GDS_START 1530778
<< end >>

