magic
tech sky130A
magscale 1 2
timestamp 1636387369
<< locali >>
rect 232421 471631 232455 471801
rect 237757 471631 237791 471801
rect 152105 467891 152139 469013
rect 282193 39287 282227 40001
rect 330493 39831 330527 39933
rect 403081 39627 403115 39865
rect 31033 3247 31067 4029
rect 42809 3519 42843 3689
rect 38117 3179 38151 3349
rect 53757 3043 53791 3485
rect 57069 3315 57103 3825
rect 74733 3655 74767 3961
rect 307677 3111 307711 3417
rect 350365 3315 350399 4097
rect 358921 3859 358955 3961
rect 350365 3281 350549 3315
<< viali >>
rect 232421 471801 232455 471835
rect 232421 471597 232455 471631
rect 237757 471801 237791 471835
rect 237757 471597 237791 471631
rect 152105 469013 152139 469047
rect 152105 467857 152139 467891
rect 282193 40001 282227 40035
rect 330493 39933 330527 39967
rect 330493 39797 330527 39831
rect 403081 39865 403115 39899
rect 403081 39593 403115 39627
rect 282193 39253 282227 39287
rect 350365 4097 350399 4131
rect 31033 4029 31067 4063
rect 74733 3961 74767 3995
rect 57069 3825 57103 3859
rect 42809 3689 42843 3723
rect 42809 3485 42843 3519
rect 53757 3485 53791 3519
rect 31033 3213 31067 3247
rect 38117 3349 38151 3383
rect 38117 3145 38151 3179
rect 74733 3621 74767 3655
rect 57069 3281 57103 3315
rect 307677 3417 307711 3451
rect 358921 3961 358955 3995
rect 358921 3825 358955 3859
rect 350549 3281 350583 3315
rect 307677 3077 307711 3111
rect 53757 3009 53791 3043
<< metal1 >>
rect 238662 700952 238668 701004
rect 238720 700992 238726 701004
rect 397454 700992 397460 701004
rect 238720 700964 397460 700992
rect 238720 700952 238726 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 241422 700884 241428 700936
rect 241480 700924 241486 700936
rect 413646 700924 413652 700936
rect 241480 700896 413652 700924
rect 241480 700884 241486 700896
rect 413646 700884 413652 700896
rect 413704 700884 413710 700936
rect 89162 700816 89168 700868
rect 89220 700856 89226 700868
rect 296714 700856 296720 700868
rect 89220 700828 296720 700856
rect 89220 700816 89226 700828
rect 296714 700816 296720 700828
rect 296772 700816 296778 700868
rect 72970 700748 72976 700800
rect 73028 700788 73034 700800
rect 292574 700788 292580 700800
rect 73028 700760 292580 700788
rect 73028 700748 73034 700760
rect 292574 700748 292580 700760
rect 292632 700748 292638 700800
rect 227622 700680 227628 700732
rect 227680 700720 227686 700732
rect 462314 700720 462320 700732
rect 227680 700692 462320 700720
rect 227680 700680 227686 700692
rect 462314 700680 462320 700692
rect 462372 700680 462378 700732
rect 230382 700612 230388 700664
rect 230440 700652 230446 700664
rect 478506 700652 478512 700664
rect 230440 700624 478512 700652
rect 230440 700612 230446 700624
rect 478506 700612 478512 700624
rect 478564 700612 478570 700664
rect 40494 700544 40500 700596
rect 40552 700584 40558 700596
rect 300854 700584 300860 700596
rect 40552 700556 300860 700584
rect 40552 700544 40558 700556
rect 300854 700544 300860 700556
rect 300912 700544 300918 700596
rect 24302 700476 24308 700528
rect 24360 700516 24366 700528
rect 307754 700516 307760 700528
rect 24360 700488 307760 700516
rect 24360 700476 24366 700488
rect 307754 700476 307760 700488
rect 307812 700476 307818 700528
rect 8110 700408 8116 700460
rect 8168 700448 8174 700460
rect 303614 700448 303620 700460
rect 8168 700420 303620 700448
rect 8168 700408 8174 700420
rect 303614 700408 303620 700420
rect 303672 700408 303678 700460
rect 215202 700340 215208 700392
rect 215260 700380 215266 700392
rect 527174 700380 527180 700392
rect 215260 700352 527180 700380
rect 215260 700340 215266 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 219342 700272 219348 700324
rect 219400 700312 219406 700324
rect 543458 700312 543464 700324
rect 219400 700284 543464 700312
rect 219400 700272 219406 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 137830 700204 137836 700256
rect 137888 700244 137894 700256
rect 281534 700244 281540 700256
rect 137888 700216 281540 700244
rect 137888 700204 137894 700216
rect 281534 700204 281540 700216
rect 281592 700204 281598 700256
rect 154114 700136 154120 700188
rect 154172 700176 154178 700188
rect 285674 700176 285680 700188
rect 154172 700148 285680 700176
rect 154172 700136 154178 700148
rect 285674 700136 285680 700148
rect 285732 700136 285738 700188
rect 252462 700068 252468 700120
rect 252520 700108 252526 700120
rect 348786 700108 348792 700120
rect 252520 700080 348792 700108
rect 252520 700068 252526 700080
rect 348786 700068 348792 700080
rect 348844 700068 348850 700120
rect 249702 700000 249708 700052
rect 249760 700040 249766 700052
rect 332502 700040 332508 700052
rect 249760 700012 332508 700040
rect 249760 700000 249766 700012
rect 332502 700000 332508 700012
rect 332560 700000 332566 700052
rect 202782 699932 202788 699984
rect 202840 699972 202846 699984
rect 270494 699972 270500 699984
rect 202840 699944 270500 699972
rect 202840 699932 202846 699944
rect 270494 699932 270500 699944
rect 270552 699932 270558 699984
rect 218974 699864 218980 699916
rect 219032 699904 219038 699916
rect 274634 699904 274640 699916
rect 219032 699876 274640 699904
rect 219032 699864 219038 699876
rect 274634 699864 274640 699876
rect 274692 699864 274698 699916
rect 264882 699796 264888 699848
rect 264940 699836 264946 699848
rect 283834 699836 283840 699848
rect 264940 699808 283840 699836
rect 264940 699796 264946 699808
rect 283834 699796 283840 699808
rect 283892 699796 283898 699848
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 260742 699660 260748 699712
rect 260800 699700 260806 699712
rect 267642 699700 267648 699712
rect 260800 699672 267648 699700
rect 260800 699660 260806 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 204162 696940 204168 696992
rect 204220 696980 204226 696992
rect 580166 696980 580172 696992
rect 204220 696952 580172 696980
rect 204220 696940 204226 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 311894 683244 311900 683256
rect 3476 683216 311900 683244
rect 3476 683204 3482 683216
rect 311894 683204 311900 683216
rect 311952 683204 311958 683256
rect 208302 683136 208308 683188
rect 208360 683176 208366 683188
rect 580166 683176 580172 683188
rect 208360 683148 580172 683176
rect 208360 683136 208366 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3418 670760 3424 670812
rect 3476 670800 3482 670812
rect 318794 670800 318800 670812
rect 3476 670772 318800 670800
rect 3476 670760 3482 670772
rect 318794 670760 318800 670772
rect 318852 670760 318858 670812
rect 201402 670692 201408 670744
rect 201460 670732 201466 670744
rect 580166 670732 580172 670744
rect 201460 670704 580172 670732
rect 201460 670692 201466 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 314654 656928 314660 656940
rect 3476 656900 314660 656928
rect 3476 656888 3482 656900
rect 314654 656888 314660 656900
rect 314712 656888 314718 656940
rect 193122 643084 193128 643136
rect 193180 643124 193186 643136
rect 580166 643124 580172 643136
rect 193180 643096 580172 643124
rect 193180 643084 193186 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 322934 632108 322940 632120
rect 3476 632080 322940 632108
rect 3476 632068 3482 632080
rect 322934 632068 322940 632080
rect 322992 632068 322998 632120
rect 197262 630640 197268 630692
rect 197320 630680 197326 630692
rect 580166 630680 580172 630692
rect 197320 630652 580172 630680
rect 197320 630640 197326 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 329834 618304 329840 618316
rect 3200 618276 329840 618304
rect 3200 618264 3206 618276
rect 329834 618264 329840 618276
rect 329892 618264 329898 618316
rect 190362 616836 190368 616888
rect 190420 616876 190426 616888
rect 580166 616876 580172 616888
rect 190420 616848 580172 616876
rect 190420 616836 190426 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 325694 605860 325700 605872
rect 3292 605832 325700 605860
rect 3292 605820 3298 605832
rect 325694 605820 325700 605832
rect 325752 605820 325758 605872
rect 182082 590656 182088 590708
rect 182140 590696 182146 590708
rect 579798 590696 579804 590708
rect 182140 590668 579804 590696
rect 182140 590656 182146 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 333974 579680 333980 579692
rect 3384 579652 333980 579680
rect 3384 579640 3390 579652
rect 333974 579640 333980 579652
rect 334032 579640 334038 579692
rect 186222 576852 186228 576904
rect 186280 576892 186286 576904
rect 580166 576892 580172 576904
rect 186280 576864 580172 576892
rect 186280 576852 186286 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 340874 565876 340880 565888
rect 3476 565848 340880 565876
rect 3476 565836 3482 565848
rect 340874 565836 340880 565848
rect 340932 565836 340938 565888
rect 177942 563048 177948 563100
rect 178000 563088 178006 563100
rect 579798 563088 579804 563100
rect 178000 563060 579804 563088
rect 178000 563048 178006 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 338114 553432 338120 553444
rect 3476 553404 338120 553432
rect 3476 553392 3482 553404
rect 338114 553392 338120 553404
rect 338172 553392 338178 553444
rect 170950 536800 170956 536852
rect 171008 536840 171014 536852
rect 580166 536840 580172 536852
rect 171008 536812 580172 536840
rect 171008 536800 171014 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 345014 527184 345020 527196
rect 3476 527156 345020 527184
rect 3476 527144 3482 527156
rect 345014 527144 345020 527156
rect 345072 527144 345078 527196
rect 175182 524424 175188 524476
rect 175240 524464 175246 524476
rect 580166 524464 580172 524476
rect 175240 524436 580172 524464
rect 175240 524424 175246 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 351914 514808 351920 514820
rect 3476 514780 351920 514808
rect 3476 514768 3482 514780
rect 351914 514768 351920 514780
rect 351972 514768 351978 514820
rect 166902 510620 166908 510672
rect 166960 510660 166966 510672
rect 580166 510660 580172 510672
rect 166960 510632 580172 510660
rect 166960 510620 166966 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 349154 501004 349160 501016
rect 3108 500976 349160 501004
rect 3108 500964 3114 500976
rect 349154 500964 349160 500976
rect 349212 500964 349218 501016
rect 160002 484372 160008 484424
rect 160060 484412 160066 484424
rect 580166 484412 580172 484424
rect 160060 484384 580172 484412
rect 160060 484372 160066 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 356238 474756 356244 474768
rect 3476 474728 356244 474756
rect 3476 474716 3482 474728
rect 356238 474716 356244 474728
rect 356296 474716 356302 474768
rect 22830 472132 22836 472184
rect 22888 472172 22894 472184
rect 386414 472172 386420 472184
rect 22888 472144 386420 472172
rect 22888 472132 22894 472144
rect 386414 472132 386420 472144
rect 386472 472132 386478 472184
rect 129642 472064 129648 472116
rect 129700 472104 129706 472116
rect 512638 472104 512644 472116
rect 129700 472076 512644 472104
rect 129700 472064 129706 472076
rect 512638 472064 512644 472076
rect 512696 472064 512702 472116
rect 85114 471996 85120 472048
rect 85172 472036 85178 472048
rect 511258 472036 511264 472048
rect 85172 472008 511264 472036
rect 85172 471996 85178 472008
rect 511258 471996 511264 472008
rect 511316 471996 511322 472048
rect 159542 471928 159548 471980
rect 159600 471968 159606 471980
rect 160002 471968 160008 471980
rect 159600 471940 160008 471968
rect 159600 471928 159606 471940
rect 160002 471928 160008 471940
rect 160060 471928 160066 471980
rect 174446 471928 174452 471980
rect 174504 471968 174510 471980
rect 175182 471968 175188 471980
rect 174504 471940 175188 471968
rect 174504 471928 174510 471940
rect 175182 471928 175188 471940
rect 175240 471928 175246 471980
rect 185670 471928 185676 471980
rect 185728 471968 185734 471980
rect 186222 471968 186228 471980
rect 185728 471940 186228 471968
rect 185728 471928 185734 471940
rect 186222 471928 186228 471940
rect 186280 471928 186286 471980
rect 189350 471928 189356 471980
rect 189408 471968 189414 471980
rect 190362 471968 190368 471980
rect 189408 471940 190368 471968
rect 189408 471928 189414 471940
rect 190362 471928 190368 471940
rect 190420 471928 190426 471980
rect 196802 471928 196808 471980
rect 196860 471968 196866 471980
rect 197262 471968 197268 471980
rect 196860 471940 197268 471968
rect 196860 471928 196866 471940
rect 197262 471928 197268 471940
rect 197320 471928 197326 471980
rect 200574 471928 200580 471980
rect 200632 471968 200638 471980
rect 201402 471968 201408 471980
rect 200632 471940 201408 471968
rect 200632 471928 200638 471940
rect 201402 471928 201408 471940
rect 201460 471928 201466 471980
rect 226610 471928 226616 471980
rect 226668 471968 226674 471980
rect 227622 471968 227628 471980
rect 226668 471940 227628 471968
rect 226668 471928 226674 471940
rect 227622 471928 227628 471940
rect 227680 471928 227686 471980
rect 248966 471928 248972 471980
rect 249024 471968 249030 471980
rect 249702 471968 249708 471980
rect 249024 471940 249708 471968
rect 249024 471928 249030 471940
rect 249702 471928 249708 471940
rect 249760 471928 249766 471980
rect 260098 471928 260104 471980
rect 260156 471968 260162 471980
rect 260742 471968 260748 471980
rect 260156 471940 260748 471968
rect 260156 471928 260162 471940
rect 260742 471928 260748 471940
rect 260800 471928 260806 471980
rect 263870 471928 263876 471980
rect 263928 471968 263934 471980
rect 264882 471968 264888 471980
rect 263928 471940 264888 471968
rect 263928 471928 263934 471940
rect 264882 471928 264888 471940
rect 264940 471928 264946 471980
rect 235902 471860 235908 471912
rect 235960 471900 235966 471912
rect 266906 471900 266912 471912
rect 235960 471872 266912 471900
rect 235960 471860 235966 471872
rect 266906 471860 266912 471872
rect 266964 471860 266970 471912
rect 232409 471835 232467 471841
rect 232409 471801 232421 471835
rect 232455 471832 232467 471835
rect 237745 471835 237803 471841
rect 237745 471832 237757 471835
rect 232455 471804 237757 471832
rect 232455 471801 232467 471804
rect 232409 471795 232467 471801
rect 237745 471801 237757 471804
rect 237791 471801 237803 471835
rect 237745 471795 237803 471801
rect 256418 471792 256424 471844
rect 256476 471832 256482 471844
rect 299474 471832 299480 471844
rect 256476 471804 299480 471832
rect 256476 471792 256482 471804
rect 299474 471792 299480 471804
rect 299532 471792 299538 471844
rect 171042 471724 171048 471776
rect 171100 471764 171106 471776
rect 278130 471764 278136 471776
rect 171100 471736 278136 471764
rect 171100 471724 171106 471736
rect 278130 471724 278136 471736
rect 278188 471724 278194 471776
rect 81342 471656 81348 471708
rect 81400 471696 81406 471708
rect 81400 471668 232544 471696
rect 81400 471656 81406 471668
rect 106182 471588 106188 471640
rect 106240 471628 106246 471640
rect 232409 471631 232467 471637
rect 232409 471628 232421 471631
rect 106240 471600 232421 471628
rect 106240 471588 106246 471600
rect 232409 471597 232421 471600
rect 232455 471597 232467 471631
rect 232409 471591 232467 471597
rect 148410 471520 148416 471572
rect 148468 471560 148474 471572
rect 223390 471560 223396 471572
rect 148468 471532 223396 471560
rect 148468 471520 148474 471532
rect 223390 471520 223396 471532
rect 223448 471520 223454 471572
rect 232516 471560 232544 471668
rect 234062 471656 234068 471708
rect 234120 471696 234126 471708
rect 234120 471668 237696 471696
rect 234120 471656 234126 471668
rect 234982 471560 234988 471572
rect 232516 471532 234988 471560
rect 234982 471520 234988 471532
rect 235040 471520 235046 471572
rect 237668 471560 237696 471668
rect 237834 471656 237840 471708
rect 237892 471696 237898 471708
rect 238662 471696 238668 471708
rect 237892 471668 238668 471696
rect 237892 471656 237898 471668
rect 238662 471656 238668 471668
rect 238720 471656 238726 471708
rect 245286 471656 245292 471708
rect 245344 471696 245350 471708
rect 364334 471696 364340 471708
rect 245344 471668 364340 471696
rect 245344 471656 245350 471668
rect 364334 471656 364340 471668
rect 364392 471656 364398 471708
rect 237745 471631 237803 471637
rect 237745 471597 237757 471631
rect 237791 471628 237803 471631
rect 289262 471628 289268 471640
rect 237791 471600 289268 471628
rect 237791 471597 237803 471600
rect 237745 471591 237803 471597
rect 289262 471588 289268 471600
rect 289320 471588 289326 471640
rect 429194 471560 429200 471572
rect 237668 471532 429200 471560
rect 429194 471520 429200 471532
rect 429252 471520 429258 471572
rect 222930 471452 222936 471504
rect 222988 471492 222994 471504
rect 494054 471492 494060 471504
rect 222988 471464 494060 471492
rect 222988 471452 222994 471464
rect 494054 471452 494060 471464
rect 494112 471452 494118 471504
rect 140682 471384 140688 471436
rect 140740 471424 140746 471436
rect 467374 471424 467380 471436
rect 140740 471396 467380 471424
rect 140740 471384 140746 471396
rect 467374 471384 467380 471396
rect 467432 471384 467438 471436
rect 211706 471316 211712 471368
rect 211764 471356 211770 471368
rect 558914 471356 558920 471368
rect 211764 471328 558920 471356
rect 211764 471316 211770 471328
rect 558914 471316 558920 471328
rect 558972 471316 558978 471368
rect 118602 471248 118608 471300
rect 118660 471288 118666 471300
rect 467282 471288 467288 471300
rect 118660 471260 467288 471288
rect 118660 471248 118666 471260
rect 467282 471248 467288 471260
rect 467340 471248 467346 471300
rect 107470 471180 107476 471232
rect 107528 471220 107534 471232
rect 467190 471220 467196 471232
rect 107528 471192 467196 471220
rect 107528 471180 107534 471192
rect 467190 471180 467196 471192
rect 467248 471180 467254 471232
rect 96246 471112 96252 471164
rect 96304 471152 96310 471164
rect 467098 471152 467104 471164
rect 96304 471124 467104 471152
rect 96304 471112 96310 471124
rect 467098 471112 467104 471124
rect 467156 471112 467162 471164
rect 29730 471044 29736 471096
rect 29788 471084 29794 471096
rect 408494 471084 408500 471096
rect 29788 471056 408500 471084
rect 29788 471044 29794 471056
rect 408494 471044 408500 471056
rect 408552 471044 408558 471096
rect 32398 470976 32404 471028
rect 32456 471016 32462 471028
rect 419626 471016 419632 471028
rect 32456 470988 419632 471016
rect 32456 470976 32462 470988
rect 419626 470976 419632 470988
rect 419684 470976 419690 471028
rect 33778 470908 33784 470960
rect 33836 470948 33842 470960
rect 430850 470948 430856 470960
rect 33836 470920 430856 470948
rect 33836 470908 33842 470920
rect 430850 470908 430856 470920
rect 430908 470908 430914 470960
rect 92382 470840 92388 470892
rect 92440 470880 92446 470892
rect 497458 470880 497464 470892
rect 92440 470852 497464 470880
rect 92440 470840 92446 470852
rect 497458 470840 497464 470852
rect 497516 470840 497522 470892
rect 35158 470772 35164 470824
rect 35216 470812 35222 470824
rect 441982 470812 441988 470824
rect 35216 470784 441988 470812
rect 35216 470772 35222 470784
rect 441982 470772 441988 470784
rect 442040 470772 442046 470824
rect 36538 470704 36544 470756
rect 36596 470744 36602 470756
rect 453206 470744 453212 470756
rect 36596 470716 453212 470744
rect 36596 470704 36602 470716
rect 453206 470704 453212 470716
rect 453264 470704 453270 470756
rect 163314 470636 163320 470688
rect 163372 470676 163378 470688
rect 580166 470676 580172 470688
rect 163372 470648 580172 470676
rect 163372 470636 163378 470648
rect 580166 470636 580172 470648
rect 580224 470636 580230 470688
rect 40678 470568 40684 470620
rect 40736 470608 40742 470620
rect 464338 470608 464344 470620
rect 40736 470580 464344 470608
rect 40736 470568 40742 470580
rect 464338 470568 464344 470580
rect 464396 470568 464402 470620
rect 155862 470364 155868 470416
rect 155920 470404 155926 470416
rect 468478 470404 468484 470416
rect 155920 470376 468484 470404
rect 155920 470364 155926 470376
rect 468478 470364 468484 470376
rect 468536 470364 468542 470416
rect 39390 470296 39396 470348
rect 39448 470336 39454 470348
rect 389818 470336 389824 470348
rect 39448 470308 389824 470336
rect 39448 470296 39454 470308
rect 389818 470296 389824 470308
rect 389876 470296 389882 470348
rect 133506 470228 133512 470280
rect 133564 470268 133570 470280
rect 486418 470268 486424 470280
rect 133564 470240 486424 470268
rect 133564 470228 133570 470240
rect 486418 470228 486424 470240
rect 486476 470228 486482 470280
rect 223390 470160 223396 470212
rect 223448 470200 223454 470212
rect 580442 470200 580448 470212
rect 223448 470172 580448 470200
rect 223448 470160 223454 470172
rect 580442 470160 580448 470172
rect 580500 470160 580506 470212
rect 3602 470092 3608 470144
rect 3660 470132 3666 470144
rect 367462 470132 367468 470144
rect 3660 470104 367468 470132
rect 3660 470092 3666 470104
rect 367462 470092 367468 470104
rect 367520 470092 367526 470144
rect 111150 470024 111156 470076
rect 111208 470064 111214 470076
rect 483658 470064 483664 470076
rect 111208 470036 483664 470064
rect 111208 470024 111214 470036
rect 483658 470024 483664 470036
rect 483716 470024 483722 470076
rect 15838 469956 15844 470008
rect 15896 469996 15902 470008
rect 393590 469996 393596 470008
rect 15896 469968 393596 469996
rect 15896 469956 15902 469968
rect 393590 469956 393596 469968
rect 393648 469956 393654 470008
rect 88794 469888 88800 469940
rect 88852 469928 88858 469940
rect 479518 469928 479524 469940
rect 88852 469900 479524 469928
rect 88852 469888 88858 469900
rect 479518 469888 479524 469900
rect 479576 469888 479582 469940
rect 18598 469820 18604 469872
rect 18656 469860 18662 469872
rect 412174 469860 412180 469872
rect 18656 469832 412180 469860
rect 18656 469820 18662 469832
rect 412174 469820 412180 469832
rect 412232 469820 412238 469872
rect 103238 469752 103244 469804
rect 103296 469792 103302 469804
rect 500218 469792 500224 469804
rect 103296 469764 500224 469792
rect 103296 469752 103302 469764
rect 500218 469752 500224 469764
rect 500276 469752 500282 469804
rect 17218 469684 17224 469736
rect 17276 469724 17282 469736
rect 415946 469724 415952 469736
rect 17276 469696 415952 469724
rect 17276 469684 17282 469696
rect 415946 469684 415952 469696
rect 416004 469684 416010 469736
rect 65978 469616 65984 469668
rect 66036 469656 66042 469668
rect 472618 469656 472624 469668
rect 66036 469628 472624 469656
rect 66036 469616 66042 469628
rect 472618 469616 472624 469628
rect 472676 469616 472682 469668
rect 21358 469548 21364 469600
rect 21416 469588 21422 469600
rect 434714 469588 434720 469600
rect 21416 469560 434720 469588
rect 21416 469548 21422 469560
rect 434714 469548 434720 469560
rect 434772 469548 434778 469600
rect 70210 469480 70216 469532
rect 70268 469520 70274 469532
rect 493318 469520 493324 469532
rect 70268 469492 493324 469520
rect 70268 469480 70274 469492
rect 493318 469480 493324 469492
rect 493376 469480 493382 469532
rect 7558 469412 7564 469464
rect 7616 469452 7622 469464
rect 438302 469452 438308 469464
rect 7616 469424 438308 469452
rect 7616 469412 7622 469424
rect 438302 469412 438308 469424
rect 438360 469412 438366 469464
rect 29638 469344 29644 469396
rect 29696 469384 29702 469396
rect 461118 469384 461124 469396
rect 29696 469356 461124 469384
rect 29696 469344 29702 469356
rect 461118 469344 461124 469356
rect 461176 469344 461182 469396
rect 58986 469276 58992 469328
rect 59044 469316 59050 469328
rect 490558 469316 490564 469328
rect 59044 469288 490564 469316
rect 59044 469276 59050 469288
rect 490558 469276 490564 469288
rect 490616 469276 490622 469328
rect 11698 469208 11704 469260
rect 11756 469248 11762 469260
rect 456886 469248 456892 469260
rect 11756 469220 456892 469248
rect 11756 469208 11762 469220
rect 456886 469208 456892 469220
rect 456944 469208 456950 469260
rect 152090 469044 152096 469056
rect 152051 469016 152096 469044
rect 152090 469004 152096 469016
rect 152148 469004 152154 469056
rect 234982 469004 234988 469056
rect 235040 469044 235046 469056
rect 580258 469044 580264 469056
rect 235040 469016 580264 469044
rect 235040 469004 235046 469016
rect 580258 469004 580264 469016
rect 580316 469004 580322 469056
rect 15930 468936 15936 468988
rect 15988 468976 15994 468988
rect 360194 468976 360200 468988
rect 15988 468948 360200 468976
rect 15988 468936 15994 468948
rect 360194 468936 360200 468948
rect 360252 468936 360258 468988
rect 144730 468868 144736 468920
rect 144788 468908 144794 468920
rect 489178 468908 489184 468920
rect 144788 468880 489184 468908
rect 144788 468868 144794 468880
rect 489178 468868 489184 468880
rect 489236 468868 489242 468920
rect 17310 468800 17316 468852
rect 17368 468840 17374 468852
rect 371556 468840 371562 468852
rect 17368 468812 371562 468840
rect 17368 468800 17374 468812
rect 371556 468800 371562 468812
rect 371614 468800 371620 468852
rect 122374 468732 122380 468784
rect 122432 468772 122438 468784
rect 485038 468772 485044 468784
rect 122432 468744 485044 468772
rect 122432 468732 122438 468744
rect 485038 468732 485044 468744
rect 485096 468732 485102 468784
rect 4890 468664 4896 468716
rect 4948 468704 4954 468716
rect 378686 468704 378692 468716
rect 4948 468676 378692 468704
rect 4948 468664 4954 468676
rect 378686 468664 378692 468676
rect 378744 468664 378750 468716
rect 7650 468596 7656 468648
rect 7708 468636 7714 468648
rect 382366 468636 382372 468648
rect 7708 468608 382372 468636
rect 7708 468596 7714 468608
rect 382366 468596 382372 468608
rect 382424 468596 382430 468648
rect 100018 468528 100024 468580
rect 100076 468568 100082 468580
rect 482278 468568 482284 468580
rect 100076 468540 482284 468568
rect 100076 468528 100082 468540
rect 482278 468528 482284 468540
rect 482336 468528 482342 468580
rect 14458 468460 14464 468512
rect 14516 468500 14522 468512
rect 401042 468500 401048 468512
rect 14516 468472 401048 468500
rect 14516 468460 14522 468472
rect 401042 468460 401048 468472
rect 401100 468460 401106 468512
rect 114922 468392 114928 468444
rect 114980 468432 114986 468444
rect 501598 468432 501604 468444
rect 114980 468404 501604 468432
rect 114980 468392 114986 468404
rect 501598 468392 501604 468404
rect 501656 468392 501662 468444
rect 77662 468324 77668 468376
rect 77720 468364 77726 468376
rect 475378 468364 475384 468376
rect 77720 468336 475384 468364
rect 77720 468324 77726 468336
rect 475378 468324 475384 468336
rect 475436 468324 475442 468376
rect 25498 468256 25504 468308
rect 25556 468296 25562 468308
rect 423582 468296 423588 468308
rect 25556 468268 423588 468296
rect 25556 468256 25562 468268
rect 423582 468256 423588 468268
rect 423640 468256 423646 468308
rect 3510 468188 3516 468240
rect 3568 468228 3574 468240
rect 404722 468228 404728 468240
rect 3568 468200 404728 468228
rect 3568 468188 3574 468200
rect 404722 468188 404728 468200
rect 404780 468188 404786 468240
rect 39298 468120 39304 468172
rect 39356 468160 39362 468172
rect 449434 468160 449440 468172
rect 39356 468132 449440 468160
rect 39356 468120 39362 468132
rect 449434 468120 449440 468132
rect 449492 468120 449498 468172
rect 55122 468052 55128 468104
rect 55180 468092 55186 468104
rect 471238 468092 471244 468104
rect 55180 468064 471244 468092
rect 55180 468052 55186 468064
rect 471238 468052 471244 468064
rect 471296 468052 471302 468104
rect 4798 467984 4804 468036
rect 4856 468024 4862 468036
rect 427078 468024 427084 468036
rect 4856 467996 427084 468024
rect 4856 467984 4862 467996
rect 427078 467984 427084 467996
rect 427136 467984 427142 468036
rect 445754 468024 445760 468036
rect 431926 467996 445760 468024
rect 22738 467916 22744 467968
rect 22796 467956 22802 467968
rect 431926 467956 431954 467996
rect 445754 467984 445760 467996
rect 445812 467984 445818 468036
rect 22796 467928 431954 467956
rect 22796 467916 22802 467928
rect 152093 467891 152151 467897
rect 152093 467857 152105 467891
rect 152139 467888 152151 467891
rect 580350 467888 580356 467900
rect 152139 467860 580356 467888
rect 152139 467857 152151 467860
rect 152093 467851 152151 467857
rect 580350 467848 580356 467860
rect 580408 467848 580414 467900
rect 3418 463632 3424 463684
rect 3476 463672 3482 463684
rect 13814 463672 13820 463684
rect 3476 463644 13820 463672
rect 3476 463632 3482 463644
rect 13814 463632 13820 463644
rect 13872 463632 13878 463684
rect 468478 458124 468484 458176
rect 468536 458164 468542 458176
rect 580166 458164 580172 458176
rect 468536 458136 580172 458164
rect 468536 458124 468542 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 15930 449868 15936 449880
rect 3384 449840 15936 449868
rect 3384 449828 3390 449840
rect 15930 449828 15936 449840
rect 15988 449828 15994 449880
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 40770 411244 40776 411256
rect 3016 411216 40776 411244
rect 3016 411204 3022 411216
rect 40770 411204 40776 411216
rect 40828 411204 40834 411256
rect 489178 405628 489184 405680
rect 489236 405668 489242 405680
rect 579614 405668 579620 405680
rect 489236 405640 579620 405668
rect 489236 405628 489242 405640
rect 579614 405628 579620 405640
rect 579672 405628 579678 405680
rect 3234 398760 3240 398812
rect 3292 398800 3298 398812
rect 17310 398800 17316 398812
rect 3292 398772 17316 398800
rect 3292 398760 3298 398772
rect 17310 398760 17316 398772
rect 17368 398760 17374 398812
rect 504358 379448 504364 379500
rect 504416 379488 504422 379500
rect 580166 379488 580172 379500
rect 504416 379460 580172 379488
rect 504416 379448 504422 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 2774 371356 2780 371408
rect 2832 371396 2838 371408
rect 4890 371396 4896 371408
rect 2832 371368 4896 371396
rect 2832 371356 2838 371368
rect 4890 371356 4896 371368
rect 4948 371356 4954 371408
rect 467374 365644 467380 365696
rect 467432 365684 467438 365696
rect 580166 365684 580172 365696
rect 467432 365656 580172 365684
rect 467432 365644 467438 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 22830 358748 22836 358760
rect 3384 358720 22836 358748
rect 3384 358708 3390 358720
rect 22830 358708 22836 358720
rect 22888 358708 22894 358760
rect 486418 353200 486424 353252
rect 486476 353240 486482 353252
rect 580166 353240 580172 353252
rect 486476 353212 580172 353240
rect 486476 353200 486482 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 7650 346372 7656 346384
rect 3200 346344 7656 346372
rect 3200 346332 3206 346344
rect 7650 346332 7656 346344
rect 7708 346332 7714 346384
rect 502978 325592 502984 325644
rect 503036 325632 503042 325644
rect 579890 325632 579896 325644
rect 503036 325604 579896 325632
rect 503036 325592 503042 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 3510 320084 3516 320136
rect 3568 320124 3574 320136
rect 39390 320124 39396 320136
rect 3568 320096 39396 320124
rect 3568 320084 3574 320096
rect 39390 320084 39396 320096
rect 39448 320084 39454 320136
rect 512638 313216 512644 313268
rect 512696 313256 512702 313268
rect 580166 313256 580172 313268
rect 512696 313228 580172 313256
rect 512696 313216 512702 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 35250 306320 35256 306332
rect 3568 306292 35256 306320
rect 3568 306280 3574 306292
rect 35250 306280 35256 306292
rect 35308 306280 35314 306332
rect 485038 299412 485044 299464
rect 485096 299452 485102 299464
rect 579614 299452 579620 299464
rect 485096 299424 579620 299452
rect 485096 299412 485102 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 15838 293944 15844 293956
rect 3108 293916 15844 293944
rect 3108 293904 3114 293916
rect 15838 293904 15844 293916
rect 15896 293904 15902 293956
rect 501598 273164 501604 273216
rect 501656 273204 501662 273216
rect 579890 273204 579896 273216
rect 501656 273176 579896 273204
rect 501656 273164 501662 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 14458 267696 14464 267708
rect 3568 267668 14464 267696
rect 3568 267656 3574 267668
rect 14458 267656 14464 267668
rect 14516 267656 14522 267708
rect 467282 259360 467288 259412
rect 467340 259400 467346 259412
rect 579798 259400 579804 259412
rect 467340 259372 579804 259400
rect 467340 259360 467346 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 29730 255252 29736 255264
rect 3200 255224 29736 255252
rect 3200 255212 3206 255224
rect 29730 255212 29736 255224
rect 29788 255212 29794 255264
rect 483658 245556 483664 245608
rect 483716 245596 483722 245608
rect 580166 245596 580172 245608
rect 483716 245568 580172 245596
rect 483716 245556 483722 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 500218 233180 500224 233232
rect 500276 233220 500282 233232
rect 580166 233220 580172 233232
rect 500276 233192 580172 233220
rect 500276 233180 500282 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 467190 219376 467196 219428
rect 467248 219416 467254 219428
rect 579890 219416 579896 219428
rect 467248 219388 579896 219416
rect 467248 219376 467254 219388
rect 579890 219376 579896 219388
rect 579948 219376 579954 219428
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 18598 215268 18604 215280
rect 3384 215240 18604 215268
rect 3384 215228 3390 215240
rect 18598 215228 18604 215240
rect 18656 215228 18662 215280
rect 482278 206932 482284 206984
rect 482336 206972 482342 206984
rect 580166 206972 580172 206984
rect 482336 206944 580172 206972
rect 482336 206932 482342 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 32398 202824 32404 202836
rect 3476 202796 32404 202824
rect 3476 202784 3482 202796
rect 32398 202784 32404 202796
rect 32456 202784 32462 202836
rect 497458 193128 497464 193180
rect 497516 193168 497522 193180
rect 580166 193168 580172 193180
rect 497516 193140 580172 193168
rect 497516 193128 497522 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 17218 189020 17224 189032
rect 3476 188992 17224 189020
rect 3476 188980 3482 188992
rect 17218 188980 17224 188992
rect 17276 188980 17282 189032
rect 467098 179324 467104 179376
rect 467156 179364 467162 179376
rect 579982 179364 579988 179376
rect 467156 179336 579988 179364
rect 467156 179324 467162 179336
rect 579982 179324 579988 179336
rect 580040 179324 580046 179376
rect 479518 166948 479524 167000
rect 479576 166988 479582 167000
rect 580166 166988 580172 167000
rect 479576 166960 580172 166988
rect 479576 166948 479582 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 25498 164200 25504 164212
rect 3292 164172 25504 164200
rect 3292 164160 3298 164172
rect 25498 164160 25504 164172
rect 25556 164160 25562 164212
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 33778 150396 33784 150408
rect 3476 150368 33784 150396
rect 3476 150356 3482 150368
rect 33778 150356 33784 150368
rect 33836 150356 33842 150408
rect 511258 139340 511264 139392
rect 511316 139380 511322 139392
rect 580166 139380 580172 139392
rect 511316 139352 580172 139380
rect 511316 139340 511322 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 2774 137096 2780 137148
rect 2832 137136 2838 137148
rect 4798 137136 4804 137148
rect 2832 137108 4804 137136
rect 2832 137096 2838 137108
rect 4798 137096 4804 137108
rect 4856 137096 4862 137148
rect 475378 126896 475384 126948
rect 475436 126936 475442 126948
rect 580166 126936 580172 126948
rect 475436 126908 580172 126936
rect 475436 126896 475442 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 493318 113092 493324 113144
rect 493376 113132 493382 113144
rect 579798 113132 579804 113144
rect 493376 113104 579804 113132
rect 493376 113092 493382 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 21358 111772 21364 111784
rect 3476 111744 21364 111772
rect 3476 111732 3482 111744
rect 21358 111732 21364 111744
rect 21416 111732 21422 111784
rect 508498 100648 508504 100700
rect 508556 100688 508562 100700
rect 580166 100688 580172 100700
rect 508556 100660 580172 100688
rect 508556 100648 508562 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 35158 97968 35164 97980
rect 3476 97940 35164 97968
rect 3476 97928 3482 97940
rect 35158 97928 35164 97940
rect 35216 97928 35222 97980
rect 472618 86912 472624 86964
rect 472676 86952 472682 86964
rect 580166 86952 580172 86964
rect 472676 86924 580172 86952
rect 472676 86912 472682 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 7558 85524 7564 85536
rect 3200 85496 7564 85524
rect 3200 85484 3206 85496
rect 7558 85484 7564 85496
rect 7616 85484 7622 85536
rect 490558 73108 490564 73160
rect 490616 73148 490622 73160
rect 580166 73148 580172 73160
rect 490616 73120 580172 73148
rect 490616 73108 490622 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 22738 71720 22744 71732
rect 3476 71692 22744 71720
rect 3476 71680 3482 71692
rect 22738 71680 22744 71692
rect 22796 71680 22802 71732
rect 507118 60664 507124 60716
rect 507176 60704 507182 60716
rect 580166 60704 580172 60716
rect 507176 60676 580172 60704
rect 507176 60664 507182 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 36538 59344 36544 59356
rect 3108 59316 36544 59344
rect 3108 59304 3114 59316
rect 36538 59304 36544 59316
rect 36596 59304 36602 59356
rect 471238 46860 471244 46912
rect 471296 46900 471302 46912
rect 580166 46900 580172 46912
rect 471296 46872 580172 46900
rect 471296 46860 471302 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 39298 45540 39304 45552
rect 3476 45512 39304 45540
rect 3476 45500 3482 45512
rect 39298 45500 39304 45512
rect 39356 45500 39362 45552
rect 56594 41828 56600 41880
rect 56652 41868 56658 41880
rect 57836 41868 57842 41880
rect 56652 41840 57842 41868
rect 56652 41828 56658 41840
rect 57836 41828 57842 41840
rect 57894 41828 57900 41880
rect 70486 41828 70492 41880
rect 70544 41868 70550 41880
rect 71636 41868 71642 41880
rect 70544 41840 71642 41868
rect 70544 41828 70550 41840
rect 71636 41828 71642 41840
rect 71694 41828 71700 41880
rect 26142 39992 26148 40044
rect 26200 40032 26206 40044
rect 60366 40032 60372 40044
rect 26200 40004 60372 40032
rect 26200 39992 26206 40004
rect 60366 39992 60372 40004
rect 60424 39992 60430 40044
rect 67542 39992 67548 40044
rect 67600 40032 67606 40044
rect 90542 40032 90548 40044
rect 67600 40004 90548 40032
rect 67600 39992 67606 40004
rect 90542 39992 90548 40004
rect 90600 39992 90606 40044
rect 95050 39992 95056 40044
rect 95108 40032 95114 40044
rect 111150 40032 111156 40044
rect 95108 40004 111156 40032
rect 95108 39992 95114 40004
rect 111150 39992 111156 40004
rect 111208 39992 111214 40044
rect 111610 39992 111616 40044
rect 111668 40032 111674 40044
rect 122374 40032 122380 40044
rect 111668 40004 122380 40032
rect 111668 39992 111674 40004
rect 122374 39992 122380 40004
rect 122432 39992 122438 40044
rect 128262 39992 128268 40044
rect 128320 40032 128326 40044
rect 134426 40032 134432 40044
rect 128320 40004 134432 40032
rect 128320 39992 128326 40004
rect 134426 39992 134432 40004
rect 134484 39992 134490 40044
rect 142062 39992 142068 40044
rect 142120 40032 142126 40044
rect 144730 40032 144736 40044
rect 142120 40004 144736 40032
rect 142120 39992 142126 40004
rect 144730 39992 144736 40004
rect 144788 39992 144794 40044
rect 266262 39992 266268 40044
rect 266320 40032 266326 40044
rect 282181 40035 282239 40041
rect 282181 40032 282193 40035
rect 266320 40004 282193 40032
rect 266320 39992 266326 40004
rect 282181 40001 282193 40004
rect 282227 40001 282239 40035
rect 282181 39995 282239 40001
rect 297266 39992 297272 40044
rect 297324 40032 297330 40044
rect 299198 40032 299204 40044
rect 297324 40004 299204 40032
rect 297324 39992 297330 40004
rect 299198 39992 299204 40004
rect 299256 39992 299262 40044
rect 301590 39992 301596 40044
rect 301648 40032 301654 40044
rect 322198 40032 322204 40044
rect 301648 40004 322204 40032
rect 301648 39992 301654 40004
rect 322198 39992 322204 40004
rect 322256 39992 322262 40044
rect 327442 39992 327448 40044
rect 327500 40032 327506 40044
rect 342898 40032 342904 40044
rect 327500 40004 342904 40032
rect 327500 39992 327506 40004
rect 342898 39992 342904 40004
rect 342956 39992 342962 40044
rect 393774 39992 393780 40044
rect 393832 40032 393838 40044
rect 481634 40032 481640 40044
rect 393832 40004 481640 40032
rect 393832 39992 393838 40004
rect 481634 39992 481640 40004
rect 481692 39992 481698 40044
rect 28902 39924 28908 39976
rect 28960 39964 28966 39976
rect 62114 39964 62120 39976
rect 28960 39936 62120 39964
rect 28960 39924 28966 39936
rect 62114 39924 62120 39936
rect 62172 39924 62178 39976
rect 64782 39924 64788 39976
rect 64840 39964 64846 39976
rect 88794 39964 88800 39976
rect 64840 39936 88800 39964
rect 64840 39924 64846 39936
rect 88794 39924 88800 39936
rect 88852 39924 88858 39976
rect 89622 39924 89628 39976
rect 89680 39964 89686 39976
rect 106918 39964 106924 39976
rect 89680 39936 106924 39964
rect 89680 39924 89686 39936
rect 106918 39924 106924 39936
rect 106976 39924 106982 39976
rect 108942 39924 108948 39976
rect 109000 39964 109006 39976
rect 120626 39964 120632 39976
rect 109000 39936 120632 39964
rect 109000 39924 109006 39936
rect 120626 39924 120632 39936
rect 120684 39924 120690 39976
rect 140682 39924 140688 39976
rect 140740 39964 140746 39976
rect 143902 39964 143908 39976
rect 140740 39936 143908 39964
rect 140740 39924 140746 39936
rect 143902 39924 143908 39936
rect 143960 39924 143966 39976
rect 255130 39924 255136 39976
rect 255188 39964 255194 39976
rect 255188 39936 258074 39964
rect 255188 39924 255194 39936
rect 24762 39856 24768 39908
rect 24820 39896 24826 39908
rect 59538 39896 59544 39908
rect 24820 39868 59544 39896
rect 24820 39856 24826 39868
rect 59538 39856 59544 39868
rect 59596 39856 59602 39908
rect 62022 39856 62028 39908
rect 62080 39896 62086 39908
rect 86218 39896 86224 39908
rect 62080 39868 86224 39896
rect 62080 39856 62086 39868
rect 86218 39856 86224 39868
rect 86276 39856 86282 39908
rect 86862 39856 86868 39908
rect 86920 39896 86926 39908
rect 104250 39896 104256 39908
rect 86920 39868 104256 39896
rect 86920 39856 86926 39868
rect 104250 39856 104256 39868
rect 104308 39856 104314 39908
rect 107562 39856 107568 39908
rect 107620 39896 107626 39908
rect 119798 39896 119804 39908
rect 107620 39868 119804 39896
rect 107620 39856 107626 39868
rect 119798 39856 119804 39868
rect 119856 39856 119862 39908
rect 126882 39856 126888 39908
rect 126940 39896 126946 39908
rect 133598 39896 133604 39908
rect 126940 39868 133604 39896
rect 126940 39856 126946 39868
rect 133598 39856 133604 39868
rect 133656 39856 133662 39908
rect 137922 39856 137928 39908
rect 137980 39896 137986 39908
rect 142154 39896 142160 39908
rect 137980 39868 142160 39896
rect 137980 39856 137986 39868
rect 142154 39856 142160 39868
rect 142212 39856 142218 39908
rect 258046 39896 258074 39936
rect 268010 39924 268016 39976
rect 268068 39964 268074 39976
rect 304258 39964 304264 39976
rect 268068 39936 304264 39964
rect 268068 39924 268074 39936
rect 304258 39924 304264 39936
rect 304316 39924 304322 39976
rect 319714 39924 319720 39976
rect 319772 39964 319778 39976
rect 330481 39967 330539 39973
rect 330481 39964 330493 39967
rect 319772 39936 330493 39964
rect 319772 39924 319778 39936
rect 330481 39933 330493 39936
rect 330527 39933 330539 39967
rect 330481 39927 330539 39933
rect 343818 39924 343824 39976
rect 343876 39964 343882 39976
rect 352558 39964 352564 39976
rect 343876 39936 352564 39964
rect 343876 39924 343882 39936
rect 352558 39924 352564 39936
rect 352616 39924 352622 39976
rect 391198 39924 391204 39976
rect 391256 39964 391262 39976
rect 478874 39964 478880 39976
rect 391256 39936 478880 39964
rect 391256 39924 391262 39936
rect 478874 39924 478880 39936
rect 478932 39924 478938 39976
rect 269666 39896 269672 39908
rect 258046 39868 269672 39896
rect 269666 39856 269672 39868
rect 269724 39856 269730 39908
rect 318058 39896 318064 39908
rect 277366 39868 318064 39896
rect 23382 39788 23388 39840
rect 23440 39828 23446 39840
rect 58618 39828 58624 39840
rect 23440 39800 58624 39828
rect 23440 39788 23446 39800
rect 58618 39788 58624 39800
rect 58676 39788 58682 39840
rect 60642 39788 60648 39840
rect 60700 39828 60706 39840
rect 85390 39828 85396 39840
rect 60700 39800 85396 39828
rect 60700 39788 60706 39800
rect 85390 39788 85396 39800
rect 85448 39788 85454 39840
rect 91002 39788 91008 39840
rect 91060 39828 91066 39840
rect 107746 39828 107752 39840
rect 91060 39800 107752 39828
rect 91060 39788 91066 39800
rect 107746 39788 107752 39800
rect 107804 39788 107810 39840
rect 110322 39788 110328 39840
rect 110380 39828 110386 39840
rect 121546 39828 121552 39840
rect 110380 39800 121552 39828
rect 110380 39788 110386 39800
rect 121546 39788 121552 39800
rect 121604 39788 121610 39840
rect 122742 39788 122748 39840
rect 122800 39828 122806 39840
rect 131114 39828 131120 39840
rect 122800 39800 131120 39828
rect 122800 39788 122806 39800
rect 131114 39788 131120 39800
rect 131172 39788 131178 39840
rect 244734 39788 244740 39840
rect 244792 39828 244798 39840
rect 262858 39828 262864 39840
rect 244792 39800 262864 39828
rect 244792 39788 244798 39800
rect 262858 39788 262864 39800
rect 262916 39788 262922 39840
rect 275738 39788 275744 39840
rect 275796 39828 275802 39840
rect 277366 39828 277394 39868
rect 318058 39856 318064 39868
rect 318116 39856 318122 39908
rect 325694 39856 325700 39908
rect 325752 39896 325758 39908
rect 359550 39896 359556 39908
rect 325752 39868 359556 39896
rect 325752 39856 325758 39868
rect 359550 39856 359556 39868
rect 359608 39856 359614 39908
rect 403069 39899 403127 39905
rect 403069 39865 403081 39899
rect 403115 39896 403127 39899
rect 486418 39896 486424 39908
rect 403115 39868 486424 39896
rect 403115 39865 403127 39868
rect 403069 39859 403127 39865
rect 486418 39856 486424 39868
rect 486476 39856 486482 39908
rect 275796 39800 277394 39828
rect 275796 39788 275802 39800
rect 281810 39788 281816 39840
rect 281868 39828 281874 39840
rect 327718 39828 327724 39840
rect 281868 39800 327724 39828
rect 281868 39788 281874 39800
rect 327718 39788 327724 39800
rect 327776 39788 327782 39840
rect 330481 39831 330539 39837
rect 330481 39797 330493 39831
rect 330527 39828 330539 39831
rect 335998 39828 336004 39840
rect 330527 39800 336004 39828
rect 330527 39797 330539 39800
rect 330481 39791 330539 39797
rect 335998 39788 336004 39800
rect 336056 39788 336062 39840
rect 348970 39788 348976 39840
rect 349028 39828 349034 39840
rect 363506 39828 363512 39840
rect 349028 39800 363512 39828
rect 349028 39788 349034 39800
rect 363506 39788 363512 39800
rect 363564 39788 363570 39840
rect 369670 39788 369676 39840
rect 369728 39828 369734 39840
rect 381538 39828 381544 39840
rect 369728 39800 381544 39828
rect 369728 39788 369734 39800
rect 381538 39788 381544 39800
rect 381596 39788 381602 39840
rect 398926 39788 398932 39840
rect 398984 39828 398990 39840
rect 489914 39828 489920 39840
rect 398984 39800 489920 39828
rect 398984 39788 398990 39800
rect 489914 39788 489920 39800
rect 489972 39788 489978 39840
rect 16482 39720 16488 39772
rect 16540 39760 16546 39772
rect 53466 39760 53472 39772
rect 16540 39732 53472 39760
rect 16540 39720 16546 39732
rect 53466 39720 53472 39732
rect 53524 39720 53530 39772
rect 63402 39720 63408 39772
rect 63460 39760 63466 39772
rect 87966 39760 87972 39772
rect 63460 39732 87972 39760
rect 63460 39720 63466 39732
rect 87966 39720 87972 39732
rect 88024 39720 88030 39772
rect 88242 39720 88248 39772
rect 88300 39760 88306 39772
rect 105998 39760 106004 39772
rect 88300 39732 106004 39760
rect 88300 39720 88306 39732
rect 105998 39720 106004 39732
rect 106056 39720 106062 39772
rect 111702 39720 111708 39772
rect 111760 39760 111766 39772
rect 123202 39760 123208 39772
rect 111760 39732 123208 39760
rect 111760 39720 111766 39732
rect 123202 39720 123208 39732
rect 123260 39720 123266 39772
rect 125502 39720 125508 39772
rect 125560 39760 125566 39772
rect 132678 39760 132684 39772
rect 125560 39732 132684 39760
rect 125560 39720 125566 39732
rect 132678 39720 132684 39732
rect 132736 39720 132742 39772
rect 257706 39720 257712 39772
rect 257764 39760 257770 39772
rect 276566 39760 276572 39772
rect 257764 39732 276572 39760
rect 257764 39720 257770 39732
rect 276566 39720 276572 39732
rect 276624 39720 276630 39772
rect 280062 39720 280068 39772
rect 280120 39760 280126 39772
rect 325694 39760 325700 39772
rect 280120 39732 325700 39760
rect 280120 39720 280126 39732
rect 325694 39720 325700 39732
rect 325752 39720 325758 39772
rect 326614 39720 326620 39772
rect 326672 39760 326678 39772
rect 359458 39760 359464 39772
rect 326672 39732 359464 39760
rect 326672 39720 326678 39732
rect 359458 39720 359464 39732
rect 359516 39720 359522 39772
rect 361850 39720 361856 39772
rect 361908 39760 361914 39772
rect 377306 39760 377312 39772
rect 361908 39732 377312 39760
rect 361908 39720 361914 39732
rect 377306 39720 377312 39732
rect 377364 39720 377370 39772
rect 402330 39720 402336 39772
rect 402388 39760 402394 39772
rect 493318 39760 493324 39772
rect 402388 39732 493324 39760
rect 402388 39720 402394 39732
rect 493318 39720 493324 39732
rect 493376 39720 493382 39772
rect 19242 39652 19248 39704
rect 19300 39692 19306 39704
rect 55214 39692 55220 39704
rect 19300 39664 55220 39692
rect 19300 39652 19306 39664
rect 55214 39652 55220 39664
rect 55272 39652 55278 39704
rect 57882 39652 57888 39704
rect 57940 39692 57946 39704
rect 83642 39692 83648 39704
rect 57940 39664 83648 39692
rect 57940 39652 57946 39664
rect 83642 39652 83648 39664
rect 83700 39652 83706 39704
rect 85482 39652 85488 39704
rect 85540 39692 85546 39704
rect 103514 39692 103520 39704
rect 85540 39664 103520 39692
rect 85540 39652 85546 39664
rect 103514 39652 103520 39664
rect 103572 39652 103578 39704
rect 104802 39652 104808 39704
rect 104860 39692 104866 39704
rect 118050 39692 118056 39704
rect 104860 39664 118056 39692
rect 104860 39652 104866 39664
rect 118050 39652 118056 39664
rect 118108 39652 118114 39704
rect 119982 39652 119988 39704
rect 120040 39692 120046 39704
rect 128446 39692 128452 39704
rect 120040 39664 128452 39692
rect 120040 39652 120046 39664
rect 128446 39652 128452 39664
rect 128504 39652 128510 39704
rect 242158 39652 242164 39704
rect 242216 39692 242222 39704
rect 251818 39692 251824 39704
rect 242216 39664 251824 39692
rect 242216 39652 242222 39664
rect 251818 39652 251824 39664
rect 251876 39652 251882 39704
rect 252554 39652 252560 39704
rect 252612 39692 252618 39704
rect 273898 39692 273904 39704
rect 252612 39664 273904 39692
rect 252612 39652 252618 39664
rect 273898 39652 273904 39664
rect 273956 39652 273962 39704
rect 283558 39652 283564 39704
rect 283616 39692 283622 39704
rect 331214 39692 331220 39704
rect 283616 39664 331220 39692
rect 283616 39652 283622 39664
rect 331214 39652 331220 39664
rect 331272 39652 331278 39704
rect 333514 39652 333520 39704
rect 333572 39692 333578 39704
rect 349706 39692 349712 39704
rect 333572 39664 349712 39692
rect 333572 39652 333578 39664
rect 349706 39652 349712 39664
rect 349764 39652 349770 39704
rect 351546 39652 351552 39704
rect 351604 39692 351610 39704
rect 396718 39692 396724 39704
rect 351604 39664 396724 39692
rect 351604 39652 351610 39664
rect 396718 39652 396724 39664
rect 396776 39652 396782 39704
rect 404078 39652 404084 39704
rect 404136 39692 404142 39704
rect 496814 39692 496820 39704
rect 404136 39664 496820 39692
rect 404136 39652 404142 39664
rect 496814 39652 496820 39664
rect 496872 39652 496878 39704
rect 15102 39584 15108 39636
rect 15160 39624 15166 39636
rect 52638 39624 52644 39636
rect 15160 39596 52644 39624
rect 15160 39584 15166 39596
rect 52638 39584 52644 39596
rect 52696 39584 52702 39636
rect 53742 39584 53748 39636
rect 53800 39624 53806 39636
rect 81066 39624 81072 39636
rect 53800 39596 81072 39624
rect 53800 39584 53806 39596
rect 81066 39584 81072 39596
rect 81124 39584 81130 39636
rect 84102 39584 84108 39636
rect 84160 39624 84166 39636
rect 102594 39624 102600 39636
rect 84160 39596 102600 39624
rect 84160 39584 84166 39596
rect 102594 39584 102600 39596
rect 102652 39584 102658 39636
rect 103330 39584 103336 39636
rect 103388 39624 103394 39636
rect 116394 39624 116400 39636
rect 103388 39596 116400 39624
rect 103388 39584 103394 39596
rect 116394 39584 116400 39596
rect 116452 39584 116458 39636
rect 118602 39584 118608 39636
rect 118660 39624 118666 39636
rect 127526 39624 127532 39636
rect 118660 39596 127532 39624
rect 118660 39584 118666 39596
rect 127526 39584 127532 39596
rect 127584 39584 127590 39636
rect 129642 39584 129648 39636
rect 129700 39624 129706 39636
rect 136174 39624 136180 39636
rect 129700 39596 136180 39624
rect 129700 39584 129706 39596
rect 136174 39584 136180 39596
rect 136232 39584 136238 39636
rect 247310 39584 247316 39636
rect 247368 39624 247374 39636
rect 248966 39624 248972 39636
rect 247368 39596 248972 39624
rect 247368 39584 247374 39596
rect 248966 39584 248972 39596
rect 249024 39584 249030 39636
rect 262766 39584 262772 39636
rect 262824 39624 262830 39636
rect 287698 39624 287704 39636
rect 262824 39596 287704 39624
rect 262824 39584 262830 39596
rect 287698 39584 287704 39596
rect 287756 39584 287762 39636
rect 289538 39584 289544 39636
rect 289596 39624 289602 39636
rect 338758 39624 338764 39636
rect 289596 39596 338764 39624
rect 289596 39584 289602 39596
rect 338758 39584 338764 39596
rect 338816 39584 338822 39636
rect 346394 39584 346400 39636
rect 346452 39624 346458 39636
rect 395338 39624 395344 39636
rect 346452 39596 395344 39624
rect 346452 39584 346458 39596
rect 395338 39584 395344 39596
rect 395396 39584 395402 39636
rect 397178 39584 397184 39636
rect 397236 39624 397242 39636
rect 403069 39627 403127 39633
rect 403069 39624 403081 39627
rect 397236 39596 403081 39624
rect 397236 39584 397242 39596
rect 403069 39593 403081 39596
rect 403115 39593 403127 39627
rect 503714 39624 503720 39636
rect 403069 39587 403127 39593
rect 414308 39596 503720 39624
rect 13722 39516 13728 39568
rect 13780 39556 13786 39568
rect 51718 39556 51724 39568
rect 13780 39528 51724 39556
rect 13780 39516 13786 39528
rect 51718 39516 51724 39528
rect 51776 39516 51782 39568
rect 56502 39516 56508 39568
rect 56560 39556 56566 39568
rect 82814 39556 82820 39568
rect 56560 39528 82820 39556
rect 56560 39516 56566 39528
rect 82814 39516 82820 39528
rect 82872 39516 82878 39568
rect 86770 39516 86776 39568
rect 86828 39556 86834 39568
rect 105170 39556 105176 39568
rect 86828 39528 105176 39556
rect 86828 39516 86834 39528
rect 105170 39516 105176 39528
rect 105228 39516 105234 39568
rect 106182 39516 106188 39568
rect 106240 39556 106246 39568
rect 118970 39556 118976 39568
rect 106240 39528 118976 39556
rect 106240 39516 106246 39528
rect 118970 39516 118976 39528
rect 119028 39516 119034 39568
rect 121362 39516 121368 39568
rect 121420 39556 121426 39568
rect 130102 39556 130108 39568
rect 121420 39528 130108 39556
rect 121420 39516 121426 39528
rect 130102 39516 130108 39528
rect 130160 39516 130166 39568
rect 132402 39516 132408 39568
rect 132460 39556 132466 39568
rect 138014 39556 138020 39568
rect 132460 39528 138020 39556
rect 132460 39516 132466 39528
rect 138014 39516 138020 39528
rect 138072 39516 138078 39568
rect 224126 39516 224132 39568
rect 224184 39556 224190 39568
rect 244918 39556 244924 39568
rect 224184 39528 244924 39556
rect 224184 39516 224190 39528
rect 244918 39516 244924 39528
rect 244976 39516 244982 39568
rect 256786 39516 256792 39568
rect 256844 39556 256850 39568
rect 293954 39556 293960 39568
rect 256844 39528 293960 39556
rect 256844 39516 256850 39528
rect 293954 39516 293960 39528
rect 294012 39516 294018 39568
rect 307662 39516 307668 39568
rect 307720 39556 307726 39568
rect 356606 39556 356612 39568
rect 307720 39528 356612 39556
rect 307720 39516 307726 39528
rect 356606 39516 356612 39528
rect 356664 39516 356670 39568
rect 364518 39516 364524 39568
rect 364576 39556 364582 39568
rect 413278 39556 413284 39568
rect 364576 39528 413284 39556
rect 364576 39516 364582 39528
rect 413278 39516 413284 39528
rect 413336 39516 413342 39568
rect 6822 39448 6828 39500
rect 6880 39488 6886 39500
rect 46566 39488 46572 39500
rect 6880 39460 46572 39488
rect 6880 39448 6886 39460
rect 46566 39448 46572 39460
rect 46624 39448 46630 39500
rect 53650 39448 53656 39500
rect 53708 39488 53714 39500
rect 80146 39488 80152 39500
rect 53708 39460 80152 39488
rect 53708 39448 53714 39460
rect 80146 39448 80152 39460
rect 80204 39448 80210 39500
rect 81342 39448 81348 39500
rect 81400 39488 81406 39500
rect 100846 39488 100852 39500
rect 81400 39460 100852 39488
rect 81400 39448 81406 39460
rect 100846 39448 100852 39460
rect 100904 39448 100910 39500
rect 103422 39448 103428 39500
rect 103480 39488 103486 39500
rect 117314 39488 117320 39500
rect 103480 39460 117320 39488
rect 103480 39448 103486 39460
rect 117314 39448 117320 39460
rect 117372 39448 117378 39500
rect 119890 39448 119896 39500
rect 119948 39488 119954 39500
rect 129274 39488 129280 39500
rect 119948 39460 129280 39488
rect 119948 39448 119954 39460
rect 129274 39448 129280 39460
rect 129332 39448 129338 39500
rect 131022 39448 131028 39500
rect 131080 39488 131086 39500
rect 137002 39488 137008 39500
rect 131080 39460 137008 39488
rect 131080 39448 131086 39460
rect 137002 39448 137008 39460
rect 137060 39448 137066 39500
rect 218974 39448 218980 39500
rect 219032 39488 219038 39500
rect 224218 39488 224224 39500
rect 219032 39460 224224 39488
rect 219032 39448 219038 39460
rect 224218 39448 224224 39460
rect 224276 39448 224282 39500
rect 237006 39448 237012 39500
rect 237064 39488 237070 39500
rect 267090 39488 267096 39500
rect 237064 39460 267096 39488
rect 237064 39448 237070 39460
rect 267090 39448 267096 39460
rect 267148 39448 267154 39500
rect 273162 39448 273168 39500
rect 273220 39488 273226 39500
rect 282178 39488 282184 39500
rect 273220 39460 282184 39488
rect 273220 39448 273226 39460
rect 282178 39448 282184 39460
rect 282236 39448 282242 39500
rect 293862 39448 293868 39500
rect 293920 39488 293926 39500
rect 345014 39488 345020 39500
rect 293920 39460 345020 39488
rect 293920 39448 293926 39460
rect 345014 39448 345020 39460
rect 345072 39448 345078 39500
rect 359274 39448 359280 39500
rect 359332 39488 359338 39500
rect 411898 39488 411904 39500
rect 359332 39460 411904 39488
rect 359332 39448 359338 39460
rect 411898 39448 411904 39460
rect 411956 39448 411962 39500
rect 9582 39380 9588 39432
rect 9640 39420 9646 39432
rect 48314 39420 48320 39432
rect 9640 39392 48320 39420
rect 9640 39380 9646 39392
rect 48314 39380 48320 39392
rect 48372 39380 48378 39432
rect 49602 39380 49608 39432
rect 49660 39420 49666 39432
rect 77570 39420 77576 39432
rect 49660 39392 77576 39420
rect 49660 39380 49666 39392
rect 77570 39380 77576 39392
rect 77628 39380 77634 39432
rect 78490 39380 78496 39432
rect 78548 39420 78554 39432
rect 98270 39420 98276 39432
rect 78548 39392 98276 39420
rect 78548 39380 78554 39392
rect 98270 39380 98276 39392
rect 98328 39380 98334 39432
rect 99282 39380 99288 39432
rect 99340 39420 99346 39432
rect 113726 39420 113732 39432
rect 99340 39392 113732 39420
rect 99340 39380 99346 39392
rect 113726 39380 113732 39392
rect 113784 39380 113790 39432
rect 115842 39380 115848 39432
rect 115900 39420 115906 39432
rect 125870 39420 125876 39432
rect 115900 39392 125876 39420
rect 115900 39380 115906 39392
rect 125870 39380 125876 39392
rect 125928 39380 125934 39432
rect 229278 39380 229284 39432
rect 229336 39420 229342 39432
rect 255866 39420 255872 39432
rect 229336 39392 255872 39420
rect 229336 39380 229342 39392
rect 255866 39380 255872 39392
rect 255924 39380 255930 39432
rect 267182 39380 267188 39432
rect 267240 39420 267246 39432
rect 307754 39420 307760 39432
rect 267240 39392 307760 39420
rect 267240 39380 267246 39392
rect 307754 39380 307760 39392
rect 307812 39380 307818 39432
rect 315390 39380 315396 39432
rect 315448 39420 315454 39432
rect 370406 39420 370412 39432
rect 315448 39392 370412 39420
rect 315448 39380 315454 39392
rect 370406 39380 370412 39392
rect 370464 39380 370470 39432
rect 379974 39380 379980 39432
rect 380032 39420 380038 39432
rect 388438 39420 388444 39432
rect 380032 39392 388444 39420
rect 380032 39380 380038 39392
rect 388438 39380 388444 39392
rect 388496 39380 388502 39432
rect 409230 39380 409236 39432
rect 409288 39420 409294 39432
rect 414308 39420 414336 39596
rect 503714 39584 503720 39596
rect 503772 39584 503778 39636
rect 414382 39516 414388 39568
rect 414440 39556 414446 39568
rect 510614 39556 510620 39568
rect 414440 39528 510620 39556
rect 414440 39516 414446 39528
rect 510614 39516 510620 39528
rect 510672 39516 510678 39568
rect 512638 39488 512644 39500
rect 427096 39460 512644 39488
rect 427096 39420 427124 39460
rect 512638 39448 512644 39460
rect 512696 39448 512702 39500
rect 522298 39420 522304 39432
rect 409288 39392 414336 39420
rect 422266 39392 427124 39420
rect 431926 39392 522304 39420
rect 409288 39380 409294 39392
rect 4062 39312 4068 39364
rect 4120 39352 4126 39364
rect 44910 39352 44916 39364
rect 4120 39324 44916 39352
rect 4120 39312 4126 39324
rect 44910 39312 44916 39324
rect 44968 39312 44974 39364
rect 45462 39312 45468 39364
rect 45520 39352 45526 39364
rect 74994 39352 75000 39364
rect 45520 39324 75000 39352
rect 45520 39312 45526 39324
rect 74994 39312 75000 39324
rect 75052 39312 75058 39364
rect 75822 39312 75828 39364
rect 75880 39352 75886 39364
rect 96614 39352 96620 39364
rect 75880 39324 96620 39352
rect 75880 39312 75886 39324
rect 96614 39312 96620 39324
rect 96672 39312 96678 39364
rect 97902 39312 97908 39364
rect 97960 39352 97966 39364
rect 112898 39352 112904 39364
rect 97960 39324 112904 39352
rect 97960 39312 97966 39324
rect 112898 39312 112904 39324
rect 112956 39312 112962 39364
rect 113082 39312 113088 39364
rect 113140 39352 113146 39364
rect 124214 39352 124220 39364
rect 113140 39324 124220 39352
rect 113140 39312 113146 39324
rect 124214 39312 124220 39324
rect 124272 39312 124278 39364
rect 128170 39312 128176 39364
rect 128228 39352 128234 39364
rect 135254 39352 135260 39364
rect 128228 39324 135260 39352
rect 128228 39312 128234 39324
rect 135254 39312 135260 39324
rect 135312 39312 135318 39364
rect 216306 39312 216312 39364
rect 216364 39352 216370 39364
rect 238018 39352 238024 39364
rect 216364 39324 238024 39352
rect 216364 39312 216370 39324
rect 238018 39312 238024 39324
rect 238076 39312 238082 39364
rect 246482 39312 246488 39364
rect 246540 39352 246546 39364
rect 280246 39352 280252 39364
rect 246540 39324 280252 39352
rect 246540 39312 246546 39324
rect 280246 39312 280252 39324
rect 280304 39312 280310 39364
rect 282638 39312 282644 39364
rect 282696 39352 282702 39364
rect 329926 39352 329932 39364
rect 282696 39324 329932 39352
rect 282696 39312 282702 39324
rect 329926 39312 329932 39324
rect 329984 39312 329990 39364
rect 393958 39352 393964 39364
rect 335326 39324 393964 39352
rect 31662 39244 31668 39296
rect 31720 39284 31726 39296
rect 64690 39284 64696 39296
rect 31720 39256 64696 39284
rect 31720 39244 31726 39256
rect 64690 39244 64696 39256
rect 64748 39244 64754 39296
rect 70302 39244 70308 39296
rect 70360 39284 70366 39296
rect 93118 39284 93124 39296
rect 70360 39256 93124 39284
rect 70360 39244 70366 39256
rect 93118 39244 93124 39256
rect 93176 39244 93182 39296
rect 95142 39244 95148 39296
rect 95200 39284 95206 39296
rect 110414 39284 110420 39296
rect 95200 39256 110420 39284
rect 95200 39244 95206 39256
rect 110414 39244 110420 39256
rect 110472 39244 110478 39296
rect 117222 39244 117228 39296
rect 117280 39284 117286 39296
rect 126698 39284 126704 39296
rect 117280 39256 126704 39284
rect 117280 39244 117286 39256
rect 126698 39244 126704 39256
rect 126756 39244 126762 39296
rect 258534 39244 258540 39296
rect 258592 39284 258598 39296
rect 268378 39284 268384 39296
rect 258592 39256 268384 39284
rect 258592 39244 258598 39256
rect 268378 39244 268384 39256
rect 268436 39244 268442 39296
rect 282181 39287 282239 39293
rect 282181 39253 282193 39287
rect 282227 39284 282239 39287
rect 289078 39284 289084 39296
rect 282227 39256 289084 39284
rect 282227 39253 282239 39256
rect 282181 39247 282239 39253
rect 289078 39244 289084 39256
rect 289136 39244 289142 39296
rect 294690 39244 294696 39296
rect 294748 39284 294754 39296
rect 307018 39284 307024 39296
rect 294748 39256 307024 39284
rect 294748 39244 294754 39256
rect 307018 39244 307024 39256
rect 307076 39244 307082 39296
rect 311986 39244 311992 39296
rect 312044 39284 312050 39296
rect 324958 39284 324964 39296
rect 312044 39256 324964 39284
rect 312044 39244 312050 39256
rect 324958 39244 324964 39256
rect 325016 39244 325022 39296
rect 330846 39244 330852 39296
rect 330904 39284 330910 39296
rect 335326 39284 335354 39324
rect 393958 39312 393964 39324
rect 394016 39312 394022 39364
rect 416130 39312 416136 39364
rect 416188 39352 416194 39364
rect 422266 39352 422294 39392
rect 416188 39324 422294 39352
rect 416188 39312 416194 39324
rect 423858 39312 423864 39364
rect 423916 39352 423922 39364
rect 431926 39352 431954 39392
rect 522298 39380 522304 39392
rect 522356 39380 522362 39432
rect 423916 39324 431954 39352
rect 423916 39312 423922 39324
rect 434254 39312 434260 39364
rect 434312 39352 434318 39364
rect 437290 39352 437296 39364
rect 434312 39324 437296 39352
rect 434312 39312 434318 39324
rect 437290 39312 437296 39324
rect 437348 39312 437354 39364
rect 441982 39312 441988 39364
rect 442040 39352 442046 39364
rect 444190 39352 444196 39364
rect 442040 39324 444196 39352
rect 442040 39312 442046 39324
rect 444190 39312 444196 39324
rect 444248 39312 444254 39364
rect 462682 39312 462688 39364
rect 462740 39352 462746 39364
rect 574738 39352 574744 39364
rect 462740 39324 574744 39352
rect 462740 39312 462746 39324
rect 574738 39312 574744 39324
rect 574796 39312 574802 39364
rect 330904 39256 335354 39284
rect 330904 39244 330910 39256
rect 387702 39244 387708 39296
rect 387760 39284 387766 39296
rect 473354 39284 473360 39296
rect 387760 39256 473360 39284
rect 387760 39244 387766 39256
rect 473354 39244 473360 39256
rect 473412 39244 473418 39296
rect 33042 39176 33048 39228
rect 33100 39216 33106 39228
rect 65518 39216 65524 39228
rect 33100 39188 65524 39216
rect 33100 39176 33106 39188
rect 65518 39176 65524 39188
rect 65576 39176 65582 39228
rect 71682 39176 71688 39228
rect 71740 39216 71746 39228
rect 93946 39216 93952 39228
rect 71740 39188 93952 39216
rect 71740 39176 71746 39188
rect 93946 39176 93952 39188
rect 94004 39176 94010 39228
rect 96522 39176 96528 39228
rect 96580 39216 96586 39228
rect 112070 39216 112076 39228
rect 96580 39188 112076 39216
rect 96580 39176 96586 39188
rect 112070 39176 112076 39188
rect 112128 39176 112134 39228
rect 114462 39176 114468 39228
rect 114520 39216 114526 39228
rect 124950 39216 124956 39228
rect 114520 39188 124956 39216
rect 114520 39176 114526 39188
rect 124950 39176 124956 39188
rect 125008 39176 125014 39228
rect 404998 39176 405004 39228
rect 405056 39216 405062 39228
rect 489178 39216 489184 39228
rect 405056 39188 489184 39216
rect 405056 39176 405062 39188
rect 489178 39176 489184 39188
rect 489236 39176 489242 39228
rect 38562 39108 38568 39160
rect 38620 39148 38626 39160
rect 69842 39148 69848 39160
rect 38620 39120 69848 39148
rect 38620 39108 38626 39120
rect 69842 39108 69848 39120
rect 69900 39108 69906 39160
rect 74442 39108 74448 39160
rect 74500 39148 74506 39160
rect 95694 39148 95700 39160
rect 74500 39120 95700 39148
rect 74500 39108 74506 39120
rect 95694 39108 95700 39120
rect 95752 39108 95758 39160
rect 100662 39108 100668 39160
rect 100720 39148 100726 39160
rect 114646 39148 114652 39160
rect 100720 39120 114652 39148
rect 100720 39108 100726 39120
rect 114646 39108 114652 39120
rect 114704 39108 114710 39160
rect 392026 39108 392032 39160
rect 392084 39148 392090 39160
rect 475378 39148 475384 39160
rect 392084 39120 475384 39148
rect 392084 39108 392090 39120
rect 475378 39108 475384 39120
rect 475436 39108 475442 39160
rect 35802 39040 35808 39092
rect 35860 39080 35866 39092
rect 67266 39080 67272 39092
rect 35860 39052 67272 39080
rect 35860 39040 35866 39052
rect 67266 39040 67272 39052
rect 67324 39040 67330 39092
rect 68922 39040 68928 39092
rect 68980 39080 68986 39092
rect 91094 39080 91100 39092
rect 68980 39052 91100 39080
rect 68980 39040 68986 39052
rect 91094 39040 91100 39052
rect 91152 39040 91158 39092
rect 92382 39040 92388 39092
rect 92440 39080 92446 39092
rect 108574 39080 108580 39092
rect 92440 39052 108580 39080
rect 92440 39040 92446 39052
rect 108574 39040 108580 39052
rect 108632 39040 108638 39092
rect 136542 39040 136548 39092
rect 136600 39080 136606 39092
rect 141326 39080 141332 39092
rect 136600 39052 141332 39080
rect 136600 39040 136606 39052
rect 141326 39040 141332 39052
rect 141384 39040 141390 39092
rect 239582 39040 239588 39092
rect 239640 39080 239646 39092
rect 242158 39080 242164 39092
rect 239640 39052 242164 39080
rect 239640 39040 239646 39052
rect 242158 39040 242164 39052
rect 242216 39040 242222 39092
rect 410150 39040 410156 39092
rect 410208 39080 410214 39092
rect 467098 39080 467104 39092
rect 410208 39052 467104 39080
rect 410208 39040 410214 39052
rect 467098 39040 467104 39052
rect 467156 39040 467162 39092
rect 39942 38972 39948 39024
rect 40000 39012 40006 39024
rect 70670 39012 70676 39024
rect 40000 38984 70676 39012
rect 40000 38972 40006 38984
rect 70670 38972 70676 38984
rect 70728 38972 70734 39024
rect 73062 38972 73068 39024
rect 73120 39012 73126 39024
rect 94866 39012 94872 39024
rect 73120 38984 94872 39012
rect 73120 38972 73126 38984
rect 94866 38972 94872 38984
rect 94924 38972 94930 39024
rect 102042 38972 102048 39024
rect 102100 39012 102106 39024
rect 115474 39012 115480 39024
rect 102100 38984 115480 39012
rect 102100 38972 102106 38984
rect 115474 38972 115480 38984
rect 115532 38972 115538 39024
rect 139302 38972 139308 39024
rect 139360 39012 139366 39024
rect 143074 39012 143080 39024
rect 139360 38984 143080 39012
rect 139360 38972 139366 38984
rect 143074 38972 143080 38984
rect 143132 38972 143138 39024
rect 143442 38972 143448 39024
rect 143500 39012 143506 39024
rect 145650 39012 145656 39024
rect 143500 38984 145656 39012
rect 143500 38972 143506 38984
rect 145650 38972 145656 38984
rect 145708 38972 145714 39024
rect 146202 38972 146208 39024
rect 146260 39012 146266 39024
rect 148226 39012 148232 39024
rect 146260 38984 148232 39012
rect 146260 38972 146266 38984
rect 148226 38972 148232 38984
rect 148284 38972 148290 39024
rect 148962 38972 148968 39024
rect 149020 39012 149026 39024
rect 149974 39012 149980 39024
rect 149020 38984 149980 39012
rect 149020 38972 149026 38984
rect 149974 38972 149980 38984
rect 150032 38972 150038 39024
rect 151814 38972 151820 39024
rect 151872 39012 151878 39024
rect 152550 39012 152556 39024
rect 151872 38984 152556 39012
rect 151872 38972 151878 38984
rect 152550 38972 152556 38984
rect 152608 38972 152614 39024
rect 157794 38972 157800 39024
rect 157852 39012 157858 39024
rect 158530 39012 158536 39024
rect 157852 38984 158536 39012
rect 157852 38972 157858 38984
rect 158530 38972 158536 38984
rect 158588 38972 158594 39024
rect 159542 38972 159548 39024
rect 159600 39012 159606 39024
rect 160002 39012 160008 39024
rect 159600 38984 160008 39012
rect 159600 38972 159606 38984
rect 160002 38972 160008 38984
rect 160060 38972 160066 39024
rect 162118 38972 162124 39024
rect 162176 39012 162182 39024
rect 162762 39012 162768 39024
rect 162176 38984 162768 39012
rect 162176 38972 162182 38984
rect 162762 38972 162768 38984
rect 162820 38972 162826 39024
rect 162946 38972 162952 39024
rect 163004 39012 163010 39024
rect 165706 39012 165712 39024
rect 163004 38984 165712 39012
rect 163004 38972 163010 38984
rect 165706 38972 165712 38984
rect 165764 38972 165770 39024
rect 166350 38972 166356 39024
rect 166408 39012 166414 39024
rect 166902 39012 166908 39024
rect 166408 38984 166908 39012
rect 166408 38972 166414 38984
rect 166902 38972 166908 38984
rect 166960 38972 166966 39024
rect 167270 38972 167276 39024
rect 167328 39012 167334 39024
rect 168282 39012 168288 39024
rect 167328 38984 168288 39012
rect 167328 38972 167334 38984
rect 168282 38972 168288 38984
rect 168340 38972 168346 39024
rect 169018 38972 169024 39024
rect 169076 39012 169082 39024
rect 169662 39012 169668 39024
rect 169076 38984 169668 39012
rect 169076 38972 169082 38984
rect 169662 38972 169668 38984
rect 169720 38972 169726 39024
rect 169846 38972 169852 39024
rect 169904 39012 169910 39024
rect 170950 39012 170956 39024
rect 169904 38984 170956 39012
rect 169904 38972 169910 38984
rect 170950 38972 170956 38984
rect 171008 38972 171014 39024
rect 171594 38972 171600 39024
rect 171652 39012 171658 39024
rect 172330 39012 172336 39024
rect 171652 38984 172336 39012
rect 171652 38972 171658 38984
rect 172330 38972 172336 38984
rect 172388 38972 172394 39024
rect 173250 38972 173256 39024
rect 173308 39012 173314 39024
rect 173802 39012 173808 39024
rect 173308 38984 173808 39012
rect 173308 38972 173314 38984
rect 173802 38972 173808 38984
rect 173860 38972 173866 39024
rect 175826 38972 175832 39024
rect 175884 39012 175890 39024
rect 176562 39012 176568 39024
rect 175884 38984 176568 39012
rect 175884 38972 175890 38984
rect 176562 38972 176568 38984
rect 176620 38972 176626 39024
rect 178494 38972 178500 39024
rect 178552 39012 178558 39024
rect 179322 39012 179328 39024
rect 178552 38984 179328 39012
rect 178552 38972 178558 38984
rect 179322 38972 179328 38984
rect 179380 38972 179386 39024
rect 180150 38972 180156 39024
rect 180208 39012 180214 39024
rect 180702 39012 180708 39024
rect 180208 38984 180708 39012
rect 180208 38972 180214 38984
rect 180702 38972 180708 38984
rect 180760 38972 180766 39024
rect 181070 38972 181076 39024
rect 181128 39012 181134 39024
rect 182082 39012 182088 39024
rect 181128 38984 182088 39012
rect 181128 38972 181134 38984
rect 182082 38972 182088 38984
rect 182140 38972 182146 39024
rect 182726 38972 182732 39024
rect 182784 39012 182790 39024
rect 183462 39012 183468 39024
rect 182784 38984 183468 39012
rect 182784 38972 182790 38984
rect 183462 38972 183468 38984
rect 183520 38972 183526 39024
rect 183646 38972 183652 39024
rect 183704 39012 183710 39024
rect 184842 39012 184848 39024
rect 183704 38984 184848 39012
rect 183704 38972 183710 38984
rect 184842 38972 184848 38984
rect 184900 38972 184906 39024
rect 185302 38972 185308 39024
rect 185360 39012 185366 39024
rect 186130 39012 186136 39024
rect 185360 38984 186136 39012
rect 185360 38972 185366 38984
rect 186130 38972 186136 38984
rect 186188 38972 186194 39024
rect 187050 38972 187056 39024
rect 187108 39012 187114 39024
rect 187602 39012 187608 39024
rect 187108 38984 187608 39012
rect 187108 38972 187114 38984
rect 187602 38972 187608 38984
rect 187660 38972 187666 39024
rect 187970 38972 187976 39024
rect 188028 39012 188034 39024
rect 188890 39012 188896 39024
rect 188028 38984 188896 39012
rect 188028 38972 188034 38984
rect 188890 38972 188896 38984
rect 188948 38972 188954 39024
rect 189626 38972 189632 39024
rect 189684 39012 189690 39024
rect 190362 39012 190368 39024
rect 189684 38984 190368 39012
rect 189684 38972 189690 38984
rect 190362 38972 190368 38984
rect 190420 38972 190426 39024
rect 190546 38972 190552 39024
rect 190604 39012 190610 39024
rect 191650 39012 191656 39024
rect 190604 38984 191656 39012
rect 190604 38972 190610 38984
rect 191650 38972 191656 38984
rect 191708 38972 191714 39024
rect 192202 38972 192208 39024
rect 192260 39012 192266 39024
rect 193122 39012 193128 39024
rect 192260 38984 193128 39012
rect 192260 38972 192266 38984
rect 193122 38972 193128 38984
rect 193180 38972 193186 39024
rect 193950 38972 193956 39024
rect 194008 39012 194014 39024
rect 194502 39012 194508 39024
rect 194008 38984 194508 39012
rect 194008 38972 194014 38984
rect 194502 38972 194508 38984
rect 194560 38972 194566 39024
rect 194778 38972 194784 39024
rect 194836 39012 194842 39024
rect 195790 39012 195796 39024
rect 194836 38984 195796 39012
rect 194836 38972 194842 38984
rect 195790 38972 195796 38984
rect 195848 38972 195854 39024
rect 196526 38972 196532 39024
rect 196584 39012 196590 39024
rect 197262 39012 197268 39024
rect 196584 38984 197268 39012
rect 196584 38972 196590 38984
rect 197262 38972 197268 38984
rect 197320 38972 197326 39024
rect 197354 38972 197360 39024
rect 197412 39012 197418 39024
rect 198642 39012 198648 39024
rect 197412 38984 198648 39012
rect 197412 38972 197418 38984
rect 198642 38972 198648 38984
rect 198700 38972 198706 39024
rect 199102 38972 199108 39024
rect 199160 39012 199166 39024
rect 200022 39012 200028 39024
rect 199160 38984 200028 39012
rect 199160 38972 199166 38984
rect 200022 38972 200028 38984
rect 200080 38972 200086 39024
rect 200850 38972 200856 39024
rect 200908 39012 200914 39024
rect 201402 39012 201408 39024
rect 200908 38984 201408 39012
rect 200908 38972 200914 38984
rect 201402 38972 201408 38984
rect 201460 38972 201466 39024
rect 201678 38972 201684 39024
rect 201736 39012 201742 39024
rect 202782 39012 202788 39024
rect 201736 38984 202788 39012
rect 201736 38972 201742 38984
rect 202782 38972 202788 38984
rect 202840 38972 202846 39024
rect 203426 38972 203432 39024
rect 203484 39012 203490 39024
rect 204162 39012 204168 39024
rect 203484 38984 204168 39012
rect 203484 38972 203490 38984
rect 204162 38972 204168 38984
rect 204220 38972 204226 39024
rect 206002 38972 206008 39024
rect 206060 39012 206066 39024
rect 206830 39012 206836 39024
rect 206060 38984 206836 39012
rect 206060 38972 206066 38984
rect 206830 38972 206836 38984
rect 206888 38972 206894 39024
rect 207750 38972 207756 39024
rect 207808 39012 207814 39024
rect 208302 39012 208308 39024
rect 207808 38984 208308 39012
rect 207808 38972 207814 38984
rect 208302 38972 208308 38984
rect 208360 38972 208366 39024
rect 208578 38972 208584 39024
rect 208636 39012 208642 39024
rect 209590 39012 209596 39024
rect 208636 38984 209596 39012
rect 208636 38972 208642 38984
rect 209590 38972 209596 38984
rect 209648 38972 209654 39024
rect 210326 38972 210332 39024
rect 210384 39012 210390 39024
rect 211062 39012 211068 39024
rect 210384 38984 211068 39012
rect 210384 38972 210390 38984
rect 211062 38972 211068 38984
rect 211120 38972 211126 39024
rect 211154 38972 211160 39024
rect 211212 39012 211218 39024
rect 212350 39012 212356 39024
rect 211212 38984 212356 39012
rect 211212 38972 211218 38984
rect 212350 38972 212356 38984
rect 212408 38972 212414 39024
rect 212902 38972 212908 39024
rect 212960 39012 212966 39024
rect 213822 39012 213828 39024
rect 212960 38984 213828 39012
rect 212960 38972 212966 38984
rect 213822 38972 213828 38984
rect 213880 38972 213886 39024
rect 214650 38972 214656 39024
rect 214708 39012 214714 39024
rect 215202 39012 215208 39024
rect 214708 38984 215208 39012
rect 214708 38972 214714 38984
rect 215202 38972 215208 38984
rect 215260 38972 215266 39024
rect 215478 38972 215484 39024
rect 215536 39012 215542 39024
rect 216582 39012 216588 39024
rect 215536 38984 216588 39012
rect 215536 38972 215542 38984
rect 216582 38972 216588 38984
rect 216640 38972 216646 39024
rect 217226 38972 217232 39024
rect 217284 39012 217290 39024
rect 217962 39012 217968 39024
rect 217284 38984 217968 39012
rect 217284 38972 217290 38984
rect 217962 38972 217968 38984
rect 218020 38972 218026 39024
rect 218054 38972 218060 39024
rect 218112 39012 218118 39024
rect 219342 39012 219348 39024
rect 218112 38984 219348 39012
rect 218112 38972 218118 38984
rect 219342 38972 219348 38984
rect 219400 38972 219406 39024
rect 219802 38972 219808 39024
rect 219860 39012 219866 39024
rect 220722 39012 220728 39024
rect 219860 38984 220728 39012
rect 219860 38972 219866 38984
rect 220722 38972 220728 38984
rect 220780 38972 220786 39024
rect 224954 38972 224960 39024
rect 225012 39012 225018 39024
rect 226242 39012 226248 39024
rect 225012 38984 226248 39012
rect 225012 38972 225018 38984
rect 226242 38972 226248 38984
rect 226300 38972 226306 39024
rect 226702 38972 226708 39024
rect 226760 39012 226766 39024
rect 227530 39012 227536 39024
rect 226760 38984 227536 39012
rect 226760 38972 226766 38984
rect 227530 38972 227536 38984
rect 227588 38972 227594 39024
rect 228358 38972 228364 39024
rect 228416 39012 228422 39024
rect 229002 39012 229008 39024
rect 228416 38984 229008 39012
rect 228416 38972 228422 38984
rect 229002 38972 229008 38984
rect 229060 38972 229066 39024
rect 231026 38972 231032 39024
rect 231084 39012 231090 39024
rect 231762 39012 231768 39024
rect 231084 38984 231768 39012
rect 231084 38972 231090 38984
rect 231762 38972 231768 38984
rect 231820 38972 231826 39024
rect 232682 38972 232688 39024
rect 232740 39012 232746 39024
rect 233142 39012 233148 39024
rect 232740 38984 233148 39012
rect 232740 38972 232746 38984
rect 233142 38972 233148 38984
rect 233200 38972 233206 39024
rect 235258 38972 235264 39024
rect 235316 39012 235322 39024
rect 235902 39012 235908 39024
rect 235316 38984 235908 39012
rect 235316 38972 235322 38984
rect 235902 38972 235908 38984
rect 235960 38972 235966 39024
rect 236178 38972 236184 39024
rect 236236 39012 236242 39024
rect 237282 39012 237288 39024
rect 236236 38984 237288 39012
rect 236236 38972 236242 38984
rect 237282 38972 237288 38984
rect 237340 38972 237346 39024
rect 237834 38972 237840 39024
rect 237892 39012 237898 39024
rect 238662 39012 238668 39024
rect 237892 38984 238668 39012
rect 237892 38972 237898 38984
rect 238662 38972 238668 38984
rect 238720 38972 238726 39024
rect 238754 38972 238760 39024
rect 238812 39012 238818 39024
rect 240042 39012 240048 39024
rect 238812 38984 240048 39012
rect 238812 38972 238818 38984
rect 240042 38972 240048 38984
rect 240100 38972 240106 39024
rect 240502 38972 240508 39024
rect 240560 39012 240566 39024
rect 241422 39012 241428 39024
rect 240560 38984 241428 39012
rect 240560 38972 240566 38984
rect 241422 38972 241428 38984
rect 241480 38972 241486 39024
rect 243078 38972 243084 39024
rect 243136 39012 243142 39024
rect 244182 39012 244188 39024
rect 243136 38984 244188 39012
rect 243136 38972 243142 38984
rect 244182 38972 244188 38984
rect 244240 38972 244246 39024
rect 245654 38972 245660 39024
rect 245712 39012 245718 39024
rect 246942 39012 246948 39024
rect 245712 38984 246948 39012
rect 245712 38972 245718 38984
rect 246942 38972 246948 38984
rect 247000 38972 247006 39024
rect 249058 38972 249064 39024
rect 249116 39012 249122 39024
rect 249702 39012 249708 39024
rect 249116 38984 249708 39012
rect 249116 38972 249122 38984
rect 249702 38972 249708 38984
rect 249760 38972 249766 39024
rect 249978 38972 249984 39024
rect 250036 39012 250042 39024
rect 250990 39012 250996 39024
rect 250036 38984 250996 39012
rect 250036 38972 250042 38984
rect 250990 38972 250996 38984
rect 251048 38972 251054 39024
rect 251634 38972 251640 39024
rect 251692 39012 251698 39024
rect 252462 39012 252468 39024
rect 251692 38984 252468 39012
rect 251692 38972 251698 38984
rect 252462 38972 252468 38984
rect 252520 38972 252526 39024
rect 253382 38972 253388 39024
rect 253440 39012 253446 39024
rect 253842 39012 253848 39024
rect 253440 38984 253848 39012
rect 253440 38972 253446 38984
rect 253842 38972 253848 38984
rect 253900 38972 253906 39024
rect 254210 38972 254216 39024
rect 254268 39012 254274 39024
rect 255222 39012 255228 39024
rect 254268 38984 255228 39012
rect 254268 38972 254274 38984
rect 255222 38972 255228 38984
rect 255280 38972 255286 39024
rect 255958 38972 255964 39024
rect 256016 39012 256022 39024
rect 256602 39012 256608 39024
rect 256016 38984 256608 39012
rect 256016 38972 256022 38984
rect 256602 38972 256608 38984
rect 256660 38972 256666 39024
rect 260282 38972 260288 39024
rect 260340 39012 260346 39024
rect 260742 39012 260748 39024
rect 260340 38984 260748 39012
rect 260340 38972 260346 38984
rect 260742 38972 260748 38984
rect 260800 38972 260806 39024
rect 261110 38972 261116 39024
rect 261168 39012 261174 39024
rect 262950 39012 262956 39024
rect 261168 38984 262956 39012
rect 261168 38972 261174 38984
rect 262950 38972 262956 38984
rect 263008 38972 263014 39024
rect 263686 38972 263692 39024
rect 263744 39012 263750 39024
rect 264790 39012 264796 39024
rect 263744 38984 264796 39012
rect 263744 38972 263750 38984
rect 264790 38972 264796 38984
rect 264848 38972 264854 39024
rect 265434 38972 265440 39024
rect 265492 39012 265498 39024
rect 266998 39012 267004 39024
rect 265492 38984 267004 39012
rect 265492 38972 265498 38984
rect 266998 38972 267004 38984
rect 267056 38972 267062 39024
rect 269758 38972 269764 39024
rect 269816 39012 269822 39024
rect 270402 39012 270408 39024
rect 269816 38984 270408 39012
rect 269816 38972 269822 38984
rect 270402 38972 270408 38984
rect 270460 38972 270466 39024
rect 270586 38972 270592 39024
rect 270644 39012 270650 39024
rect 271782 39012 271788 39024
rect 270644 38984 271788 39012
rect 270644 38972 270650 38984
rect 271782 38972 271788 38984
rect 271840 38972 271846 39024
rect 272334 38972 272340 39024
rect 272392 39012 272398 39024
rect 273162 39012 273168 39024
rect 272392 38984 273168 39012
rect 272392 38972 272398 38984
rect 273162 38972 273168 38984
rect 273220 38972 273226 39024
rect 274082 38972 274088 39024
rect 274140 39012 274146 39024
rect 274542 39012 274548 39024
rect 274140 38984 274548 39012
rect 274140 38972 274146 38984
rect 274542 38972 274548 38984
rect 274600 38972 274606 39024
rect 274910 38972 274916 39024
rect 274968 39012 274974 39024
rect 275922 39012 275928 39024
rect 274968 38984 275928 39012
rect 274968 38972 274974 38984
rect 275922 38972 275928 38984
rect 275980 38972 275986 39024
rect 276658 38972 276664 39024
rect 276716 39012 276722 39024
rect 277302 39012 277308 39024
rect 276716 38984 277308 39012
rect 276716 38972 276722 38984
rect 277302 38972 277308 38984
rect 277360 38972 277366 39024
rect 277486 38972 277492 39024
rect 277544 39012 277550 39024
rect 278682 39012 278688 39024
rect 277544 38984 278688 39012
rect 277544 38972 277550 38984
rect 278682 38972 278688 38984
rect 278740 38972 278746 39024
rect 279234 38972 279240 39024
rect 279292 39012 279298 39024
rect 280798 39012 280804 39024
rect 279292 38984 280804 39012
rect 279292 38972 279298 38984
rect 280798 38972 280804 38984
rect 280856 38972 280862 39024
rect 280982 38972 280988 39024
rect 281040 39012 281046 39024
rect 281442 39012 281448 39024
rect 281040 38984 281448 39012
rect 281040 38972 281046 38984
rect 281442 38972 281448 38984
rect 281500 38972 281506 39024
rect 286134 38972 286140 39024
rect 286192 39012 286198 39024
rect 286962 39012 286968 39024
rect 286192 38984 286968 39012
rect 286192 38972 286198 38984
rect 286962 38972 286968 38984
rect 287020 38972 287026 39024
rect 288710 38972 288716 39024
rect 288768 39012 288774 39024
rect 289722 39012 289728 39024
rect 288768 38984 289728 39012
rect 288768 38972 288774 38984
rect 289722 38972 289728 38984
rect 289780 38972 289786 39024
rect 290366 38972 290372 39024
rect 290424 39012 290430 39024
rect 291102 39012 291108 39024
rect 290424 38984 291108 39012
rect 290424 38972 290430 38984
rect 291102 38972 291108 38984
rect 291160 38972 291166 39024
rect 291286 38972 291292 39024
rect 291344 39012 291350 39024
rect 292482 39012 292488 39024
rect 291344 38984 292488 39012
rect 291344 38972 291350 38984
rect 292482 38972 292488 38984
rect 292540 38972 292546 39024
rect 293034 38972 293040 39024
rect 293092 39012 293098 39024
rect 293862 39012 293868 39024
rect 293092 38984 293868 39012
rect 293092 38972 293098 38984
rect 293862 38972 293868 38984
rect 293920 38972 293926 39024
rect 295610 38972 295616 39024
rect 295668 39012 295674 39024
rect 296622 39012 296628 39024
rect 295668 38984 296628 39012
rect 295668 38972 295674 38984
rect 296622 38972 296628 38984
rect 296680 38972 296686 39024
rect 298186 38972 298192 39024
rect 298244 39012 298250 39024
rect 299382 39012 299388 39024
rect 298244 38984 299388 39012
rect 298244 38972 298250 38984
rect 299382 38972 299388 38984
rect 299440 38972 299446 39024
rect 299842 38972 299848 39024
rect 299900 39012 299906 39024
rect 300670 39012 300676 39024
rect 299900 38984 300676 39012
rect 299900 38972 299906 38984
rect 300670 38972 300676 38984
rect 300728 38972 300734 39024
rect 302510 38972 302516 39024
rect 302568 39012 302574 39024
rect 303430 39012 303436 39024
rect 302568 38984 303436 39012
rect 302568 38972 302574 38984
rect 303430 38972 303436 38984
rect 303488 38972 303494 39024
rect 305086 38972 305092 39024
rect 305144 39012 305150 39024
rect 306190 39012 306196 39024
rect 305144 38984 306196 39012
rect 305144 38972 305150 38984
rect 306190 38972 306196 38984
rect 306248 38972 306254 39024
rect 306742 38972 306748 39024
rect 306800 39012 306806 39024
rect 307662 39012 307668 39024
rect 306800 38984 307668 39012
rect 306800 38972 306806 38984
rect 307662 38972 307668 38984
rect 307720 38972 307726 39024
rect 309318 38972 309324 39024
rect 309376 39012 309382 39024
rect 310422 39012 310428 39024
rect 309376 38984 310428 39012
rect 309376 38972 309382 38984
rect 310422 38972 310428 38984
rect 310480 38972 310486 39024
rect 311066 38972 311072 39024
rect 311124 39012 311130 39024
rect 311802 39012 311808 39024
rect 311124 38984 311808 39012
rect 311124 38972 311130 38984
rect 311802 38972 311808 38984
rect 311860 38972 311866 39024
rect 313642 38972 313648 39024
rect 313700 39012 313706 39024
rect 314562 39012 314568 39024
rect 313700 38984 314568 39012
rect 313700 38972 313706 38984
rect 314562 38972 314568 38984
rect 314620 38972 314626 39024
rect 316218 38972 316224 39024
rect 316276 39012 316282 39024
rect 317322 39012 317328 39024
rect 316276 38984 317328 39012
rect 316276 38972 316282 38984
rect 317322 38972 317328 38984
rect 317380 38972 317386 39024
rect 317966 38972 317972 39024
rect 318024 39012 318030 39024
rect 318702 39012 318708 39024
rect 318024 38984 318708 39012
rect 318024 38972 318030 38984
rect 318702 38972 318708 38984
rect 318760 38972 318766 39024
rect 318794 38972 318800 39024
rect 318852 39012 318858 39024
rect 320082 39012 320088 39024
rect 318852 38984 320088 39012
rect 318852 38972 318858 38984
rect 320082 38972 320088 38984
rect 320140 38972 320146 39024
rect 320542 38972 320548 39024
rect 320600 39012 320606 39024
rect 321370 39012 321376 39024
rect 320600 38984 321376 39012
rect 320600 38972 320606 38984
rect 321370 38972 321376 38984
rect 321428 38972 321434 39024
rect 323118 38972 323124 39024
rect 323176 39012 323182 39024
rect 324130 39012 324136 39024
rect 323176 38984 324136 39012
rect 323176 38972 323182 38984
rect 324130 38972 324136 38984
rect 324188 38972 324194 39024
rect 324866 38972 324872 39024
rect 324924 39012 324930 39024
rect 325602 39012 325608 39024
rect 324924 38984 325608 39012
rect 324924 38972 324930 38984
rect 325602 38972 325608 38984
rect 325660 38972 325666 39024
rect 329190 38972 329196 39024
rect 329248 39012 329254 39024
rect 329742 39012 329748 39024
rect 329248 38984 329748 39012
rect 329248 38972 329254 38984
rect 329742 38972 329748 38984
rect 329800 38972 329806 39024
rect 330018 38972 330024 39024
rect 330076 39012 330082 39024
rect 331122 39012 331128 39024
rect 330076 38984 331128 39012
rect 330076 38972 330082 38984
rect 331122 38972 331128 38984
rect 331180 38972 331186 39024
rect 331766 38972 331772 39024
rect 331824 39012 331830 39024
rect 332502 39012 332508 39024
rect 331824 38984 332508 39012
rect 331824 38972 331830 38984
rect 332502 38972 332508 38984
rect 332560 38972 332566 39024
rect 332594 38972 332600 39024
rect 332652 39012 332658 39024
rect 333882 39012 333888 39024
rect 332652 38984 333888 39012
rect 332652 38972 332658 38984
rect 333882 38972 333888 38984
rect 333940 38972 333946 39024
rect 334342 38972 334348 39024
rect 334400 39012 334406 39024
rect 335262 39012 335268 39024
rect 334400 38984 335268 39012
rect 334400 38972 334406 38984
rect 335262 38972 335268 38984
rect 335320 38972 335326 39024
rect 336090 38972 336096 39024
rect 336148 39012 336154 39024
rect 336642 39012 336648 39024
rect 336148 38984 336648 39012
rect 336148 38972 336154 38984
rect 336642 38972 336648 38984
rect 336700 38972 336706 39024
rect 336918 38972 336924 39024
rect 336976 39012 336982 39024
rect 338022 39012 338028 39024
rect 336976 38984 338028 39012
rect 336976 38972 336982 38984
rect 338022 38972 338028 38984
rect 338080 38972 338086 39024
rect 338666 38972 338672 39024
rect 338724 39012 338730 39024
rect 339402 39012 339408 39024
rect 338724 38984 339408 39012
rect 338724 38972 338730 38984
rect 339402 38972 339408 38984
rect 339460 38972 339466 39024
rect 339494 38972 339500 39024
rect 339552 39012 339558 39024
rect 340782 39012 340788 39024
rect 339552 38984 340788 39012
rect 339552 38972 339558 38984
rect 340782 38972 340788 38984
rect 340840 38972 340846 39024
rect 341242 38972 341248 39024
rect 341300 39012 341306 39024
rect 342070 39012 342076 39024
rect 341300 38984 342076 39012
rect 341300 38972 341306 38984
rect 342070 38972 342076 38984
rect 342128 38972 342134 39024
rect 342990 38972 342996 39024
rect 343048 39012 343054 39024
rect 343542 39012 343548 39024
rect 343048 38984 343548 39012
rect 343048 38972 343054 38984
rect 343542 38972 343548 38984
rect 343600 38972 343606 39024
rect 345566 38972 345572 39024
rect 345624 39012 345630 39024
rect 346302 39012 346308 39024
rect 345624 38984 346308 39012
rect 345624 38972 345630 38984
rect 346302 38972 346308 38984
rect 346360 38972 346366 39024
rect 347222 38972 347228 39024
rect 347280 39012 347286 39024
rect 347682 39012 347688 39024
rect 347280 38984 347688 39012
rect 347280 38972 347286 38984
rect 347682 38972 347688 38984
rect 347740 38972 347746 39024
rect 348142 38972 348148 39024
rect 348200 39012 348206 39024
rect 349062 39012 349068 39024
rect 348200 38984 349068 39012
rect 348200 38972 348206 38984
rect 349062 38972 349068 38984
rect 349120 38972 349126 39024
rect 349798 38972 349804 39024
rect 349856 39012 349862 39024
rect 350442 39012 350448 39024
rect 349856 38984 350448 39012
rect 349856 38972 349862 38984
rect 350442 38972 350448 38984
rect 350500 38972 350506 39024
rect 350718 38972 350724 39024
rect 350776 39012 350782 39024
rect 351822 39012 351828 39024
rect 350776 38984 351828 39012
rect 350776 38972 350782 38984
rect 351822 38972 351828 38984
rect 351880 38972 351886 39024
rect 352374 38972 352380 39024
rect 352432 39012 352438 39024
rect 353202 39012 353208 39024
rect 352432 38984 353208 39012
rect 352432 38972 352438 38984
rect 353202 38972 353208 38984
rect 353260 38972 353266 39024
rect 353294 38972 353300 39024
rect 353352 39012 353358 39024
rect 354582 39012 354588 39024
rect 353352 38984 354588 39012
rect 353352 38972 353358 38984
rect 354582 38972 354588 38984
rect 354640 38972 354646 39024
rect 355042 38972 355048 39024
rect 355100 39012 355106 39024
rect 355962 39012 355968 39024
rect 355100 38984 355968 39012
rect 355100 38972 355106 38984
rect 355962 38972 355968 38984
rect 356020 38972 356026 39024
rect 356698 38972 356704 39024
rect 356756 39012 356762 39024
rect 357342 39012 357348 39024
rect 356756 38984 357348 39012
rect 356756 38972 356762 38984
rect 357342 38972 357348 38984
rect 357400 38972 357406 39024
rect 357618 38972 357624 39024
rect 357676 39012 357682 39024
rect 358722 39012 358728 39024
rect 357676 38984 358728 39012
rect 357676 38972 357682 38984
rect 358722 38972 358728 38984
rect 358780 38972 358786 39024
rect 360194 38972 360200 39024
rect 360252 39012 360258 39024
rect 361482 39012 361488 39024
rect 360252 38984 361488 39012
rect 360252 38972 360258 38984
rect 361482 38972 361488 38984
rect 361540 38972 361546 39024
rect 363598 38972 363604 39024
rect 363656 39012 363662 39024
rect 364242 39012 364248 39024
rect 363656 38984 364248 39012
rect 363656 38972 363662 38984
rect 364242 38972 364248 38984
rect 364300 38972 364306 39024
rect 366174 38972 366180 39024
rect 366232 39012 366238 39024
rect 367002 39012 367008 39024
rect 366232 38984 367008 39012
rect 366232 38972 366238 38984
rect 367002 38972 367008 38984
rect 367060 38972 367066 39024
rect 367922 38972 367928 39024
rect 367980 39012 367986 39024
rect 368382 39012 368388 39024
rect 367980 38984 368388 39012
rect 367980 38972 367986 38984
rect 368382 38972 368388 38984
rect 368440 38972 368446 39024
rect 368750 38972 368756 39024
rect 368808 39012 368814 39024
rect 369762 39012 369768 39024
rect 368808 38984 369768 39012
rect 368808 38972 368814 38984
rect 369762 38972 369768 38984
rect 369820 38972 369826 39024
rect 370498 38972 370504 39024
rect 370556 39012 370562 39024
rect 371142 39012 371148 39024
rect 370556 38984 371148 39012
rect 370556 38972 370562 38984
rect 371142 38972 371148 38984
rect 371200 38972 371206 39024
rect 373074 38972 373080 39024
rect 373132 39012 373138 39024
rect 373902 39012 373908 39024
rect 373132 38984 373908 39012
rect 373132 38972 373138 38984
rect 373902 38972 373908 38984
rect 373960 38972 373966 39024
rect 373994 38972 374000 39024
rect 374052 39012 374058 39024
rect 375282 39012 375288 39024
rect 374052 38984 375288 39012
rect 374052 38972 374058 38984
rect 375282 38972 375288 38984
rect 375340 38972 375346 39024
rect 375650 38972 375656 39024
rect 375708 39012 375714 39024
rect 376662 39012 376668 39024
rect 375708 38984 376668 39012
rect 375708 38972 375714 38984
rect 376662 38972 376668 38984
rect 376720 38972 376726 39024
rect 377398 38972 377404 39024
rect 377456 39012 377462 39024
rect 378042 39012 378048 39024
rect 377456 38984 378048 39012
rect 377456 38972 377462 38984
rect 378042 38972 378048 38984
rect 378100 38972 378106 39024
rect 382550 38972 382556 39024
rect 382608 39012 382614 39024
rect 383470 39012 383476 39024
rect 382608 38984 383476 39012
rect 382608 38972 382614 38984
rect 383470 38972 383476 38984
rect 383528 38972 383534 39024
rect 384298 38972 384304 39024
rect 384356 39012 384362 39024
rect 384942 39012 384948 39024
rect 384356 38984 384948 39012
rect 384356 38972 384362 38984
rect 384942 38972 384948 38984
rect 385000 38972 385006 39024
rect 388622 38972 388628 39024
rect 388680 39012 388686 39024
rect 389082 39012 389088 39024
rect 388680 38984 389088 39012
rect 388680 38972 388686 38984
rect 389082 38972 389088 38984
rect 389140 38972 389146 39024
rect 389450 38972 389456 39024
rect 389508 39012 389514 39024
rect 390462 39012 390468 39024
rect 389508 38984 390468 39012
rect 389508 38972 389514 38984
rect 390462 38972 390468 38984
rect 390520 38972 390526 39024
rect 395522 38972 395528 39024
rect 395580 39012 395586 39024
rect 395982 39012 395988 39024
rect 395580 38984 395988 39012
rect 395580 38972 395586 38984
rect 395982 38972 395988 38984
rect 396040 38972 396046 39024
rect 396350 38972 396356 39024
rect 396408 39012 396414 39024
rect 397362 39012 397368 39024
rect 396408 38984 397368 39012
rect 396408 38972 396414 38984
rect 397362 38972 397368 38984
rect 397420 38972 397426 39024
rect 398098 38972 398104 39024
rect 398156 39012 398162 39024
rect 398742 39012 398748 39024
rect 398156 38984 398748 39012
rect 398156 38972 398162 38984
rect 398742 38972 398748 38984
rect 398800 38972 398806 39024
rect 400674 38972 400680 39024
rect 400732 39012 400738 39024
rect 401502 39012 401508 39024
rect 400732 38984 401508 39012
rect 400732 38972 400738 38984
rect 401502 38972 401508 38984
rect 401560 38972 401566 39024
rect 403250 38972 403256 39024
rect 403308 39012 403314 39024
rect 404262 39012 404268 39024
rect 403308 38984 404268 39012
rect 403308 38972 403314 38984
rect 404262 38972 404268 38984
rect 404320 38972 404326 39024
rect 405826 38972 405832 39024
rect 405884 39012 405890 39024
rect 407022 39012 407028 39024
rect 405884 38984 407028 39012
rect 405884 38972 405890 38984
rect 407022 38972 407028 38984
rect 407080 38972 407086 39024
rect 417050 38972 417056 39024
rect 417108 39012 417114 39024
rect 417970 39012 417976 39024
rect 417108 38984 417976 39012
rect 417108 38972 417114 38984
rect 417970 38972 417976 38984
rect 418028 38972 418034 39024
rect 418706 38972 418712 39024
rect 418764 39012 418770 39024
rect 419442 39012 419448 39024
rect 418764 38984 419448 39012
rect 418764 38972 418770 38984
rect 419442 38972 419448 38984
rect 419500 38972 419506 39024
rect 419626 38972 419632 39024
rect 419684 39012 419690 39024
rect 420822 39012 420828 39024
rect 419684 38984 420828 39012
rect 419684 38972 419690 38984
rect 420822 38972 420828 38984
rect 420880 38972 420886 39024
rect 423030 38972 423036 39024
rect 423088 39012 423094 39024
rect 423582 39012 423588 39024
rect 423088 38984 423588 39012
rect 423088 38972 423094 38984
rect 423582 38972 423588 38984
rect 423640 38972 423646 39024
rect 425606 38972 425612 39024
rect 425664 39012 425670 39024
rect 426342 39012 426348 39024
rect 425664 38984 426348 39012
rect 425664 38972 425670 38984
rect 426342 38972 426348 38984
rect 426400 38972 426406 39024
rect 428182 38972 428188 39024
rect 428240 39012 428246 39024
rect 429102 39012 429108 39024
rect 428240 38984 429108 39012
rect 428240 38972 428246 38984
rect 429102 38972 429108 38984
rect 429160 38972 429166 39024
rect 429930 38972 429936 39024
rect 429988 39012 429994 39024
rect 430482 39012 430488 39024
rect 429988 38984 430488 39012
rect 429988 38972 429994 38984
rect 430482 38972 430488 38984
rect 430540 38972 430546 39024
rect 430758 38972 430764 39024
rect 430816 39012 430822 39024
rect 431862 39012 431868 39024
rect 430816 38984 431868 39012
rect 430816 38972 430822 38984
rect 431862 38972 431868 38984
rect 431920 38972 431926 39024
rect 432506 38972 432512 39024
rect 432564 39012 432570 39024
rect 433242 39012 433248 39024
rect 432564 38984 433248 39012
rect 432564 38972 432570 38984
rect 433242 38972 433248 38984
rect 433300 38972 433306 39024
rect 433334 38972 433340 39024
rect 433392 39012 433398 39024
rect 434622 39012 434628 39024
rect 433392 38984 434628 39012
rect 433392 38972 433398 38984
rect 434622 38972 434628 38984
rect 434680 38972 434686 39024
rect 435082 38972 435088 39024
rect 435140 39012 435146 39024
rect 436002 39012 436008 39024
rect 435140 38984 436008 39012
rect 435140 38972 435146 38984
rect 436002 38972 436008 38984
rect 436060 38972 436066 39024
rect 436830 38972 436836 39024
rect 436888 39012 436894 39024
rect 437382 39012 437388 39024
rect 436888 38984 437388 39012
rect 436888 38972 436894 38984
rect 437382 38972 437388 38984
rect 437440 38972 437446 39024
rect 437658 38972 437664 39024
rect 437716 39012 437722 39024
rect 438762 39012 438768 39024
rect 437716 38984 438768 39012
rect 437716 38972 437722 38984
rect 438762 38972 438768 38984
rect 438820 38972 438826 39024
rect 440234 38972 440240 39024
rect 440292 39012 440298 39024
rect 441522 39012 441528 39024
rect 440292 38984 441528 39012
rect 440292 38972 440298 38984
rect 441522 38972 441528 38984
rect 441580 38972 441586 39024
rect 443730 38972 443736 39024
rect 443788 39012 443794 39024
rect 444282 39012 444288 39024
rect 443788 38984 444288 39012
rect 443788 38972 443794 38984
rect 444282 38972 444288 38984
rect 444340 38972 444346 39024
rect 446306 38972 446312 39024
rect 446364 39012 446370 39024
rect 447042 39012 447048 39024
rect 446364 38984 447048 39012
rect 446364 38972 446370 38984
rect 447042 38972 447048 38984
rect 447100 38972 447106 39024
rect 448882 38972 448888 39024
rect 448940 39012 448946 39024
rect 449802 39012 449808 39024
rect 448940 38984 449808 39012
rect 448940 38972 448946 38984
rect 449802 38972 449808 38984
rect 449860 38972 449866 39024
rect 450630 38972 450636 39024
rect 450688 39012 450694 39024
rect 451182 39012 451188 39024
rect 450688 38984 451188 39012
rect 450688 38972 450694 38984
rect 451182 38972 451188 38984
rect 451240 38972 451246 39024
rect 451458 38972 451464 39024
rect 451516 39012 451522 39024
rect 452470 39012 452476 39024
rect 451516 38984 452476 39012
rect 451516 38972 451522 38984
rect 452470 38972 452476 38984
rect 452528 38972 452534 39024
rect 453206 38972 453212 39024
rect 453264 39012 453270 39024
rect 453942 39012 453948 39024
rect 453264 38984 453948 39012
rect 453264 38972 453270 38984
rect 453942 38972 453948 38984
rect 454000 38972 454006 39024
rect 454034 38972 454040 39024
rect 454092 39012 454098 39024
rect 455322 39012 455328 39024
rect 454092 38984 455328 39012
rect 454092 38972 454098 38984
rect 455322 38972 455328 38984
rect 455380 38972 455386 39024
rect 455782 38972 455788 39024
rect 455840 39012 455846 39024
rect 456702 39012 456708 39024
rect 455840 38984 456708 39012
rect 455840 38972 455846 38984
rect 456702 38972 456708 38984
rect 456760 38972 456766 39024
rect 457530 38972 457536 39024
rect 457588 39012 457594 39024
rect 458082 39012 458088 39024
rect 457588 38984 458088 39012
rect 457588 38972 457594 38984
rect 458082 38972 458088 38984
rect 458140 38972 458146 39024
rect 458358 38972 458364 39024
rect 458416 39012 458422 39024
rect 459462 39012 459468 39024
rect 458416 38984 459468 39012
rect 458416 38972 458422 38984
rect 459462 38972 459468 38984
rect 459520 38972 459526 39024
rect 460934 38972 460940 39024
rect 460992 39012 460998 39024
rect 462222 39012 462228 39024
rect 460992 38984 462228 39012
rect 460992 38972 460998 38984
rect 462222 38972 462228 38984
rect 462280 38972 462286 39024
rect 465258 38972 465264 39024
rect 465316 39012 465322 39024
rect 466270 39012 466276 39024
rect 465316 38984 466276 39012
rect 465316 38972 465322 38984
rect 466270 38972 466276 38984
rect 466328 38972 466334 39024
rect 42702 38904 42708 38956
rect 42760 38944 42766 38956
rect 72418 38944 72424 38956
rect 42760 38916 72424 38944
rect 42760 38904 42766 38916
rect 72418 38904 72424 38916
rect 72476 38904 72482 38956
rect 77202 38904 77208 38956
rect 77260 38944 77266 38956
rect 97442 38944 97448 38956
rect 77260 38916 97448 38944
rect 77260 38904 77266 38916
rect 97442 38904 97448 38916
rect 97500 38904 97506 38956
rect 137278 38904 137284 38956
rect 137336 38944 137342 38956
rect 140498 38944 140504 38956
rect 137336 38916 140504 38944
rect 137336 38904 137342 38916
rect 140498 38904 140504 38916
rect 140556 38904 140562 38956
rect 144822 38904 144828 38956
rect 144880 38944 144886 38956
rect 146478 38944 146484 38956
rect 144880 38916 146484 38944
rect 144880 38904 144886 38916
rect 146478 38904 146484 38916
rect 146536 38904 146542 38956
rect 147582 38904 147588 38956
rect 147640 38944 147646 38956
rect 149054 38944 149060 38956
rect 147640 38916 149060 38944
rect 147640 38904 147646 38916
rect 149054 38904 149060 38916
rect 149112 38904 149118 38956
rect 154574 38904 154580 38956
rect 154632 38944 154638 38956
rect 155126 38944 155132 38956
rect 154632 38916 155132 38944
rect 154632 38904 154638 38916
rect 155126 38904 155132 38916
rect 155184 38904 155190 38956
rect 160370 38904 160376 38956
rect 160428 38944 160434 38956
rect 161382 38944 161388 38956
rect 160428 38916 161388 38944
rect 160428 38904 160434 38916
rect 161382 38904 161388 38916
rect 161440 38904 161446 38956
rect 176746 38904 176752 38956
rect 176804 38944 176810 38956
rect 177850 38944 177856 38956
rect 176804 38916 177856 38944
rect 176804 38904 176810 38916
rect 177850 38904 177856 38916
rect 177908 38904 177914 38956
rect 222378 38904 222384 38956
rect 222436 38944 222442 38956
rect 223482 38944 223488 38956
rect 222436 38916 223488 38944
rect 222436 38904 222442 38916
rect 223482 38904 223488 38916
rect 223540 38904 223546 38956
rect 231854 38904 231860 38956
rect 231912 38944 231918 38956
rect 233050 38944 233056 38956
rect 231912 38916 233056 38944
rect 231912 38904 231918 38916
rect 233050 38904 233056 38916
rect 233108 38904 233114 38956
rect 284386 38904 284392 38956
rect 284444 38944 284450 38956
rect 285490 38944 285496 38956
rect 284444 38916 285496 38944
rect 284444 38904 284450 38916
rect 285490 38904 285496 38916
rect 285548 38904 285554 38956
rect 308490 38904 308496 38956
rect 308548 38944 308554 38956
rect 309042 38944 309048 38956
rect 308548 38916 309048 38944
rect 308548 38904 308554 38916
rect 309042 38904 309048 38916
rect 309100 38904 309106 38956
rect 322290 38904 322296 38956
rect 322348 38944 322354 38956
rect 322842 38944 322848 38956
rect 322348 38916 322848 38944
rect 322348 38904 322354 38916
rect 322842 38904 322848 38916
rect 322900 38904 322906 38956
rect 367094 38904 367100 38956
rect 367152 38944 367158 38956
rect 368290 38944 368296 38956
rect 367152 38916 368296 38944
rect 367152 38904 367158 38916
rect 368290 38904 368296 38916
rect 368348 38904 368354 38956
rect 371326 38904 371332 38956
rect 371384 38944 371390 38956
rect 372522 38944 372528 38956
rect 371384 38916 372528 38944
rect 371384 38904 371390 38916
rect 372522 38904 372528 38916
rect 372580 38904 372586 38956
rect 378226 38904 378232 38956
rect 378284 38944 378290 38956
rect 379422 38944 379428 38956
rect 378284 38916 379428 38944
rect 378284 38904 378290 38916
rect 379422 38904 379428 38916
rect 379480 38904 379486 38956
rect 426526 38904 426532 38956
rect 426584 38944 426590 38956
rect 429838 38944 429844 38956
rect 426584 38916 429844 38944
rect 426584 38904 426590 38916
rect 429838 38904 429844 38916
rect 429896 38904 429902 38956
rect 464338 38904 464344 38956
rect 464396 38944 464402 38956
rect 464982 38944 464988 38956
rect 464396 38916 464988 38944
rect 464396 38904 464402 38916
rect 464982 38904 464988 38916
rect 465040 38904 465046 38956
rect 43438 38836 43444 38888
rect 43496 38876 43502 38888
rect 49142 38876 49148 38888
rect 43496 38848 49148 38876
rect 43496 38836 43502 38848
rect 49142 38836 49148 38848
rect 49200 38836 49206 38888
rect 50982 38836 50988 38888
rect 51040 38876 51046 38888
rect 78398 38876 78404 38888
rect 51040 38848 78404 38876
rect 51040 38836 51046 38848
rect 78398 38836 78404 38848
rect 78456 38836 78462 38888
rect 79962 38836 79968 38888
rect 80020 38876 80026 38888
rect 100018 38876 100024 38888
rect 80020 38848 100024 38876
rect 80020 38836 80026 38848
rect 100018 38836 100024 38848
rect 100076 38836 100082 38888
rect 133782 38836 133788 38888
rect 133840 38876 133846 38888
rect 138750 38876 138756 38888
rect 133840 38848 138756 38876
rect 133840 38836 133846 38848
rect 138750 38836 138756 38848
rect 138808 38836 138814 38888
rect 304166 38836 304172 38888
rect 304224 38876 304230 38888
rect 304902 38876 304908 38888
rect 304224 38848 304908 38876
rect 304224 38836 304230 38848
rect 304902 38836 304908 38848
rect 304960 38836 304966 38888
rect 381722 38836 381728 38888
rect 381780 38876 381786 38888
rect 382182 38876 382188 38888
rect 381780 38848 382188 38876
rect 381780 38836 381786 38848
rect 382182 38836 382188 38848
rect 382240 38836 382246 38888
rect 48958 38768 48964 38820
rect 49016 38808 49022 38820
rect 62942 38808 62948 38820
rect 49016 38780 62948 38808
rect 49016 38768 49022 38780
rect 62942 38768 62948 38780
rect 63000 38768 63006 38820
rect 64138 38768 64144 38820
rect 64196 38808 64202 38820
rect 75914 38808 75920 38820
rect 64196 38780 75920 38808
rect 64196 38768 64202 38780
rect 75914 38768 75920 38780
rect 75972 38768 75978 38820
rect 78582 38768 78588 38820
rect 78640 38808 78646 38820
rect 99098 38808 99104 38820
rect 78640 38780 99104 38808
rect 78640 38768 78646 38780
rect 99098 38768 99104 38780
rect 99156 38768 99162 38820
rect 135162 38768 135168 38820
rect 135220 38808 135226 38820
rect 139578 38808 139584 38820
rect 135220 38780 139584 38808
rect 135220 38768 135226 38780
rect 139578 38768 139584 38780
rect 139636 38768 139642 38820
rect 164694 38768 164700 38820
rect 164752 38808 164758 38820
rect 165522 38808 165528 38820
rect 164752 38780 165528 38808
rect 164752 38768 164758 38780
rect 165522 38768 165528 38780
rect 165580 38768 165586 38820
rect 168098 38768 168104 38820
rect 168156 38808 168162 38820
rect 169018 38808 169024 38820
rect 168156 38780 169024 38808
rect 168156 38768 168162 38780
rect 169018 38768 169024 38780
rect 169076 38768 169082 38820
rect 174170 38768 174176 38820
rect 174228 38808 174234 38820
rect 175090 38808 175096 38820
rect 174228 38780 175096 38808
rect 174228 38768 174234 38780
rect 175090 38768 175096 38780
rect 175148 38768 175154 38820
rect 204254 38768 204260 38820
rect 204312 38808 204318 38820
rect 205450 38808 205456 38820
rect 204312 38780 205456 38808
rect 204312 38768 204318 38780
rect 205450 38768 205456 38780
rect 205508 38768 205514 38820
rect 221550 38768 221556 38820
rect 221608 38808 221614 38820
rect 228358 38808 228364 38820
rect 221608 38780 228364 38808
rect 221608 38768 221614 38780
rect 228358 38768 228364 38780
rect 228416 38768 228422 38820
rect 233602 38768 233608 38820
rect 233660 38808 233666 38820
rect 234522 38808 234528 38820
rect 233660 38780 234528 38808
rect 233660 38768 233666 38780
rect 234522 38768 234528 38780
rect 234580 38768 234586 38820
rect 287790 38768 287796 38820
rect 287848 38808 287854 38820
rect 288342 38808 288348 38820
rect 287848 38780 288348 38808
rect 287848 38768 287854 38780
rect 288342 38768 288348 38780
rect 288400 38768 288406 38820
rect 386874 38768 386880 38820
rect 386932 38808 386938 38820
rect 387702 38808 387708 38820
rect 386932 38780 387708 38808
rect 386932 38768 386938 38780
rect 387702 38768 387708 38780
rect 387760 38768 387766 38820
rect 55858 38700 55864 38752
rect 55916 38740 55922 38752
rect 68094 38740 68100 38752
rect 55916 38712 68100 38740
rect 55916 38700 55922 38712
rect 68094 38700 68100 38712
rect 68152 38700 68158 38752
rect 82722 38700 82728 38752
rect 82780 38740 82786 38752
rect 101674 38740 101680 38752
rect 82780 38712 101680 38740
rect 82780 38700 82786 38712
rect 101674 38700 101680 38712
rect 101732 38700 101738 38752
rect 144730 38700 144736 38752
rect 144788 38740 144794 38752
rect 147398 38740 147404 38752
rect 144788 38712 147404 38740
rect 144788 38700 144794 38712
rect 147398 38700 147404 38712
rect 147456 38700 147462 38752
rect 439406 38700 439412 38752
rect 439464 38740 439470 38752
rect 440142 38740 440148 38752
rect 439464 38712 440148 38740
rect 439464 38700 439470 38712
rect 440142 38700 440148 38712
rect 440200 38700 440206 38752
rect 46198 38632 46204 38684
rect 46256 38672 46262 38684
rect 56042 38672 56048 38684
rect 46256 38644 56048 38672
rect 46256 38632 46262 38644
rect 56042 38632 56048 38644
rect 56100 38632 56106 38684
rect 62758 38632 62764 38684
rect 62816 38672 62822 38684
rect 73246 38672 73252 38684
rect 62816 38644 73252 38672
rect 62816 38632 62822 38644
rect 73246 38632 73252 38644
rect 73304 38632 73310 38684
rect 93762 38632 93768 38684
rect 93820 38672 93826 38684
rect 109494 38672 109500 38684
rect 93820 38644 109500 38672
rect 93820 38632 93826 38644
rect 109494 38632 109500 38644
rect 109552 38632 109558 38684
rect 124122 38632 124128 38684
rect 124180 38672 124186 38684
rect 131850 38672 131856 38684
rect 124180 38644 131856 38672
rect 124180 38632 124186 38644
rect 131850 38632 131856 38644
rect 131908 38632 131914 38684
rect 385126 38360 385132 38412
rect 385184 38400 385190 38412
rect 470594 38400 470600 38412
rect 385184 38372 470600 38400
rect 385184 38360 385190 38372
rect 470594 38360 470600 38372
rect 470652 38360 470658 38412
rect 407574 38292 407580 38344
rect 407632 38332 407638 38344
rect 500954 38332 500960 38344
rect 407632 38304 500960 38332
rect 407632 38292 407638 38304
rect 500954 38292 500960 38304
rect 501012 38292 501018 38344
rect 412726 38224 412732 38276
rect 412784 38264 412790 38276
rect 507854 38264 507860 38276
rect 412784 38236 507860 38264
rect 412784 38224 412790 38236
rect 507854 38224 507860 38236
rect 507912 38224 507918 38276
rect 421282 38156 421288 38208
rect 421340 38196 421346 38208
rect 520274 38196 520280 38208
rect 421340 38168 520280 38196
rect 421340 38156 421346 38168
rect 520274 38156 520280 38168
rect 520332 38156 520338 38208
rect 437290 38088 437296 38140
rect 437348 38128 437354 38140
rect 538214 38128 538220 38140
rect 437348 38100 538220 38128
rect 437348 38088 437354 38100
rect 538214 38088 538220 38100
rect 538272 38088 538278 38140
rect 444190 38020 444196 38072
rect 444248 38060 444254 38072
rect 547874 38060 547880 38072
rect 444248 38032 547880 38060
rect 444248 38020 444254 38032
rect 547874 38020 547880 38032
rect 547932 38020 547938 38072
rect 444558 37952 444564 38004
rect 444616 37992 444622 38004
rect 551278 37992 551284 38004
rect 444616 37964 551284 37992
rect 444616 37952 444622 37964
rect 551278 37952 551284 37964
rect 551336 37952 551342 38004
rect 299198 37884 299204 37936
rect 299256 37924 299262 37936
rect 349154 37924 349160 37936
rect 299256 37896 349160 37924
rect 299256 37884 299262 37896
rect 349154 37884 349160 37896
rect 349212 37884 349218 37936
rect 349706 37884 349712 37936
rect 349764 37924 349770 37936
rect 398834 37924 398840 37936
rect 349764 37896 398840 37924
rect 349764 37884 349770 37896
rect 398834 37884 398840 37896
rect 398892 37884 398898 37936
rect 452286 37884 452292 37936
rect 452344 37924 452350 37936
rect 560938 37924 560944 37936
rect 452344 37896 560944 37924
rect 452344 37884 452350 37896
rect 560938 37884 560944 37896
rect 560996 37884 561002 37936
rect 406654 36864 406660 36916
rect 406712 36904 406718 36916
rect 499574 36904 499580 36916
rect 406712 36876 499580 36904
rect 406712 36864 406718 36876
rect 499574 36864 499580 36876
rect 499632 36864 499638 36916
rect 411806 36796 411812 36848
rect 411864 36836 411870 36848
rect 506474 36836 506480 36848
rect 411864 36808 506480 36836
rect 411864 36796 411870 36808
rect 506474 36796 506480 36808
rect 506532 36796 506538 36848
rect 447134 36728 447140 36780
rect 447192 36768 447198 36780
rect 556246 36768 556252 36780
rect 447192 36740 556252 36768
rect 447192 36728 447198 36740
rect 556246 36728 556252 36740
rect 556304 36728 556310 36780
rect 449710 36660 449716 36712
rect 449768 36700 449774 36712
rect 558178 36700 558184 36712
rect 449768 36672 558184 36700
rect 449768 36660 449774 36672
rect 558178 36660 558184 36672
rect 558236 36660 558242 36712
rect 454862 36592 454868 36644
rect 454920 36632 454926 36644
rect 565814 36632 565820 36644
rect 454920 36604 565820 36632
rect 454920 36592 454926 36604
rect 565814 36592 565820 36604
rect 565872 36592 565878 36644
rect 460106 36524 460112 36576
rect 460164 36564 460170 36576
rect 572714 36564 572720 36576
rect 460164 36536 572720 36564
rect 460164 36524 460170 36536
rect 572714 36524 572720 36536
rect 572772 36524 572778 36576
rect 397362 35232 397368 35284
rect 397420 35272 397426 35284
rect 485774 35272 485780 35284
rect 397420 35244 485780 35272
rect 397420 35232 397426 35244
rect 485774 35232 485780 35244
rect 485832 35232 485838 35284
rect 417970 35164 417976 35216
rect 418028 35204 418034 35216
rect 514754 35204 514760 35216
rect 418028 35176 514760 35204
rect 418028 35164 418034 35176
rect 514754 35164 514760 35176
rect 514812 35164 514818 35216
rect 378042 33736 378048 33788
rect 378100 33776 378106 33788
rect 459554 33776 459560 33788
rect 378100 33748 459560 33776
rect 378100 33736 378106 33748
rect 459554 33736 459560 33748
rect 459612 33736 459618 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 11698 33096 11704 33108
rect 2924 33068 11704 33096
rect 2924 33056 2930 33068
rect 11698 33056 11704 33068
rect 11756 33056 11762 33108
rect 383470 31016 383476 31068
rect 383528 31056 383534 31068
rect 466454 31056 466460 31068
rect 383528 31028 466460 31056
rect 383528 31016 383534 31028
rect 466454 31016 466460 31028
rect 466512 31016 466518 31068
rect 339402 29588 339408 29640
rect 339460 29628 339466 29640
rect 407206 29628 407212 29640
rect 339460 29600 407212 29628
rect 339460 29588 339466 29600
rect 407206 29588 407212 29600
rect 407264 29588 407270 29640
rect 375190 28228 375196 28280
rect 375248 28268 375254 28280
rect 456886 28268 456892 28280
rect 375248 28240 456892 28268
rect 375248 28228 375254 28240
rect 456886 28228 456892 28240
rect 456944 28228 456950 28280
rect 372430 26868 372436 26920
rect 372488 26908 372494 26920
rect 452654 26908 452660 26920
rect 372488 26880 452660 26908
rect 372488 26868 372494 26880
rect 452654 26868 452660 26880
rect 452712 26868 452718 26920
rect 357342 25508 357348 25560
rect 357400 25548 357406 25560
rect 432046 25548 432052 25560
rect 357400 25520 432052 25548
rect 357400 25508 357406 25520
rect 432046 25508 432052 25520
rect 432104 25508 432110 25560
rect 342070 24080 342076 24132
rect 342128 24120 342134 24132
rect 409874 24120 409880 24132
rect 342128 24092 409880 24120
rect 342128 24080 342134 24092
rect 409874 24080 409880 24092
rect 409932 24080 409938 24132
rect 328362 22720 328368 22772
rect 328420 22760 328426 22772
rect 391934 22760 391940 22772
rect 328420 22732 391940 22760
rect 328420 22720 328426 22732
rect 391934 22720 391940 22732
rect 391992 22720 391998 22772
rect 401410 22720 401416 22772
rect 401468 22760 401474 22772
rect 492674 22760 492680 22772
rect 401468 22732 492680 22760
rect 401468 22720 401474 22732
rect 492674 22720 492680 22732
rect 492732 22720 492738 22772
rect 280798 21360 280804 21412
rect 280856 21400 280862 21412
rect 324314 21400 324320 21412
rect 280856 21372 324320 21400
rect 280856 21360 280862 21372
rect 324314 21360 324320 21372
rect 324372 21360 324378 21412
rect 325602 21360 325608 21412
rect 325660 21400 325666 21412
rect 387794 21400 387800 21412
rect 325660 21372 387800 21400
rect 325660 21360 325666 21372
rect 387794 21360 387800 21372
rect 387852 21360 387858 21412
rect 388438 21360 388444 21412
rect 388496 21400 388502 21412
rect 463694 21400 463700 21412
rect 388496 21372 463700 21400
rect 388496 21360 388502 21372
rect 463694 21360 463700 21372
rect 463752 21360 463758 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 40678 20652 40684 20664
rect 3476 20624 40684 20652
rect 3476 20612 3482 20624
rect 40678 20612 40684 20624
rect 40736 20612 40742 20664
rect 335998 18572 336004 18624
rect 336056 18612 336062 18624
rect 380894 18612 380900 18624
rect 336056 18584 380900 18612
rect 336056 18572 336062 18584
rect 380894 18572 380900 18584
rect 380952 18572 380958 18624
rect 381538 18572 381544 18624
rect 381596 18612 381602 18624
rect 448514 18612 448520 18624
rect 381596 18584 448520 18612
rect 381596 18572 381602 18584
rect 448514 18572 448520 18584
rect 448572 18572 448578 18624
rect 286870 17280 286876 17332
rect 286928 17320 286934 17332
rect 335354 17320 335360 17332
rect 286928 17292 335360 17320
rect 286928 17280 286934 17292
rect 335354 17280 335360 17292
rect 335412 17280 335418 17332
rect 317230 17212 317236 17264
rect 317288 17252 317294 17264
rect 376754 17252 376760 17264
rect 317288 17224 376760 17252
rect 317288 17212 317294 17224
rect 376754 17212 376760 17224
rect 376812 17212 376818 17264
rect 377398 17212 377404 17264
rect 377456 17252 377462 17264
rect 438854 17252 438860 17264
rect 377456 17224 438860 17252
rect 377456 17212 377462 17224
rect 438854 17212 438860 17224
rect 438912 17212 438918 17264
rect 289722 15920 289728 15972
rect 289780 15960 289786 15972
rect 338666 15960 338672 15972
rect 289780 15932 338672 15960
rect 289780 15920 289786 15932
rect 338666 15920 338672 15932
rect 338724 15920 338730 15972
rect 336642 15852 336648 15904
rect 336700 15892 336706 15904
rect 403618 15892 403624 15904
rect 336700 15864 403624 15892
rect 336700 15852 336706 15864
rect 403618 15852 403624 15864
rect 403676 15852 403682 15904
rect 307662 14424 307668 14476
rect 307720 14464 307726 14476
rect 363506 14464 363512 14476
rect 307720 14436 363512 14464
rect 307720 14424 307726 14436
rect 363506 14424 363512 14436
rect 363564 14424 363570 14476
rect 363598 14424 363604 14476
rect 363656 14464 363662 14476
rect 420914 14464 420920 14476
rect 363656 14436 420920 14464
rect 363656 14424 363662 14436
rect 420914 14424 420920 14436
rect 420972 14424 420978 14476
rect 299290 13064 299296 13116
rect 299348 13104 299354 13116
rect 299348 13076 335354 13104
rect 299348 13064 299354 13076
rect 335326 13036 335354 13076
rect 352558 13064 352564 13116
rect 352616 13104 352622 13116
rect 414290 13104 414296 13116
rect 352616 13076 414296 13104
rect 352616 13064 352622 13076
rect 414290 13064 414296 13076
rect 414348 13064 414354 13116
rect 352834 13036 352840 13048
rect 335326 13008 352840 13036
rect 352834 12996 352840 13008
rect 352892 12996 352898 13048
rect 304902 11704 304908 11756
rect 304960 11744 304966 11756
rect 359274 11744 359280 11756
rect 304960 11716 359280 11744
rect 304960 11704 304966 11716
rect 359274 11704 359280 11716
rect 359332 11704 359338 11756
rect 368290 11704 368296 11756
rect 368348 11744 368354 11756
rect 445754 11744 445760 11756
rect 368348 11716 445760 11744
rect 368348 11704 368354 11716
rect 445754 11704 445760 11716
rect 445812 11704 445818 11756
rect 233050 10276 233056 10328
rect 233108 10316 233114 10328
rect 260650 10316 260656 10328
rect 233108 10288 260656 10316
rect 233108 10276 233114 10288
rect 260650 10276 260656 10288
rect 260708 10276 260714 10328
rect 278590 10276 278596 10328
rect 278648 10316 278654 10328
rect 324406 10316 324412 10328
rect 278648 10288 324412 10316
rect 278648 10276 278654 10288
rect 324406 10276 324412 10288
rect 324464 10276 324470 10328
rect 324958 10276 324964 10328
rect 325016 10316 325022 10328
rect 370130 10316 370136 10328
rect 325016 10288 370136 10316
rect 325016 10276 325022 10288
rect 370130 10276 370136 10288
rect 370188 10276 370194 10328
rect 458082 10276 458088 10328
rect 458140 10316 458146 10328
rect 569218 10316 569224 10328
rect 458140 10288 569224 10316
rect 458140 10276 458146 10288
rect 569218 10276 569224 10288
rect 569276 10276 569282 10328
rect 264790 8984 264796 9036
rect 264848 9024 264854 9036
rect 304350 9024 304356 9036
rect 264848 8996 304356 9024
rect 264848 8984 264854 8996
rect 304350 8984 304356 8996
rect 304408 8984 304414 9036
rect 390370 8984 390376 9036
rect 390428 9024 390434 9036
rect 478138 9024 478144 9036
rect 390428 8996 478144 9024
rect 390428 8984 390434 8996
rect 478138 8984 478144 8996
rect 478196 8984 478202 9036
rect 296530 8916 296536 8968
rect 296588 8956 296594 8968
rect 349246 8956 349252 8968
rect 296588 8928 349252 8956
rect 296588 8916 296594 8928
rect 349246 8916 349252 8928
rect 349304 8916 349310 8968
rect 359550 8916 359556 8968
rect 359608 8956 359614 8968
rect 389450 8956 389456 8968
rect 359608 8928 389456 8956
rect 359608 8916 359614 8928
rect 389450 8916 389456 8928
rect 389508 8916 389514 8968
rect 411162 8916 411168 8968
rect 411220 8956 411226 8968
rect 506474 8956 506480 8968
rect 411220 8928 506480 8956
rect 411220 8916 411226 8928
rect 506474 8916 506480 8928
rect 506532 8916 506538 8968
rect 338758 8236 338764 8288
rect 338816 8276 338822 8288
rect 339862 8276 339868 8288
rect 338816 8248 339868 8276
rect 338816 8236 338822 8248
rect 339862 8236 339868 8248
rect 339920 8236 339926 8288
rect 411898 8236 411904 8288
rect 411956 8276 411962 8288
rect 435542 8276 435548 8288
rect 411956 8248 435548 8276
rect 411956 8236 411962 8248
rect 435542 8236 435548 8248
rect 435600 8236 435606 8288
rect 441338 8236 441344 8288
rect 441396 8276 441402 8288
rect 441522 8276 441528 8288
rect 441396 8248 441528 8276
rect 441396 8236 441402 8248
rect 441522 8236 441528 8248
rect 441580 8236 441586 8288
rect 413278 8168 413284 8220
rect 413336 8208 413342 8220
rect 442626 8208 442632 8220
rect 413336 8180 442632 8208
rect 413336 8168 413342 8180
rect 442626 8168 442632 8180
rect 442684 8168 442690 8220
rect 394602 8100 394608 8152
rect 394660 8140 394666 8152
rect 484026 8140 484032 8152
rect 394660 8112 484032 8140
rect 394660 8100 394666 8112
rect 484026 8100 484032 8112
rect 484084 8100 484090 8152
rect 400122 8032 400128 8084
rect 400180 8072 400186 8084
rect 491110 8072 491116 8084
rect 400180 8044 491116 8072
rect 400180 8032 400186 8044
rect 491110 8032 491116 8044
rect 491168 8032 491174 8084
rect 413830 7964 413836 8016
rect 413888 8004 413894 8016
rect 510062 8004 510068 8016
rect 413888 7976 510068 8004
rect 413888 7964 413894 7976
rect 510062 7964 510068 7976
rect 510120 7964 510126 8016
rect 322198 7896 322204 7948
rect 322256 7936 322262 7948
rect 356330 7936 356336 7948
rect 322256 7908 356336 7936
rect 322256 7896 322262 7908
rect 356330 7896 356336 7908
rect 356388 7896 356394 7948
rect 419442 7896 419448 7948
rect 419500 7936 419506 7948
rect 517146 7936 517152 7948
rect 419500 7908 517152 7936
rect 419500 7896 419506 7908
rect 517146 7896 517152 7908
rect 517204 7896 517210 7948
rect 310330 7828 310336 7880
rect 310388 7868 310394 7880
rect 368198 7868 368204 7880
rect 310388 7840 368204 7868
rect 310388 7828 310394 7840
rect 368198 7828 368204 7840
rect 368256 7828 368262 7880
rect 429838 7828 429844 7880
rect 429896 7868 429902 7880
rect 527818 7868 527824 7880
rect 429896 7840 527824 7868
rect 429896 7828 429902 7840
rect 527818 7828 527824 7840
rect 527876 7828 527882 7880
rect 318702 7760 318708 7812
rect 318760 7800 318766 7812
rect 378870 7800 378876 7812
rect 318760 7772 378876 7800
rect 318760 7760 318766 7772
rect 378870 7760 378876 7772
rect 378928 7760 378934 7812
rect 431770 7760 431776 7812
rect 431828 7800 431834 7812
rect 534902 7800 534908 7812
rect 431828 7772 534908 7800
rect 431828 7760 431834 7772
rect 534902 7760 534908 7772
rect 534960 7760 534966 7812
rect 321370 7692 321376 7744
rect 321428 7732 321434 7744
rect 382366 7732 382372 7744
rect 321428 7704 382372 7732
rect 321428 7692 321434 7704
rect 382366 7692 382372 7704
rect 382424 7692 382430 7744
rect 395338 7692 395344 7744
rect 395396 7732 395402 7744
rect 417878 7732 417884 7744
rect 395396 7704 417884 7732
rect 395396 7692 395402 7704
rect 417878 7692 417884 7704
rect 417936 7692 417942 7744
rect 429010 7692 429016 7744
rect 429068 7732 429074 7744
rect 531314 7732 531320 7744
rect 429068 7704 531320 7732
rect 429068 7692 429074 7704
rect 531314 7692 531320 7704
rect 531372 7692 531378 7744
rect 249058 7624 249064 7676
rect 249116 7664 249122 7676
rect 281902 7664 281908 7676
rect 249116 7636 281908 7664
rect 249116 7624 249122 7636
rect 281902 7624 281908 7636
rect 281960 7624 281966 7676
rect 282178 7624 282184 7676
rect 282236 7664 282242 7676
rect 317230 7664 317236 7676
rect 282236 7636 317236 7664
rect 282236 7624 282242 7636
rect 317230 7624 317236 7636
rect 317288 7624 317294 7676
rect 324130 7624 324136 7676
rect 324188 7664 324194 7676
rect 385954 7664 385960 7676
rect 324188 7636 385960 7664
rect 324188 7624 324194 7636
rect 385954 7624 385960 7636
rect 386012 7624 386018 7676
rect 396718 7624 396724 7676
rect 396776 7664 396782 7676
rect 424870 7664 424876 7676
rect 396776 7636 424876 7664
rect 396776 7624 396782 7636
rect 424870 7624 424876 7636
rect 424928 7624 424934 7676
rect 437382 7624 437388 7676
rect 437440 7664 437446 7676
rect 541986 7664 541992 7676
rect 437440 7636 541992 7664
rect 437440 7624 437446 7636
rect 541986 7624 541992 7636
rect 542044 7624 542050 7676
rect 228358 7556 228364 7608
rect 228416 7596 228422 7608
rect 246390 7596 246396 7608
rect 228416 7568 246396 7596
rect 228416 7556 228422 7568
rect 246390 7556 246396 7568
rect 246448 7556 246454 7608
rect 277302 7556 277308 7608
rect 277360 7596 277366 7608
rect 322106 7596 322112 7608
rect 277360 7568 322112 7596
rect 277360 7556 277366 7568
rect 322106 7556 322112 7568
rect 322164 7556 322170 7608
rect 354490 7556 354496 7608
rect 354548 7596 354554 7608
rect 428458 7596 428464 7608
rect 354548 7568 428464 7596
rect 354548 7556 354554 7568
rect 428458 7556 428464 7568
rect 428516 7556 428522 7608
rect 440142 7556 440148 7608
rect 440200 7596 440206 7608
rect 545482 7596 545488 7608
rect 440200 7568 545488 7596
rect 440200 7556 440206 7568
rect 545482 7556 545488 7568
rect 545540 7556 545546 7608
rect 370498 6876 370504 6928
rect 370556 6916 370562 6928
rect 375282 6916 375288 6928
rect 370556 6888 375288 6916
rect 370556 6876 370562 6888
rect 375282 6876 375288 6888
rect 375340 6876 375346 6928
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 29638 6848 29644 6860
rect 3476 6820 29644 6848
rect 3476 6808 3482 6820
rect 29638 6808 29644 6820
rect 29696 6808 29702 6860
rect 379330 6808 379336 6860
rect 379388 6848 379394 6860
rect 462774 6848 462780 6860
rect 379388 6820 462780 6848
rect 379388 6808 379394 6820
rect 462774 6808 462780 6820
rect 462832 6808 462838 6860
rect 467190 6808 467196 6860
rect 467248 6848 467254 6860
rect 505370 6848 505376 6860
rect 467248 6820 505376 6848
rect 467248 6808 467254 6820
rect 505370 6808 505376 6820
rect 505428 6808 505434 6860
rect 384942 6740 384948 6792
rect 385000 6780 385006 6792
rect 469858 6780 469864 6792
rect 385000 6752 469864 6780
rect 385000 6740 385006 6752
rect 469858 6740 469864 6752
rect 469916 6740 469922 6792
rect 390462 6672 390468 6724
rect 390520 6712 390526 6724
rect 476942 6712 476948 6724
rect 390520 6684 476948 6712
rect 390520 6672 390526 6684
rect 476942 6672 476948 6684
rect 477000 6672 477006 6724
rect 292390 6604 292396 6656
rect 292448 6644 292454 6656
rect 343358 6644 343364 6656
rect 292448 6616 343364 6644
rect 292448 6604 292454 6616
rect 343358 6604 343364 6616
rect 343416 6604 343422 6656
rect 356698 6604 356704 6656
rect 356756 6644 356762 6656
rect 364610 6644 364616 6656
rect 356756 6616 364616 6644
rect 356756 6604 356762 6616
rect 364610 6604 364616 6616
rect 364668 6604 364674 6656
rect 387702 6604 387708 6656
rect 387760 6644 387766 6656
rect 473446 6644 473452 6656
rect 387760 6616 473452 6644
rect 387760 6604 387766 6616
rect 473446 6604 473452 6616
rect 473504 6604 473510 6656
rect 300670 6536 300676 6588
rect 300728 6576 300734 6588
rect 354030 6576 354036 6588
rect 300728 6548 354036 6576
rect 300728 6536 300734 6548
rect 354030 6536 354036 6548
rect 354088 6536 354094 6588
rect 359366 6536 359372 6588
rect 359424 6576 359430 6588
rect 390646 6576 390652 6588
rect 359424 6548 390652 6576
rect 359424 6536 359430 6548
rect 390646 6536 390652 6548
rect 390704 6536 390710 6588
rect 395982 6536 395988 6588
rect 396040 6576 396046 6588
rect 485222 6576 485228 6588
rect 396040 6548 485228 6576
rect 396040 6536 396046 6548
rect 485222 6536 485228 6548
rect 485280 6536 485286 6588
rect 306190 6468 306196 6520
rect 306248 6508 306254 6520
rect 361114 6508 361120 6520
rect 306248 6480 361120 6508
rect 306248 6468 306254 6480
rect 361114 6468 361120 6480
rect 361172 6468 361178 6520
rect 393222 6468 393228 6520
rect 393280 6508 393286 6520
rect 481726 6508 481732 6520
rect 393280 6480 481732 6508
rect 393280 6468 393286 6480
rect 481726 6468 481732 6480
rect 481784 6468 481790 6520
rect 310422 6400 310428 6452
rect 310480 6440 310486 6452
rect 366910 6440 366916 6452
rect 310480 6412 366916 6440
rect 310480 6400 310486 6412
rect 366910 6400 366916 6412
rect 366968 6400 366974 6452
rect 401502 6400 401508 6452
rect 401560 6440 401566 6452
rect 492306 6440 492312 6452
rect 401560 6412 492312 6440
rect 401560 6400 401566 6412
rect 492306 6400 492312 6412
rect 492364 6400 492370 6452
rect 313182 6332 313188 6384
rect 313240 6372 313246 6384
rect 371694 6372 371700 6384
rect 313240 6344 371700 6372
rect 313240 6332 313246 6344
rect 371694 6332 371700 6344
rect 371752 6332 371758 6384
rect 398742 6332 398748 6384
rect 398800 6372 398806 6384
rect 488810 6372 488816 6384
rect 398800 6344 488816 6372
rect 398800 6332 398806 6344
rect 488810 6332 488816 6344
rect 488868 6332 488874 6384
rect 489178 6332 489184 6384
rect 489236 6372 489242 6384
rect 498194 6372 498200 6384
rect 489236 6344 498200 6372
rect 489236 6332 489242 6344
rect 498194 6332 498200 6344
rect 498252 6332 498258 6384
rect 262950 6264 262956 6316
rect 263008 6304 263014 6316
rect 300670 6304 300676 6316
rect 263008 6276 300676 6304
rect 263008 6264 263014 6276
rect 300670 6264 300676 6276
rect 300728 6264 300734 6316
rect 314470 6264 314476 6316
rect 314528 6304 314534 6316
rect 374086 6304 374092 6316
rect 314528 6276 374092 6304
rect 314528 6264 314534 6276
rect 374086 6264 374092 6276
rect 374144 6264 374150 6316
rect 404262 6264 404268 6316
rect 404320 6304 404326 6316
rect 495894 6304 495900 6316
rect 404320 6276 495900 6304
rect 404320 6264 404326 6276
rect 495894 6264 495900 6276
rect 495952 6264 495958 6316
rect 269022 6196 269028 6248
rect 269080 6236 269086 6248
rect 311434 6236 311440 6248
rect 269080 6208 311440 6236
rect 269080 6196 269086 6208
rect 311434 6196 311440 6208
rect 311492 6196 311498 6248
rect 322842 6196 322848 6248
rect 322900 6236 322906 6248
rect 384758 6236 384764 6248
rect 322900 6208 384764 6236
rect 322900 6196 322906 6208
rect 384758 6196 384764 6208
rect 384816 6196 384822 6248
rect 407022 6196 407028 6248
rect 407080 6236 407086 6248
rect 499390 6236 499396 6248
rect 407080 6208 499396 6236
rect 407080 6196 407086 6208
rect 499390 6196 499396 6208
rect 499448 6196 499454 6248
rect 274542 6128 274548 6180
rect 274600 6168 274606 6180
rect 318518 6168 318524 6180
rect 274600 6140 318524 6168
rect 274600 6128 274606 6140
rect 318518 6128 318524 6140
rect 318576 6128 318582 6180
rect 324222 6128 324228 6180
rect 324280 6168 324286 6180
rect 387150 6168 387156 6180
rect 324280 6140 387156 6168
rect 324280 6128 324286 6140
rect 387150 6128 387156 6140
rect 387208 6128 387214 6180
rect 408310 6128 408316 6180
rect 408368 6168 408374 6180
rect 502978 6168 502984 6180
rect 408368 6140 502984 6168
rect 408368 6128 408374 6140
rect 502978 6128 502984 6140
rect 503036 6128 503042 6180
rect 382182 6060 382188 6112
rect 382240 6100 382246 6112
rect 466270 6100 466276 6112
rect 382240 6072 466276 6100
rect 382240 6060 382246 6072
rect 466270 6060 466276 6072
rect 466328 6060 466334 6112
rect 342898 5992 342904 6044
rect 342956 6032 342962 6044
rect 391842 6032 391848 6044
rect 342956 6004 391848 6032
rect 342956 5992 342962 6004
rect 391842 5992 391848 6004
rect 391900 5992 391906 6044
rect 393958 5516 393964 5568
rect 394016 5556 394022 5568
rect 396534 5556 396540 5568
rect 394016 5528 396540 5556
rect 394016 5516 394022 5528
rect 396534 5516 396540 5528
rect 396592 5516 396598 5568
rect 475378 5516 475384 5568
rect 475436 5556 475442 5568
rect 480530 5556 480536 5568
rect 475436 5528 480536 5556
rect 475436 5516 475442 5528
rect 480530 5516 480536 5528
rect 480588 5516 480594 5568
rect 486418 5516 486424 5568
rect 486476 5556 486482 5568
rect 487614 5556 487620 5568
rect 486476 5528 487620 5556
rect 486476 5516 486482 5528
rect 487614 5516 487620 5528
rect 487672 5516 487678 5568
rect 493318 5516 493324 5568
rect 493376 5556 493382 5568
rect 494698 5556 494704 5568
rect 493376 5528 494704 5556
rect 493376 5516 493382 5528
rect 494698 5516 494704 5528
rect 494756 5516 494762 5568
rect 512638 5516 512644 5568
rect 512696 5556 512702 5568
rect 513558 5556 513564 5568
rect 512696 5528 513564 5556
rect 512696 5516 512702 5528
rect 513558 5516 513564 5528
rect 513616 5516 513622 5568
rect 269758 5448 269764 5500
rect 269816 5488 269822 5500
rect 292574 5488 292580 5500
rect 269816 5460 292580 5488
rect 269816 5448 269822 5460
rect 292574 5448 292580 5460
rect 292632 5448 292638 5500
rect 354582 5448 354588 5500
rect 354640 5488 354646 5500
rect 427262 5488 427268 5500
rect 354640 5460 427268 5488
rect 354640 5448 354646 5460
rect 427262 5448 427268 5460
rect 427320 5448 427326 5500
rect 435910 5448 435916 5500
rect 435968 5488 435974 5500
rect 540790 5488 540796 5500
rect 435968 5460 540796 5488
rect 435968 5448 435974 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 268378 5380 268384 5432
rect 268436 5420 268442 5432
rect 297266 5420 297272 5432
rect 268436 5392 297272 5420
rect 268436 5380 268442 5392
rect 297266 5380 297272 5392
rect 297324 5380 297330 5432
rect 351822 5380 351828 5432
rect 351880 5420 351886 5432
rect 423766 5420 423772 5432
rect 351880 5392 423772 5420
rect 351880 5380 351886 5392
rect 423766 5380 423772 5392
rect 423824 5380 423830 5432
rect 438670 5380 438676 5432
rect 438728 5420 438734 5432
rect 544378 5420 544384 5432
rect 438728 5392 544384 5420
rect 438728 5380 438734 5392
rect 544378 5380 544384 5392
rect 544436 5380 544442 5432
rect 256602 5312 256608 5364
rect 256660 5352 256666 5364
rect 293678 5352 293684 5364
rect 256660 5324 293684 5352
rect 256660 5312 256666 5324
rect 293678 5312 293684 5324
rect 293736 5312 293742 5364
rect 304258 5312 304264 5364
rect 304316 5352 304322 5364
rect 310238 5352 310244 5364
rect 304316 5324 310244 5352
rect 304316 5312 304322 5324
rect 310238 5312 310244 5324
rect 310296 5312 310302 5364
rect 355870 5312 355876 5364
rect 355928 5352 355934 5364
rect 430850 5352 430856 5364
rect 355928 5324 430856 5352
rect 355928 5312 355934 5324
rect 430850 5312 430856 5324
rect 430908 5312 430914 5364
rect 444282 5312 444288 5364
rect 444340 5352 444346 5364
rect 551462 5352 551468 5364
rect 444340 5324 551468 5352
rect 444340 5312 444346 5324
rect 551462 5312 551468 5324
rect 551520 5312 551526 5364
rect 266998 5244 267004 5296
rect 267056 5284 267062 5296
rect 306742 5284 306748 5296
rect 267056 5256 306748 5284
rect 267056 5244 267062 5256
rect 306742 5244 306748 5256
rect 306800 5244 306806 5296
rect 307018 5244 307024 5296
rect 307076 5284 307082 5296
rect 346946 5284 346952 5296
rect 307076 5256 346952 5284
rect 307076 5244 307082 5256
rect 346946 5244 346952 5256
rect 347004 5244 347010 5296
rect 358630 5244 358636 5296
rect 358688 5284 358694 5296
rect 434438 5284 434444 5296
rect 358688 5256 434444 5284
rect 358688 5244 358694 5256
rect 434438 5244 434444 5256
rect 434496 5244 434502 5296
rect 441430 5244 441436 5296
rect 441488 5284 441494 5296
rect 547874 5284 547880 5296
rect 441488 5256 547880 5284
rect 441488 5244 441494 5256
rect 547874 5244 547880 5256
rect 547932 5244 547938 5296
rect 271782 5176 271788 5228
rect 271840 5216 271846 5228
rect 313826 5216 313832 5228
rect 271840 5188 313832 5216
rect 271840 5176 271846 5188
rect 313826 5176 313832 5188
rect 313884 5176 313890 5228
rect 364242 5176 364248 5228
rect 364300 5216 364306 5228
rect 441522 5216 441528 5228
rect 364300 5188 441528 5216
rect 364300 5176 364306 5188
rect 441522 5176 441528 5188
rect 441580 5176 441586 5228
rect 449802 5176 449808 5228
rect 449860 5216 449866 5228
rect 558546 5216 558552 5228
rect 449860 5188 558552 5216
rect 449860 5176 449866 5188
rect 558546 5176 558552 5188
rect 558604 5176 558610 5228
rect 271690 5108 271696 5160
rect 271748 5148 271754 5160
rect 315022 5148 315028 5160
rect 271748 5120 315028 5148
rect 271748 5108 271754 5120
rect 315022 5108 315028 5120
rect 315080 5108 315086 5160
rect 361390 5108 361396 5160
rect 361448 5148 361454 5160
rect 437934 5148 437940 5160
rect 361448 5120 437940 5148
rect 361448 5108 361454 5120
rect 437934 5108 437940 5120
rect 437992 5108 437998 5160
rect 447042 5108 447048 5160
rect 447100 5148 447106 5160
rect 554958 5148 554964 5160
rect 447100 5120 554964 5148
rect 447100 5108 447106 5120
rect 554958 5108 554964 5120
rect 555016 5108 555022 5160
rect 242158 5040 242164 5092
rect 242216 5080 242222 5092
rect 271230 5080 271236 5092
rect 242216 5052 271236 5080
rect 242216 5040 242222 5052
rect 271230 5040 271236 5052
rect 271288 5040 271294 5092
rect 281442 5040 281448 5092
rect 281500 5080 281506 5092
rect 327994 5080 328000 5092
rect 281500 5052 328000 5080
rect 281500 5040 281506 5052
rect 327994 5040 328000 5052
rect 328052 5040 328058 5092
rect 367002 5040 367008 5092
rect 367060 5080 367066 5092
rect 445018 5080 445024 5092
rect 367060 5052 445024 5080
rect 367060 5040 367066 5052
rect 445018 5040 445024 5052
rect 445076 5040 445082 5092
rect 452470 5040 452476 5092
rect 452528 5080 452534 5092
rect 562042 5080 562048 5092
rect 452528 5052 562048 5080
rect 452528 5040 452534 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 234430 4972 234436 5024
rect 234488 5012 234494 5024
rect 264146 5012 264152 5024
rect 234488 4984 264152 5012
rect 234488 4972 234494 4984
rect 264146 4972 264152 4984
rect 264204 4972 264210 5024
rect 267090 4972 267096 5024
rect 267148 5012 267154 5024
rect 267734 5012 267740 5024
rect 267148 4984 267740 5012
rect 267148 4972 267154 4984
rect 267734 4972 267740 4984
rect 267792 4972 267798 5024
rect 286962 4972 286968 5024
rect 287020 5012 287026 5024
rect 335078 5012 335084 5024
rect 287020 4984 335084 5012
rect 287020 4972 287026 4984
rect 335078 4972 335084 4984
rect 335136 4972 335142 5024
rect 372522 4972 372528 5024
rect 372580 5012 372586 5024
rect 452102 5012 452108 5024
rect 372580 4984 452108 5012
rect 372580 4972 372586 4984
rect 452102 4972 452108 4984
rect 452160 4972 452166 5024
rect 455322 4972 455328 5024
rect 455380 5012 455386 5024
rect 565630 5012 565636 5024
rect 455380 4984 565636 5012
rect 455380 4972 455386 4984
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 224218 4904 224224 4956
rect 224276 4944 224282 4956
rect 242894 4944 242900 4956
rect 224276 4916 242900 4944
rect 224276 4904 224282 4916
rect 242894 4904 242900 4916
rect 242952 4904 242958 4956
rect 250990 4904 250996 4956
rect 251048 4944 251054 4956
rect 285398 4944 285404 4956
rect 251048 4916 285404 4944
rect 251048 4904 251054 4916
rect 285398 4904 285404 4916
rect 285456 4904 285462 4956
rect 285490 4904 285496 4956
rect 285548 4944 285554 4956
rect 332686 4944 332692 4956
rect 285548 4916 332692 4944
rect 285548 4904 285554 4916
rect 332686 4904 332692 4916
rect 332744 4904 332750 4956
rect 369762 4904 369768 4956
rect 369820 4944 369826 4956
rect 448606 4944 448612 4956
rect 369820 4916 448612 4944
rect 369820 4904 369826 4916
rect 448606 4904 448612 4916
rect 448664 4904 448670 4956
rect 456610 4904 456616 4956
rect 456668 4944 456674 4956
rect 569126 4944 569132 4956
rect 456668 4916 569132 4944
rect 456668 4904 456674 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 213730 4836 213736 4888
rect 213788 4876 213794 4888
rect 235810 4876 235816 4888
rect 213788 4848 235816 4876
rect 213788 4836 213794 4848
rect 235810 4836 235816 4848
rect 235868 4836 235874 4888
rect 238018 4836 238024 4888
rect 238076 4876 238082 4888
rect 239306 4876 239312 4888
rect 238076 4848 239312 4876
rect 238076 4836 238082 4848
rect 239306 4836 239312 4848
rect 239364 4836 239370 4888
rect 253842 4836 253848 4888
rect 253900 4876 253906 4888
rect 290182 4876 290188 4888
rect 253900 4848 290188 4876
rect 253900 4836 253906 4848
rect 290182 4836 290188 4848
rect 290240 4836 290246 4888
rect 292482 4836 292488 4888
rect 292540 4876 292546 4888
rect 342162 4876 342168 4888
rect 292540 4848 342168 4876
rect 292540 4836 292546 4848
rect 342162 4836 342168 4848
rect 342220 4836 342226 4888
rect 375190 4836 375196 4888
rect 375248 4876 375254 4888
rect 455690 4876 455696 4888
rect 375248 4848 455696 4876
rect 375248 4836 375254 4848
rect 455690 4836 455696 4848
rect 455748 4836 455754 4888
rect 462130 4836 462136 4888
rect 462188 4876 462194 4888
rect 576302 4876 576308 4888
rect 462188 4848 576308 4876
rect 462188 4836 462194 4848
rect 576302 4836 576308 4848
rect 576360 4836 576366 4888
rect 227530 4768 227536 4820
rect 227588 4808 227594 4820
rect 253474 4808 253480 4820
rect 227588 4780 253480 4808
rect 227588 4768 227594 4780
rect 253474 4768 253480 4780
rect 253532 4768 253538 4820
rect 260742 4768 260748 4820
rect 260800 4808 260806 4820
rect 299658 4808 299664 4820
rect 260800 4780 299664 4808
rect 260800 4768 260806 4780
rect 299658 4768 299664 4780
rect 299716 4768 299722 4820
rect 303430 4768 303436 4820
rect 303488 4808 303494 4820
rect 357526 4808 357532 4820
rect 303488 4780 357532 4808
rect 303488 4768 303494 4780
rect 357526 4768 357532 4780
rect 357584 4768 357590 4820
rect 376570 4768 376576 4820
rect 376628 4808 376634 4820
rect 459186 4808 459192 4820
rect 376628 4780 459192 4808
rect 376628 4768 376634 4780
rect 459186 4768 459192 4780
rect 459244 4768 459250 4820
rect 459370 4768 459376 4820
rect 459428 4808 459434 4820
rect 572714 4808 572720 4820
rect 459428 4780 572720 4808
rect 459428 4768 459434 4780
rect 572714 4768 572720 4780
rect 572772 4768 572778 4820
rect 251818 4700 251824 4752
rect 251876 4740 251882 4752
rect 274818 4740 274824 4752
rect 251876 4712 274824 4740
rect 251876 4700 251882 4712
rect 274818 4700 274824 4712
rect 274876 4700 274882 4752
rect 289078 4700 289084 4752
rect 289136 4740 289142 4752
rect 289136 4712 296714 4740
rect 289136 4700 289142 4712
rect 276658 4632 276664 4684
rect 276716 4672 276722 4684
rect 296070 4672 296076 4684
rect 276716 4644 296076 4672
rect 276716 4632 276722 4644
rect 296070 4632 296076 4644
rect 296128 4632 296134 4684
rect 296686 4672 296714 4712
rect 349062 4700 349068 4752
rect 349120 4740 349126 4752
rect 420178 4740 420184 4752
rect 349120 4712 420184 4740
rect 349120 4700 349126 4712
rect 420178 4700 420184 4712
rect 420236 4700 420242 4752
rect 434622 4700 434628 4752
rect 434680 4740 434686 4752
rect 537202 4740 537208 4752
rect 434680 4712 537208 4740
rect 434680 4700 434686 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 307938 4672 307944 4684
rect 296686 4644 307944 4672
rect 307938 4632 307944 4644
rect 307996 4632 308002 4684
rect 346302 4632 346308 4684
rect 346360 4672 346366 4684
rect 416682 4672 416688 4684
rect 346360 4644 416688 4672
rect 346360 4632 346366 4644
rect 416682 4632 416688 4644
rect 416740 4632 416746 4684
rect 431862 4632 431868 4684
rect 431920 4672 431926 4684
rect 533706 4672 533712 4684
rect 431920 4644 533712 4672
rect 431920 4632 431926 4644
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 273898 4564 273904 4616
rect 273956 4604 273962 4616
rect 288986 4604 288992 4616
rect 273956 4576 288992 4604
rect 273956 4564 273962 4576
rect 288986 4564 288992 4576
rect 289044 4564 289050 4616
rect 343542 4564 343548 4616
rect 343600 4604 343606 4616
rect 413094 4604 413100 4616
rect 343600 4576 413100 4604
rect 343600 4564 343606 4576
rect 413094 4564 413100 4576
rect 413152 4564 413158 4616
rect 429102 4564 429108 4616
rect 429160 4604 429166 4616
rect 530118 4604 530124 4616
rect 429160 4576 530124 4604
rect 429160 4564 429166 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 262858 4496 262864 4548
rect 262916 4536 262922 4548
rect 278314 4536 278320 4548
rect 262916 4508 278320 4536
rect 262916 4496 262922 4508
rect 278314 4496 278320 4508
rect 278372 4496 278378 4548
rect 287698 4496 287704 4548
rect 287756 4536 287762 4548
rect 303154 4536 303160 4548
rect 287756 4508 303160 4536
rect 287756 4496 287762 4508
rect 303154 4496 303160 4508
rect 303212 4496 303218 4548
rect 337930 4496 337936 4548
rect 337988 4536 337994 4548
rect 406010 4536 406016 4548
rect 337988 4508 406016 4536
rect 337988 4496 337994 4508
rect 406010 4496 406016 4508
rect 406068 4496 406074 4548
rect 423582 4496 423588 4548
rect 423640 4536 423646 4548
rect 523034 4536 523040 4548
rect 423640 4508 523040 4536
rect 423640 4496 423646 4508
rect 523034 4496 523040 4508
rect 523092 4496 523098 4548
rect 340690 4428 340696 4480
rect 340748 4468 340754 4480
rect 409598 4468 409604 4480
rect 340748 4440 409604 4468
rect 340748 4428 340754 4440
rect 409598 4428 409604 4440
rect 409656 4428 409662 4480
rect 426342 4428 426348 4480
rect 426400 4468 426406 4480
rect 526622 4468 526628 4480
rect 426400 4440 526628 4468
rect 426400 4428 426406 4440
rect 526622 4428 526628 4440
rect 526680 4428 526686 4480
rect 244918 4360 244924 4412
rect 244976 4400 244982 4412
rect 249978 4400 249984 4412
rect 244976 4372 249984 4400
rect 244976 4360 244982 4372
rect 249978 4360 249984 4372
rect 250036 4360 250042 4412
rect 335170 4360 335176 4412
rect 335228 4400 335234 4412
rect 402514 4400 402520 4412
rect 335228 4372 402520 4400
rect 335228 4360 335234 4372
rect 402514 4360 402520 4372
rect 402572 4360 402578 4412
rect 420730 4360 420736 4412
rect 420788 4400 420794 4412
rect 519538 4400 519544 4412
rect 420788 4372 519544 4400
rect 420788 4360 420794 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 333882 4292 333888 4344
rect 333940 4332 333946 4344
rect 398926 4332 398932 4344
rect 333940 4304 398932 4332
rect 333940 4292 333946 4304
rect 398926 4292 398932 4304
rect 398984 4292 398990 4344
rect 418062 4292 418068 4344
rect 418120 4332 418126 4344
rect 515950 4332 515956 4344
rect 418120 4304 515956 4332
rect 418120 4292 418126 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 331122 4224 331128 4276
rect 331180 4264 331186 4276
rect 395338 4264 395344 4276
rect 331180 4236 395344 4264
rect 331180 4224 331186 4236
rect 395338 4224 395344 4236
rect 395396 4224 395402 4276
rect 415302 4224 415308 4276
rect 415360 4264 415366 4276
rect 512454 4264 512460 4276
rect 415360 4236 512460 4264
rect 415360 4224 415366 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 255958 4156 255964 4208
rect 256016 4196 256022 4208
rect 257062 4196 257068 4208
rect 256016 4168 257068 4196
rect 256016 4156 256022 4168
rect 257062 4156 257068 4168
rect 257120 4156 257126 4208
rect 318058 4156 318064 4208
rect 318116 4196 318122 4208
rect 320910 4196 320916 4208
rect 318116 4168 320916 4196
rect 318116 4156 318122 4168
rect 320910 4156 320916 4168
rect 320968 4156 320974 4208
rect 327718 4156 327724 4208
rect 327776 4196 327782 4208
rect 329190 4196 329196 4208
rect 327776 4168 329196 4196
rect 327776 4156 327782 4168
rect 329190 4156 329196 4168
rect 329248 4156 329254 4208
rect 522298 4156 522304 4208
rect 522356 4196 522362 4208
rect 524230 4196 524236 4208
rect 522356 4168 524236 4196
rect 522356 4156 522362 4168
rect 524230 4156 524236 4168
rect 524288 4156 524294 4208
rect 26510 4088 26516 4140
rect 26568 4128 26574 4140
rect 60734 4128 60740 4140
rect 26568 4100 60740 4128
rect 26568 4088 26574 4100
rect 60734 4088 60740 4100
rect 60792 4088 60798 4140
rect 168282 4088 168288 4140
rect 168340 4128 168346 4140
rect 171962 4128 171968 4140
rect 168340 4100 171968 4128
rect 168340 4088 168346 4100
rect 171962 4088 171968 4100
rect 172020 4088 172026 4140
rect 186130 4088 186136 4140
rect 186188 4128 186194 4140
rect 196802 4128 196808 4140
rect 186188 4100 196808 4128
rect 186188 4088 186194 4100
rect 196802 4088 196808 4100
rect 196860 4088 196866 4140
rect 204162 4088 204168 4140
rect 204220 4128 204226 4140
rect 221550 4128 221556 4140
rect 204220 4100 221556 4128
rect 204220 4088 204226 4100
rect 221550 4088 221556 4100
rect 221608 4088 221614 4140
rect 223482 4088 223488 4140
rect 223540 4128 223546 4140
rect 247586 4128 247592 4140
rect 223540 4100 247592 4128
rect 223540 4088 223546 4100
rect 247586 4088 247592 4100
rect 247644 4088 247650 4140
rect 248322 4088 248328 4140
rect 248380 4128 248386 4140
rect 283098 4128 283104 4140
rect 248380 4100 283104 4128
rect 248380 4088 248386 4100
rect 283098 4088 283104 4100
rect 283156 4088 283162 4140
rect 291102 4088 291108 4140
rect 291160 4128 291166 4140
rect 340966 4128 340972 4140
rect 291160 4100 340972 4128
rect 291160 4088 291166 4100
rect 340966 4088 340972 4100
rect 341024 4088 341030 4140
rect 347682 4088 347688 4140
rect 347740 4128 347746 4140
rect 350353 4131 350411 4137
rect 350353 4128 350365 4131
rect 347740 4100 350365 4128
rect 347740 4088 347746 4100
rect 350353 4097 350365 4100
rect 350399 4097 350411 4131
rect 350353 4091 350411 4097
rect 350442 4088 350448 4140
rect 350500 4128 350506 4140
rect 422570 4128 422576 4140
rect 350500 4100 422576 4128
rect 350500 4088 350506 4100
rect 422570 4088 422576 4100
rect 422628 4088 422634 4140
rect 424778 4088 424784 4140
rect 424836 4128 424842 4140
rect 424962 4128 424968 4140
rect 424836 4100 424968 4128
rect 424836 4088 424842 4100
rect 424962 4088 424968 4100
rect 425020 4088 425026 4140
rect 441338 4088 441344 4140
rect 441396 4128 441402 4140
rect 546678 4128 546684 4140
rect 441396 4100 546684 4128
rect 441396 4088 441402 4100
rect 546678 4088 546684 4100
rect 546736 4088 546742 4140
rect 574738 4088 574744 4140
rect 574796 4128 574802 4140
rect 577406 4128 577412 4140
rect 574796 4100 577412 4128
rect 574796 4088 574802 4100
rect 577406 4088 577412 4100
rect 577464 4088 577470 4140
rect 31021 4063 31079 4069
rect 31021 4029 31033 4063
rect 31067 4060 31079 4063
rect 31067 4032 55214 4060
rect 31067 4029 31079 4032
rect 31021 4023 31079 4029
rect 17034 3952 17040 4004
rect 17092 3992 17098 4004
rect 53834 3992 53840 4004
rect 17092 3964 53840 3992
rect 17092 3952 17098 3964
rect 53834 3952 53840 3964
rect 53892 3952 53898 4004
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 55186 3924 55214 4032
rect 182082 4020 182088 4072
rect 182140 4060 182146 4072
rect 190822 4060 190828 4072
rect 182140 4032 190828 4060
rect 182140 4020 182146 4032
rect 190822 4020 190828 4032
rect 190880 4020 190886 4072
rect 191650 4020 191656 4072
rect 191708 4060 191714 4072
rect 203886 4060 203892 4072
rect 191708 4032 203892 4060
rect 191708 4020 191714 4032
rect 203886 4020 203892 4032
rect 203944 4020 203950 4072
rect 205542 4020 205548 4072
rect 205600 4060 205606 4072
rect 223942 4060 223948 4072
rect 205600 4032 223948 4060
rect 205600 4020 205606 4032
rect 223942 4020 223948 4032
rect 224000 4020 224006 4072
rect 226150 4020 226156 4072
rect 226208 4060 226214 4072
rect 252370 4060 252376 4072
rect 226208 4032 252376 4060
rect 226208 4020 226214 4032
rect 252370 4020 252376 4032
rect 252428 4020 252434 4072
rect 252462 4020 252468 4072
rect 252520 4060 252526 4072
rect 287790 4060 287796 4072
rect 252520 4032 287796 4060
rect 252520 4020 252526 4032
rect 287790 4020 287796 4032
rect 287848 4020 287854 4072
rect 299382 4020 299388 4072
rect 299440 4060 299446 4072
rect 351638 4060 351644 4072
rect 299440 4032 351644 4060
rect 299440 4020 299446 4032
rect 351638 4020 351644 4032
rect 351696 4020 351702 4072
rect 353202 4020 353208 4072
rect 353260 4060 353266 4072
rect 426158 4060 426164 4072
rect 353260 4032 426164 4060
rect 353260 4020 353266 4032
rect 426158 4020 426164 4032
rect 426216 4020 426222 4072
rect 442902 4020 442908 4072
rect 442960 4060 442966 4072
rect 550266 4060 550272 4072
rect 442960 4032 550272 4060
rect 442960 4020 442966 4032
rect 550266 4020 550272 4032
rect 550324 4020 550330 4072
rect 74721 3995 74779 4001
rect 74721 3961 74733 3995
rect 74767 3992 74779 3995
rect 81434 3992 81440 4004
rect 74767 3964 81440 3992
rect 74767 3961 74779 3964
rect 74721 3955 74779 3961
rect 81434 3952 81440 3964
rect 81492 3952 81498 4004
rect 161290 3952 161296 4004
rect 161348 3992 161354 4004
rect 163682 3992 163688 4004
rect 161348 3964 163688 3992
rect 161348 3952 161354 3964
rect 163682 3952 163688 3964
rect 163740 3952 163746 4004
rect 169018 3952 169024 4004
rect 169076 3992 169082 4004
rect 173158 3992 173164 4004
rect 169076 3964 173164 3992
rect 169076 3952 169082 3964
rect 173158 3952 173164 3964
rect 173216 3952 173222 4004
rect 179322 3952 179328 4004
rect 179380 3992 179386 4004
rect 187326 3992 187332 4004
rect 179380 3964 187332 3992
rect 179380 3952 179386 3964
rect 187326 3952 187332 3964
rect 187384 3952 187390 4004
rect 190362 3952 190368 4004
rect 190420 3992 190426 4004
rect 202598 3992 202604 4004
rect 190420 3964 202604 3992
rect 190420 3952 190426 3964
rect 202598 3952 202604 3964
rect 202656 3952 202662 4004
rect 202690 3952 202696 4004
rect 202748 3992 202754 4004
rect 220446 3992 220452 4004
rect 202748 3964 220452 3992
rect 202748 3952 202754 3964
rect 220446 3952 220452 3964
rect 220504 3952 220510 4004
rect 220630 3952 220636 4004
rect 220688 3992 220694 4004
rect 245194 3992 245200 4004
rect 220688 3964 245200 3992
rect 220688 3952 220694 3964
rect 245194 3952 245200 3964
rect 245252 3952 245258 4004
rect 249702 3952 249708 4004
rect 249760 3992 249766 4004
rect 284294 3992 284300 4004
rect 249760 3964 284300 3992
rect 249760 3952 249766 3964
rect 284294 3952 284300 3964
rect 284352 3952 284358 4004
rect 296622 3952 296628 4004
rect 296680 3992 296686 4004
rect 348050 3992 348056 4004
rect 296680 3964 348056 3992
rect 296680 3952 296686 3964
rect 348050 3952 348056 3964
rect 348108 3952 348114 4004
rect 358630 3952 358636 4004
rect 358688 3992 358694 4004
rect 358909 3995 358967 4001
rect 358688 3964 358860 3992
rect 358688 3952 358694 3964
rect 56594 3924 56600 3936
rect 20680 3896 50384 3924
rect 55186 3896 56600 3924
rect 20680 3884 20686 3896
rect 11146 3816 11152 3868
rect 11204 3856 11210 3868
rect 49694 3856 49700 3868
rect 11204 3828 49700 3856
rect 11204 3816 11210 3828
rect 49694 3816 49700 3828
rect 49752 3816 49758 3868
rect 50356 3856 50384 3896
rect 56594 3884 56600 3896
rect 56652 3884 56658 3936
rect 69106 3884 69112 3936
rect 69164 3924 69170 3936
rect 91186 3924 91192 3936
rect 69164 3896 91192 3924
rect 69164 3884 69170 3896
rect 91186 3884 91192 3896
rect 91244 3884 91250 3936
rect 177942 3884 177948 3936
rect 178000 3924 178006 3936
rect 186130 3924 186136 3936
rect 178000 3896 186136 3924
rect 178000 3884 178006 3896
rect 186130 3884 186136 3896
rect 186188 3884 186194 3936
rect 188890 3884 188896 3936
rect 188948 3924 188954 3936
rect 200298 3924 200304 3936
rect 188948 3896 200304 3924
rect 188948 3884 188954 3896
rect 200298 3884 200304 3896
rect 200356 3884 200362 3936
rect 205450 3884 205456 3936
rect 205508 3924 205514 3936
rect 222746 3924 222752 3936
rect 205508 3896 222752 3924
rect 205508 3884 205514 3896
rect 222746 3884 222752 3896
rect 222804 3884 222810 3936
rect 223390 3884 223396 3936
rect 223448 3924 223454 3936
rect 248782 3924 248788 3936
rect 223448 3896 248788 3924
rect 223448 3884 223454 3896
rect 248782 3884 248788 3896
rect 248840 3884 248846 3936
rect 251082 3884 251088 3936
rect 251140 3924 251146 3936
rect 286594 3924 286600 3936
rect 251140 3896 286600 3924
rect 251140 3884 251146 3896
rect 286594 3884 286600 3896
rect 286652 3884 286658 3936
rect 303522 3884 303528 3936
rect 303580 3924 303586 3936
rect 358722 3924 358728 3936
rect 303580 3896 358728 3924
rect 303580 3884 303586 3896
rect 358722 3884 358728 3896
rect 358780 3884 358786 3936
rect 358832 3924 358860 3964
rect 358909 3961 358921 3995
rect 358955 3992 358967 3995
rect 429654 3992 429660 4004
rect 358955 3964 429660 3992
rect 358955 3961 358967 3964
rect 358909 3955 358967 3961
rect 429654 3952 429660 3964
rect 429712 3952 429718 4004
rect 448422 3952 448428 4004
rect 448480 3992 448486 4004
rect 557350 3992 557356 4004
rect 448480 3964 557356 3992
rect 448480 3952 448486 3964
rect 557350 3952 557356 3964
rect 557408 3952 557414 4004
rect 433242 3924 433248 3936
rect 358832 3896 433248 3924
rect 433242 3884 433248 3896
rect 433300 3884 433306 3936
rect 445570 3884 445576 3936
rect 445628 3924 445634 3936
rect 553762 3924 553768 3936
rect 445628 3896 553768 3924
rect 445628 3884 445634 3896
rect 553762 3884 553768 3896
rect 553820 3884 553826 3936
rect 57057 3859 57115 3865
rect 50356 3828 55214 3856
rect 12342 3748 12348 3800
rect 12400 3788 12406 3800
rect 12400 3760 45554 3788
rect 12400 3748 12406 3760
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 42797 3723 42855 3729
rect 42797 3720 42809 3723
rect 7708 3692 42809 3720
rect 7708 3680 7714 3692
rect 42797 3689 42809 3692
rect 42843 3689 42855 3723
rect 42797 3683 42855 3689
rect 2866 3612 2872 3664
rect 2924 3652 2930 3664
rect 42886 3652 42892 3664
rect 2924 3624 42892 3652
rect 2924 3612 2930 3624
rect 42886 3612 42892 3624
rect 42944 3612 42950 3664
rect 45526 3652 45554 3760
rect 55186 3720 55214 3828
rect 57057 3825 57069 3859
rect 57103 3856 57115 3859
rect 64138 3856 64144 3868
rect 57103 3828 64144 3856
rect 57103 3825 57115 3828
rect 57057 3819 57115 3825
rect 64138 3816 64144 3828
rect 64196 3816 64202 3868
rect 65518 3816 65524 3868
rect 65576 3856 65582 3868
rect 89714 3856 89720 3868
rect 65576 3828 89720 3856
rect 65576 3816 65582 3828
rect 89714 3816 89720 3828
rect 89772 3816 89778 3868
rect 180702 3816 180708 3868
rect 180760 3856 180766 3868
rect 189718 3856 189724 3868
rect 180760 3828 189724 3856
rect 180760 3816 180766 3828
rect 189718 3816 189724 3828
rect 189776 3816 189782 3868
rect 191742 3816 191748 3868
rect 191800 3856 191806 3868
rect 205082 3856 205088 3868
rect 191800 3828 205088 3856
rect 191800 3816 191806 3828
rect 205082 3816 205088 3828
rect 205140 3816 205146 3868
rect 206830 3816 206836 3868
rect 206888 3856 206894 3868
rect 225138 3856 225144 3868
rect 206888 3828 225144 3856
rect 206888 3816 206894 3828
rect 225138 3816 225144 3828
rect 225196 3816 225202 3868
rect 227622 3816 227628 3868
rect 227680 3856 227686 3868
rect 254670 3856 254676 3868
rect 227680 3828 254676 3856
rect 227680 3816 227686 3828
rect 254670 3816 254676 3828
rect 254728 3816 254734 3868
rect 255222 3816 255228 3868
rect 255280 3856 255286 3868
rect 291378 3856 291384 3868
rect 255280 3828 291384 3856
rect 255280 3816 255286 3828
rect 291378 3816 291384 3828
rect 291436 3816 291442 3868
rect 300762 3816 300768 3868
rect 300820 3856 300826 3868
rect 355226 3856 355232 3868
rect 300820 3828 355232 3856
rect 300820 3816 300826 3828
rect 355226 3816 355232 3828
rect 355284 3816 355290 3868
rect 355962 3816 355968 3868
rect 356020 3856 356026 3868
rect 358909 3859 358967 3865
rect 358909 3856 358921 3859
rect 356020 3828 358921 3856
rect 356020 3816 356026 3828
rect 358909 3825 358921 3828
rect 358955 3825 358967 3859
rect 358909 3819 358967 3825
rect 361482 3816 361488 3868
rect 361540 3856 361546 3868
rect 436738 3856 436744 3868
rect 361540 3828 436744 3856
rect 361540 3816 361546 3828
rect 436738 3816 436744 3828
rect 436796 3816 436802 3868
rect 451182 3816 451188 3868
rect 451240 3856 451246 3868
rect 560846 3856 560852 3868
rect 451240 3828 560852 3856
rect 451240 3816 451246 3828
rect 560846 3816 560852 3828
rect 560904 3816 560910 3868
rect 56042 3748 56048 3800
rect 56100 3788 56106 3800
rect 56502 3788 56508 3800
rect 56100 3760 56508 3788
rect 56100 3748 56106 3760
rect 56502 3748 56508 3760
rect 56560 3748 56566 3800
rect 61930 3748 61936 3800
rect 61988 3788 61994 3800
rect 87046 3788 87052 3800
rect 61988 3760 87052 3788
rect 61988 3748 61994 3760
rect 87046 3748 87052 3760
rect 87104 3748 87110 3800
rect 183462 3748 183468 3800
rect 183520 3788 183526 3800
rect 193214 3788 193220 3800
rect 183520 3760 193220 3788
rect 183520 3748 183526 3760
rect 193214 3748 193220 3760
rect 193272 3748 193278 3800
rect 194502 3748 194508 3800
rect 194560 3788 194566 3800
rect 208578 3788 208584 3800
rect 194560 3760 208584 3788
rect 194560 3748 194566 3760
rect 208578 3748 208584 3760
rect 208636 3748 208642 3800
rect 211062 3748 211068 3800
rect 211120 3788 211126 3800
rect 231026 3788 231032 3800
rect 211120 3760 231032 3788
rect 211120 3748 211126 3760
rect 231026 3748 231032 3760
rect 231084 3748 231090 3800
rect 231762 3748 231768 3800
rect 231820 3788 231826 3800
rect 259454 3788 259460 3800
rect 231820 3760 259460 3788
rect 231820 3748 231826 3760
rect 259454 3748 259460 3760
rect 259512 3748 259518 3800
rect 262122 3748 262128 3800
rect 262180 3788 262186 3800
rect 301958 3788 301964 3800
rect 262180 3760 301964 3788
rect 262180 3748 262186 3760
rect 301958 3748 301964 3760
rect 302016 3748 302022 3800
rect 306282 3748 306288 3800
rect 306340 3788 306346 3800
rect 362310 3788 362316 3800
rect 306340 3760 362316 3788
rect 306340 3748 306346 3760
rect 362310 3748 362316 3760
rect 362368 3748 362374 3800
rect 362862 3748 362868 3800
rect 362920 3788 362926 3800
rect 440326 3788 440332 3800
rect 362920 3760 440332 3788
rect 362920 3748 362926 3760
rect 440326 3748 440332 3760
rect 440384 3748 440390 3800
rect 453942 3748 453948 3800
rect 454000 3788 454006 3800
rect 564434 3788 564440 3800
rect 454000 3760 564440 3788
rect 454000 3748 454006 3760
rect 564434 3748 564440 3760
rect 564492 3748 564498 3800
rect 56686 3720 56692 3732
rect 55186 3692 56692 3720
rect 56686 3680 56692 3692
rect 56744 3680 56750 3732
rect 58434 3680 58440 3732
rect 58492 3720 58498 3732
rect 84286 3720 84292 3732
rect 58492 3692 84292 3720
rect 58492 3680 58498 3692
rect 84286 3680 84292 3692
rect 84344 3680 84350 3732
rect 179230 3680 179236 3732
rect 179288 3720 179294 3732
rect 188522 3720 188528 3732
rect 179288 3692 188528 3720
rect 179288 3680 179294 3692
rect 188522 3680 188528 3692
rect 188580 3680 188586 3732
rect 188982 3680 188988 3732
rect 189040 3720 189046 3732
rect 201494 3720 201500 3732
rect 189040 3692 201500 3720
rect 189040 3680 189046 3692
rect 201494 3680 201500 3692
rect 201552 3680 201558 3732
rect 206922 3680 206928 3732
rect 206980 3720 206986 3732
rect 226334 3720 226340 3732
rect 206980 3692 226340 3720
rect 206980 3680 206986 3692
rect 226334 3680 226340 3692
rect 226392 3680 226398 3732
rect 230382 3680 230388 3732
rect 230440 3720 230446 3732
rect 258258 3720 258264 3732
rect 230440 3692 258264 3720
rect 230440 3680 230446 3692
rect 258258 3680 258264 3692
rect 258316 3680 258322 3732
rect 259362 3680 259368 3732
rect 259420 3720 259426 3732
rect 298462 3720 298468 3732
rect 259420 3692 298468 3720
rect 259420 3680 259426 3692
rect 298462 3680 298468 3692
rect 298520 3680 298526 3732
rect 311802 3680 311808 3732
rect 311860 3720 311866 3732
rect 369394 3720 369400 3732
rect 311860 3692 369400 3720
rect 311860 3680 311866 3692
rect 369394 3680 369400 3692
rect 369452 3680 369458 3732
rect 371142 3680 371148 3732
rect 371200 3720 371206 3732
rect 450906 3720 450912 3732
rect 371200 3692 450912 3720
rect 371200 3680 371206 3692
rect 450906 3680 450912 3692
rect 450964 3680 450970 3732
rect 456702 3680 456708 3732
rect 456760 3720 456766 3732
rect 568022 3720 568028 3732
rect 456760 3692 568028 3720
rect 456760 3680 456766 3692
rect 568022 3680 568028 3692
rect 568080 3680 568086 3732
rect 49786 3652 49792 3664
rect 45526 3624 49792 3652
rect 49786 3612 49792 3624
rect 49844 3612 49850 3664
rect 54938 3612 54944 3664
rect 54996 3652 55002 3664
rect 74721 3655 74779 3661
rect 74721 3652 74733 3655
rect 54996 3624 74733 3652
rect 54996 3612 55002 3624
rect 74721 3621 74733 3624
rect 74767 3621 74779 3655
rect 78674 3652 78680 3664
rect 74721 3615 74779 3621
rect 74828 3624 78680 3652
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 45646 3584 45652 3596
rect 5316 3556 45652 3584
rect 5316 3544 5322 3556
rect 45646 3544 45652 3556
rect 45704 3544 45710 3596
rect 51350 3544 51356 3596
rect 51408 3584 51414 3596
rect 74828 3584 74856 3624
rect 78674 3612 78680 3624
rect 78732 3612 78738 3664
rect 85666 3612 85672 3664
rect 85724 3652 85730 3664
rect 86770 3652 86776 3664
rect 85724 3624 86776 3652
rect 85724 3612 85730 3624
rect 86770 3612 86776 3624
rect 86828 3612 86834 3664
rect 170950 3612 170956 3664
rect 171008 3652 171014 3664
rect 175458 3652 175464 3664
rect 171008 3624 175464 3652
rect 171008 3612 171014 3624
rect 175458 3612 175464 3624
rect 175516 3612 175522 3664
rect 176562 3612 176568 3664
rect 176620 3652 176626 3664
rect 183738 3652 183744 3664
rect 176620 3624 183744 3652
rect 176620 3612 176626 3624
rect 183738 3612 183744 3624
rect 183796 3612 183802 3664
rect 184750 3612 184756 3664
rect 184808 3652 184814 3664
rect 195606 3652 195612 3664
rect 184808 3624 195612 3652
rect 184808 3612 184814 3624
rect 195606 3612 195612 3624
rect 195664 3612 195670 3664
rect 195790 3612 195796 3664
rect 195848 3652 195854 3664
rect 209774 3652 209780 3664
rect 195848 3624 209780 3652
rect 195848 3612 195854 3624
rect 209774 3612 209780 3624
rect 209832 3612 209838 3664
rect 212350 3612 212356 3664
rect 212408 3652 212414 3664
rect 232222 3652 232228 3664
rect 212408 3624 232228 3652
rect 212408 3612 212414 3624
rect 232222 3612 232228 3624
rect 232280 3612 232286 3664
rect 234522 3612 234528 3664
rect 234580 3652 234586 3664
rect 262950 3652 262956 3664
rect 234580 3624 262956 3652
rect 234580 3612 234586 3624
rect 262950 3612 262956 3624
rect 263008 3612 263014 3664
rect 264882 3612 264888 3664
rect 264940 3652 264946 3664
rect 305546 3652 305552 3664
rect 264940 3624 305552 3652
rect 264940 3612 264946 3624
rect 305546 3612 305552 3624
rect 305604 3612 305610 3664
rect 308950 3612 308956 3664
rect 309008 3652 309014 3664
rect 365806 3652 365812 3664
rect 309008 3624 365812 3652
rect 309008 3612 309014 3624
rect 365806 3612 365812 3624
rect 365864 3612 365870 3664
rect 368382 3612 368388 3664
rect 368440 3652 368446 3664
rect 447410 3652 447416 3664
rect 368440 3624 447416 3652
rect 368440 3612 368446 3624
rect 447410 3612 447416 3624
rect 447468 3612 447474 3664
rect 448514 3612 448520 3664
rect 448572 3652 448578 3664
rect 449802 3652 449808 3664
rect 448572 3624 449808 3652
rect 448572 3612 448578 3624
rect 449802 3612 449808 3624
rect 449860 3612 449866 3664
rect 459462 3612 459468 3664
rect 459520 3652 459526 3664
rect 571518 3652 571524 3664
rect 459520 3624 571524 3652
rect 459520 3612 459526 3624
rect 571518 3612 571524 3624
rect 571576 3612 571582 3664
rect 76098 3584 76104 3596
rect 51408 3556 74856 3584
rect 74920 3556 76104 3584
rect 51408 3544 51414 3556
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 1728 3488 41644 3516
rect 1728 3476 1734 3488
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 41506 3448 41512 3460
rect 624 3420 41512 3448
rect 624 3408 630 3420
rect 41506 3408 41512 3420
rect 41564 3408 41570 3460
rect 41616 3448 41644 3488
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 42797 3519 42855 3525
rect 42797 3485 42809 3519
rect 42843 3516 42855 3519
rect 46934 3516 46940 3528
rect 42843 3488 46940 3516
rect 42843 3485 42855 3488
rect 42797 3479 42855 3485
rect 46934 3476 46940 3488
rect 46992 3476 46998 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 53650 3516 53656 3528
rect 52604 3488 53656 3516
rect 52604 3476 52610 3488
rect 53650 3476 53656 3488
rect 53708 3476 53714 3528
rect 53745 3519 53803 3525
rect 53745 3485 53757 3519
rect 53791 3516 53803 3519
rect 74920 3516 74948 3556
rect 76098 3544 76104 3556
rect 76156 3544 76162 3596
rect 93946 3544 93952 3596
rect 94004 3584 94010 3596
rect 95050 3584 95056 3596
rect 94004 3556 95056 3584
rect 94004 3544 94010 3556
rect 95050 3544 95056 3556
rect 95108 3544 95114 3596
rect 161382 3544 161388 3596
rect 161440 3584 161446 3596
rect 162486 3584 162492 3596
rect 161440 3556 162492 3584
rect 161440 3544 161446 3556
rect 162486 3544 162492 3556
rect 162544 3544 162550 3596
rect 165430 3544 165436 3596
rect 165488 3584 165494 3596
rect 169570 3584 169576 3596
rect 165488 3556 169576 3584
rect 165488 3544 165494 3556
rect 169570 3544 169576 3556
rect 169628 3544 169634 3596
rect 172330 3544 172336 3596
rect 172388 3584 172394 3596
rect 177850 3584 177856 3596
rect 172388 3556 177856 3584
rect 172388 3544 172394 3556
rect 177850 3544 177856 3556
rect 177908 3544 177914 3596
rect 181990 3544 181996 3596
rect 182048 3584 182054 3596
rect 192018 3584 192024 3596
rect 182048 3556 192024 3584
rect 182048 3544 182054 3556
rect 192018 3544 192024 3556
rect 192076 3544 192082 3596
rect 193030 3544 193036 3596
rect 193088 3584 193094 3596
rect 207382 3584 207388 3596
rect 193088 3556 207388 3584
rect 193088 3544 193094 3556
rect 207382 3544 207388 3556
rect 207440 3544 207446 3596
rect 212442 3544 212448 3596
rect 212500 3584 212506 3596
rect 233418 3584 233424 3596
rect 212500 3556 233424 3584
rect 212500 3544 212506 3556
rect 233418 3544 233424 3556
rect 233476 3544 233482 3596
rect 241330 3544 241336 3596
rect 241388 3584 241394 3596
rect 273622 3584 273628 3596
rect 241388 3556 273628 3584
rect 241388 3544 241394 3556
rect 273622 3544 273628 3556
rect 273680 3544 273686 3596
rect 275922 3544 275928 3596
rect 275980 3584 275986 3596
rect 319714 3584 319720 3596
rect 275980 3556 319720 3584
rect 275980 3544 275986 3556
rect 319714 3544 319720 3556
rect 319772 3544 319778 3596
rect 320082 3544 320088 3596
rect 320140 3584 320146 3596
rect 379974 3584 379980 3596
rect 320140 3556 379980 3584
rect 320140 3544 320146 3556
rect 379974 3544 379980 3556
rect 380032 3544 380038 3596
rect 380802 3544 380808 3596
rect 380860 3584 380866 3596
rect 465166 3584 465172 3596
rect 380860 3556 465172 3584
rect 380860 3544 380866 3556
rect 465166 3544 465172 3556
rect 465224 3544 465230 3596
rect 466178 3544 466184 3596
rect 466236 3584 466242 3596
rect 582190 3584 582196 3596
rect 466236 3556 582196 3584
rect 466236 3544 466242 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 53791 3488 74948 3516
rect 53791 3485 53803 3488
rect 53745 3479 53803 3485
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 77386 3476 77392 3528
rect 77444 3516 77450 3528
rect 78490 3516 78496 3528
rect 77444 3488 78496 3516
rect 77444 3476 77450 3488
rect 78490 3476 78496 3488
rect 78548 3476 78554 3528
rect 80882 3476 80888 3528
rect 80940 3516 80946 3528
rect 81342 3516 81348 3528
rect 80940 3488 81348 3516
rect 80940 3476 80946 3488
rect 81342 3476 81348 3488
rect 81400 3476 81406 3528
rect 82078 3476 82084 3528
rect 82136 3516 82142 3528
rect 82722 3516 82728 3528
rect 82136 3488 82728 3516
rect 82136 3476 82142 3488
rect 82722 3476 82728 3488
rect 82780 3476 82786 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 84102 3516 84108 3528
rect 83332 3488 84108 3516
rect 83332 3476 83338 3488
rect 84102 3476 84108 3488
rect 84160 3476 84166 3528
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 85482 3516 85488 3528
rect 84528 3488 85488 3516
rect 84528 3476 84534 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 89622 3516 89628 3528
rect 89220 3488 89628 3516
rect 89220 3476 89226 3488
rect 89622 3476 89628 3488
rect 89680 3476 89686 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 92382 3516 92388 3528
rect 91612 3488 92388 3516
rect 91612 3476 91618 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 102042 3516 102048 3528
rect 101088 3488 102048 3516
rect 101088 3476 101094 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 102226 3476 102232 3528
rect 102284 3516 102290 3528
rect 103238 3516 103244 3528
rect 102284 3488 103244 3516
rect 102284 3476 102290 3488
rect 103238 3476 103244 3488
rect 103296 3476 103302 3528
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 106182 3516 106188 3528
rect 105780 3488 106188 3516
rect 105780 3476 105786 3488
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 110322 3516 110328 3528
rect 109368 3488 110328 3516
rect 109368 3476 109374 3488
rect 110322 3476 110328 3488
rect 110380 3476 110386 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111518 3516 111524 3528
rect 110564 3488 111524 3516
rect 110564 3476 110570 3488
rect 111518 3476 111524 3488
rect 111576 3476 111582 3528
rect 114002 3476 114008 3528
rect 114060 3516 114066 3528
rect 114462 3516 114468 3528
rect 114060 3488 114468 3516
rect 114060 3476 114066 3488
rect 114462 3476 114468 3488
rect 114520 3476 114526 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 116394 3476 116400 3528
rect 116452 3516 116458 3528
rect 117222 3516 117228 3528
rect 116452 3488 117228 3516
rect 116452 3476 116458 3488
rect 117222 3476 117228 3488
rect 117280 3476 117286 3528
rect 117590 3476 117596 3528
rect 117648 3516 117654 3528
rect 118602 3516 118608 3528
rect 117648 3488 118608 3516
rect 117648 3476 117654 3488
rect 118602 3476 118608 3488
rect 118660 3476 118666 3528
rect 118786 3476 118792 3528
rect 118844 3516 118850 3528
rect 119982 3516 119988 3528
rect 118844 3488 119988 3516
rect 118844 3476 118850 3488
rect 119982 3476 119988 3488
rect 120040 3476 120046 3528
rect 122282 3476 122288 3528
rect 122340 3516 122346 3528
rect 122742 3516 122748 3528
rect 122340 3488 122748 3516
rect 122340 3476 122346 3488
rect 122742 3476 122748 3488
rect 122800 3476 122806 3528
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126882 3516 126888 3528
rect 125928 3488 126888 3516
rect 125928 3476 125934 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128262 3516 128268 3528
rect 127032 3488 128268 3516
rect 127032 3476 127038 3488
rect 128262 3476 128268 3488
rect 128320 3476 128326 3528
rect 130562 3476 130568 3528
rect 130620 3516 130626 3528
rect 131022 3516 131028 3528
rect 130620 3488 131028 3516
rect 130620 3476 130626 3488
rect 131022 3476 131028 3488
rect 131080 3476 131086 3528
rect 132954 3476 132960 3528
rect 133012 3516 133018 3528
rect 133782 3516 133788 3528
rect 133012 3488 133788 3516
rect 133012 3476 133018 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
rect 134150 3476 134156 3528
rect 134208 3516 134214 3528
rect 135162 3516 135168 3528
rect 134208 3488 135168 3516
rect 134208 3476 134214 3488
rect 135162 3476 135168 3488
rect 135220 3476 135226 3528
rect 135254 3476 135260 3528
rect 135312 3516 135318 3528
rect 137278 3516 137284 3528
rect 135312 3488 137284 3516
rect 135312 3476 135318 3488
rect 137278 3476 137284 3488
rect 137336 3476 137342 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 140682 3516 140688 3528
rect 140096 3488 140688 3516
rect 140096 3476 140102 3488
rect 140682 3476 140688 3488
rect 140740 3476 140746 3528
rect 142430 3476 142436 3528
rect 142488 3516 142494 3528
rect 143442 3516 143448 3528
rect 142488 3488 143448 3516
rect 142488 3476 142494 3488
rect 143442 3476 143448 3488
rect 143500 3476 143506 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
rect 150434 3516 150440 3528
rect 149572 3488 150440 3516
rect 149572 3476 149578 3488
rect 150434 3476 150440 3488
rect 150492 3476 150498 3528
rect 153286 3476 153292 3528
rect 153344 3516 153350 3528
rect 154206 3516 154212 3528
rect 153344 3488 154212 3516
rect 153344 3476 153350 3488
rect 154206 3476 154212 3488
rect 154264 3476 154270 3528
rect 155954 3476 155960 3528
rect 156012 3516 156018 3528
rect 156598 3516 156604 3528
rect 156012 3488 156604 3516
rect 156012 3476 156018 3488
rect 156598 3476 156604 3488
rect 156656 3476 156662 3528
rect 157242 3476 157248 3528
rect 157300 3516 157306 3528
rect 157794 3516 157800 3528
rect 157300 3488 157800 3516
rect 157300 3476 157306 3488
rect 157794 3476 157800 3488
rect 157852 3476 157858 3528
rect 158438 3476 158444 3528
rect 158496 3516 158502 3528
rect 158898 3516 158904 3528
rect 158496 3488 158904 3516
rect 158496 3476 158502 3488
rect 158898 3476 158904 3488
rect 158956 3476 158962 3528
rect 160002 3476 160008 3528
rect 160060 3516 160066 3528
rect 161290 3516 161296 3528
rect 160060 3488 161296 3516
rect 160060 3476 160066 3488
rect 161290 3476 161296 3488
rect 161348 3476 161354 3528
rect 164142 3476 164148 3528
rect 164200 3516 164206 3528
rect 167178 3516 167184 3528
rect 164200 3488 167184 3516
rect 164200 3476 164206 3488
rect 167178 3476 167184 3488
rect 167236 3476 167242 3528
rect 169662 3476 169668 3528
rect 169720 3516 169726 3528
rect 174262 3516 174268 3528
rect 169720 3488 174268 3516
rect 169720 3476 169726 3488
rect 174262 3476 174268 3488
rect 174320 3476 174326 3528
rect 187602 3476 187608 3528
rect 187660 3516 187666 3528
rect 199102 3516 199108 3528
rect 187660 3488 199108 3516
rect 187660 3476 187666 3488
rect 199102 3476 199108 3488
rect 199160 3476 199166 3528
rect 199930 3476 199936 3528
rect 199988 3516 199994 3528
rect 216858 3516 216864 3528
rect 199988 3488 216864 3516
rect 199988 3476 199994 3488
rect 216858 3476 216864 3488
rect 216916 3476 216922 3528
rect 217962 3476 217968 3528
rect 218020 3516 218026 3528
rect 240502 3516 240508 3528
rect 218020 3488 240508 3516
rect 218020 3476 218026 3488
rect 240502 3476 240508 3488
rect 240560 3476 240566 3528
rect 241422 3476 241428 3528
rect 241480 3516 241486 3528
rect 272426 3516 272432 3528
rect 241480 3488 272432 3516
rect 241480 3476 241486 3488
rect 272426 3476 272432 3488
rect 272484 3476 272490 3528
rect 273162 3476 273168 3528
rect 273220 3516 273226 3528
rect 316218 3516 316224 3528
rect 273220 3488 316224 3516
rect 273220 3476 273226 3488
rect 316218 3476 316224 3488
rect 316276 3476 316282 3528
rect 317414 3476 317420 3528
rect 317472 3516 317478 3528
rect 376478 3516 376484 3528
rect 317472 3488 376484 3516
rect 317472 3476 317478 3488
rect 376478 3476 376484 3488
rect 376536 3476 376542 3528
rect 376662 3476 376668 3528
rect 376720 3516 376726 3528
rect 458082 3516 458088 3528
rect 376720 3488 458088 3516
rect 376720 3476 376726 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 462222 3476 462228 3528
rect 462280 3516 462286 3528
rect 575106 3516 575112 3528
rect 462280 3488 575112 3516
rect 462280 3476 462286 3488
rect 575106 3476 575112 3488
rect 575164 3476 575170 3528
rect 42886 3448 42892 3460
rect 41616 3420 42892 3448
rect 42886 3408 42892 3420
rect 42944 3408 42950 3460
rect 44266 3408 44272 3460
rect 44324 3448 44330 3460
rect 44324 3420 66668 3448
rect 44324 3408 44330 3420
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 9582 3380 9588 3392
rect 8812 3352 9588 3380
rect 8812 3340 8818 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 16482 3380 16488 3392
rect 15988 3352 16488 3380
rect 15988 3340 15994 3352
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 19242 3380 19248 3392
rect 18288 3352 19248 3380
rect 18288 3340 18294 3352
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 24210 3340 24216 3392
rect 24268 3380 24274 3392
rect 24762 3380 24768 3392
rect 24268 3352 24768 3380
rect 24268 3340 24274 3352
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 25314 3340 25320 3392
rect 25372 3380 25378 3392
rect 26142 3380 26148 3392
rect 25372 3352 26148 3380
rect 25372 3340 25378 3352
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 28902 3380 28908 3392
rect 27764 3352 28908 3380
rect 27764 3340 27770 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 32398 3340 32404 3392
rect 32456 3380 32462 3392
rect 33042 3380 33048 3392
rect 32456 3352 33048 3380
rect 32456 3340 32462 3352
rect 33042 3340 33048 3352
rect 33100 3340 33106 3392
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 38105 3383 38163 3389
rect 38105 3349 38117 3383
rect 38151 3380 38163 3383
rect 38151 3352 57192 3380
rect 38151 3349 38163 3352
rect 38105 3343 38163 3349
rect 9950 3272 9956 3324
rect 10008 3312 10014 3324
rect 43438 3312 43444 3324
rect 10008 3284 43444 3312
rect 10008 3272 10014 3284
rect 43438 3272 43444 3284
rect 43496 3272 43502 3324
rect 46658 3272 46664 3324
rect 46716 3312 46722 3324
rect 57057 3315 57115 3321
rect 57057 3312 57069 3315
rect 46716 3284 57069 3312
rect 46716 3272 46722 3284
rect 57057 3281 57069 3284
rect 57103 3281 57115 3315
rect 57164 3312 57192 3352
rect 57238 3340 57244 3392
rect 57296 3380 57302 3392
rect 57882 3380 57888 3392
rect 57296 3352 57888 3380
rect 57296 3340 57302 3352
rect 57882 3340 57888 3352
rect 57940 3340 57946 3392
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 60642 3380 60648 3392
rect 59688 3352 60648 3380
rect 59688 3340 59694 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 60826 3340 60832 3392
rect 60884 3380 60890 3392
rect 62022 3380 62028 3392
rect 60884 3352 62028 3380
rect 60884 3340 60890 3352
rect 62022 3340 62028 3352
rect 62080 3340 62086 3392
rect 64322 3340 64328 3392
rect 64380 3380 64386 3392
rect 64782 3380 64788 3392
rect 64380 3352 64788 3380
rect 64380 3340 64386 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 66640 3380 66668 3420
rect 66714 3408 66720 3460
rect 66772 3448 66778 3460
rect 67542 3448 67548 3460
rect 66772 3420 67548 3448
rect 66772 3408 66778 3420
rect 67542 3408 67548 3420
rect 67600 3408 67606 3460
rect 67910 3408 67916 3460
rect 67968 3448 67974 3460
rect 68922 3448 68928 3460
rect 67968 3420 68928 3448
rect 67968 3408 67974 3420
rect 68922 3408 68928 3420
rect 68980 3408 68986 3460
rect 72602 3408 72608 3460
rect 72660 3448 72666 3460
rect 73062 3448 73068 3460
rect 72660 3420 73068 3448
rect 72660 3408 72666 3420
rect 73062 3408 73068 3420
rect 73120 3408 73126 3460
rect 73798 3408 73804 3460
rect 73856 3448 73862 3460
rect 74442 3448 74448 3460
rect 73856 3420 74448 3448
rect 73856 3408 73862 3420
rect 74442 3408 74448 3420
rect 74500 3408 74506 3460
rect 131758 3408 131764 3460
rect 131816 3448 131822 3460
rect 132402 3448 132408 3460
rect 131816 3420 132408 3448
rect 131816 3408 131822 3420
rect 132402 3408 132408 3420
rect 132460 3408 132466 3460
rect 158530 3408 158536 3460
rect 158588 3448 158594 3460
rect 160094 3448 160100 3460
rect 158588 3420 160100 3448
rect 158588 3408 158594 3420
rect 160094 3408 160100 3420
rect 160152 3408 160158 3460
rect 166902 3408 166908 3460
rect 166960 3448 166966 3460
rect 170766 3448 170772 3460
rect 166960 3420 170772 3448
rect 166960 3408 166966 3420
rect 170766 3408 170772 3420
rect 170824 3408 170830 3460
rect 171042 3408 171048 3460
rect 171100 3448 171106 3460
rect 176654 3448 176660 3460
rect 171100 3420 176660 3448
rect 171100 3408 171106 3420
rect 176654 3408 176660 3420
rect 176712 3408 176718 3460
rect 177758 3408 177764 3460
rect 177816 3448 177822 3460
rect 184934 3448 184940 3460
rect 177816 3420 184940 3448
rect 177816 3408 177822 3420
rect 184934 3408 184940 3420
rect 184992 3408 184998 3460
rect 186222 3408 186228 3460
rect 186280 3448 186286 3460
rect 197906 3448 197912 3460
rect 186280 3420 197912 3448
rect 186280 3408 186286 3420
rect 197906 3408 197912 3420
rect 197964 3408 197970 3460
rect 198550 3408 198556 3460
rect 198608 3448 198614 3460
rect 214466 3448 214472 3460
rect 198608 3420 214472 3448
rect 198608 3408 198614 3420
rect 214466 3408 214472 3420
rect 214524 3408 214530 3460
rect 215202 3408 215208 3460
rect 215260 3448 215266 3460
rect 237006 3448 237012 3460
rect 215260 3420 237012 3448
rect 215260 3408 215266 3420
rect 237006 3408 237012 3420
rect 237064 3408 237070 3460
rect 240042 3408 240048 3460
rect 240100 3448 240106 3460
rect 270034 3448 270040 3460
rect 240100 3420 270040 3448
rect 240100 3408 240106 3420
rect 270034 3408 270040 3420
rect 270092 3408 270098 3460
rect 270402 3408 270408 3460
rect 270460 3448 270466 3460
rect 307665 3451 307723 3457
rect 307665 3448 307677 3451
rect 270460 3420 307677 3448
rect 270460 3408 270466 3420
rect 307665 3417 307677 3420
rect 307711 3417 307723 3451
rect 307665 3411 307723 3417
rect 307754 3408 307760 3460
rect 307812 3448 307818 3460
rect 309042 3448 309048 3460
rect 307812 3420 309048 3448
rect 307812 3408 307818 3420
rect 309042 3408 309048 3420
rect 309100 3408 309106 3460
rect 314562 3408 314568 3460
rect 314620 3448 314626 3460
rect 372890 3448 372896 3460
rect 314620 3420 372896 3448
rect 314620 3408 314626 3420
rect 372890 3408 372896 3420
rect 372948 3408 372954 3460
rect 373902 3408 373908 3460
rect 373960 3448 373966 3460
rect 454494 3448 454500 3460
rect 373960 3420 454500 3448
rect 373960 3408 373966 3420
rect 454494 3408 454500 3420
rect 454552 3408 454558 3460
rect 463602 3408 463608 3460
rect 463660 3448 463666 3460
rect 578602 3448 578608 3460
rect 463660 3420 578608 3448
rect 463660 3408 463666 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 73430 3380 73436 3392
rect 66640 3352 73436 3380
rect 73430 3340 73436 3352
rect 73488 3340 73494 3392
rect 173802 3340 173808 3392
rect 173860 3380 173866 3392
rect 180242 3380 180248 3392
rect 173860 3352 180248 3380
rect 173860 3340 173866 3352
rect 180242 3340 180248 3352
rect 180300 3340 180306 3392
rect 184842 3340 184848 3392
rect 184900 3380 184906 3392
rect 194410 3380 194416 3392
rect 184900 3352 194416 3380
rect 184900 3340 184906 3352
rect 194410 3340 194416 3352
rect 194468 3340 194474 3392
rect 201402 3340 201408 3392
rect 201460 3380 201466 3392
rect 218054 3380 218060 3392
rect 201460 3352 218060 3380
rect 201460 3340 201466 3352
rect 218054 3340 218060 3352
rect 218112 3340 218118 3392
rect 219342 3340 219348 3392
rect 219400 3380 219406 3392
rect 241698 3380 241704 3392
rect 219400 3352 241704 3380
rect 219400 3340 219406 3352
rect 241698 3340 241704 3352
rect 241756 3340 241762 3392
rect 243998 3340 244004 3392
rect 244056 3380 244062 3392
rect 277118 3380 277124 3392
rect 244056 3352 277124 3380
rect 244056 3340 244062 3352
rect 277118 3340 277124 3352
rect 277176 3340 277182 3392
rect 293862 3340 293868 3392
rect 293920 3380 293926 3392
rect 344554 3380 344560 3392
rect 293920 3352 344560 3380
rect 293920 3340 293926 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 344922 3340 344928 3392
rect 344980 3380 344986 3392
rect 415486 3380 415492 3392
rect 344980 3352 415492 3380
rect 344980 3340 344986 3352
rect 415486 3340 415492 3352
rect 415544 3340 415550 3392
rect 438762 3340 438768 3392
rect 438820 3380 438826 3392
rect 543182 3380 543188 3392
rect 438820 3352 543188 3380
rect 438820 3340 438826 3352
rect 543182 3340 543188 3352
rect 543240 3340 543246 3392
rect 551278 3340 551284 3392
rect 551336 3380 551342 3392
rect 552658 3380 552664 3392
rect 551336 3352 552664 3380
rect 551336 3340 551342 3352
rect 552658 3340 552664 3352
rect 552716 3340 552722 3392
rect 558178 3340 558184 3392
rect 558236 3380 558242 3392
rect 559742 3380 559748 3392
rect 558236 3352 559748 3380
rect 558236 3340 558242 3352
rect 559742 3340 559748 3352
rect 559800 3340 559806 3392
rect 63586 3312 63592 3324
rect 57164 3284 63592 3312
rect 57057 3275 57115 3281
rect 63586 3272 63592 3284
rect 63644 3272 63650 3324
rect 138842 3272 138848 3324
rect 138900 3312 138906 3324
rect 139302 3312 139308 3324
rect 138900 3284 139308 3312
rect 138900 3272 138906 3284
rect 139302 3272 139308 3284
rect 139360 3272 139366 3324
rect 200022 3272 200028 3324
rect 200080 3312 200086 3324
rect 215662 3312 215668 3324
rect 200080 3284 215668 3312
rect 200080 3272 200086 3284
rect 215662 3272 215668 3284
rect 215720 3272 215726 3324
rect 220722 3272 220728 3324
rect 220780 3312 220786 3324
rect 244090 3312 244096 3324
rect 220780 3284 244096 3312
rect 220780 3272 220786 3284
rect 244090 3272 244096 3284
rect 244148 3272 244154 3324
rect 246942 3272 246948 3324
rect 247000 3312 247006 3324
rect 279510 3312 279516 3324
rect 247000 3284 279516 3312
rect 247000 3272 247006 3284
rect 279510 3272 279516 3284
rect 279568 3272 279574 3324
rect 288342 3272 288348 3324
rect 288400 3312 288406 3324
rect 337470 3312 337476 3324
rect 288400 3284 337476 3312
rect 288400 3272 288406 3284
rect 337470 3272 337476 3284
rect 337528 3272 337534 3324
rect 349154 3272 349160 3324
rect 349212 3312 349218 3324
rect 350442 3312 350448 3324
rect 349212 3284 350448 3312
rect 349212 3272 349218 3284
rect 350442 3272 350448 3284
rect 350500 3272 350506 3324
rect 350537 3315 350595 3321
rect 350537 3281 350549 3315
rect 350583 3312 350595 3315
rect 418982 3312 418988 3324
rect 350583 3284 418988 3312
rect 350583 3281 350595 3284
rect 350537 3275 350595 3281
rect 418982 3272 418988 3284
rect 419040 3272 419046 3324
rect 436002 3272 436008 3324
rect 436060 3312 436066 3324
rect 539594 3312 539600 3324
rect 436060 3284 539600 3312
rect 436060 3272 436066 3284
rect 539594 3272 539600 3284
rect 539652 3272 539658 3324
rect 21818 3204 21824 3256
rect 21876 3244 21882 3256
rect 31021 3247 31079 3253
rect 31021 3244 31033 3247
rect 21876 3216 31033 3244
rect 21876 3204 21882 3216
rect 31021 3213 31033 3216
rect 31067 3213 31079 3247
rect 31021 3207 31079 3213
rect 33594 3204 33600 3256
rect 33652 3244 33658 3256
rect 66346 3244 66352 3256
rect 33652 3216 66352 3244
rect 33652 3204 33658 3216
rect 66346 3204 66352 3216
rect 66404 3204 66410 3256
rect 172422 3204 172428 3256
rect 172480 3244 172486 3256
rect 179046 3244 179052 3256
rect 172480 3216 179052 3244
rect 172480 3204 172486 3216
rect 179046 3204 179052 3216
rect 179104 3204 179110 3256
rect 195882 3204 195888 3256
rect 195940 3244 195946 3256
rect 210970 3244 210976 3256
rect 195940 3216 210976 3244
rect 195940 3204 195946 3216
rect 210970 3204 210976 3216
rect 211028 3204 211034 3256
rect 216582 3204 216588 3256
rect 216640 3244 216646 3256
rect 238110 3244 238116 3256
rect 216640 3216 238116 3244
rect 216640 3204 216646 3216
rect 238110 3204 238116 3216
rect 238168 3204 238174 3256
rect 244182 3204 244188 3256
rect 244240 3244 244246 3256
rect 276014 3244 276020 3256
rect 244240 3216 276020 3244
rect 244240 3204 244246 3216
rect 276014 3204 276020 3216
rect 276072 3204 276078 3256
rect 285582 3204 285588 3256
rect 285640 3244 285646 3256
rect 333882 3244 333888 3256
rect 285640 3216 333888 3244
rect 285640 3204 285646 3216
rect 333882 3204 333888 3216
rect 333940 3204 333946 3256
rect 342070 3204 342076 3256
rect 342128 3244 342134 3256
rect 411898 3244 411904 3256
rect 342128 3216 411904 3244
rect 342128 3204 342134 3216
rect 411898 3204 411904 3216
rect 411956 3204 411962 3256
rect 433150 3204 433156 3256
rect 433208 3244 433214 3256
rect 536098 3244 536104 3256
rect 433208 3216 536104 3244
rect 433208 3204 433214 3216
rect 536098 3204 536104 3216
rect 536156 3204 536162 3256
rect 569218 3204 569224 3256
rect 569276 3244 569282 3256
rect 570322 3244 570328 3256
rect 569276 3216 570328 3244
rect 569276 3204 569282 3216
rect 570322 3204 570328 3216
rect 570380 3204 570386 3256
rect 30098 3136 30104 3188
rect 30156 3176 30162 3188
rect 38105 3179 38163 3185
rect 38105 3176 38117 3179
rect 30156 3148 38117 3176
rect 30156 3136 30162 3148
rect 38105 3145 38117 3148
rect 38151 3145 38163 3179
rect 69198 3176 69204 3188
rect 38105 3139 38163 3145
rect 38212 3148 69204 3176
rect 37182 3068 37188 3120
rect 37240 3108 37246 3120
rect 38212 3108 38240 3148
rect 69198 3136 69204 3148
rect 69256 3136 69262 3188
rect 165522 3136 165528 3188
rect 165580 3176 165586 3188
rect 168374 3176 168380 3188
rect 165580 3148 168380 3176
rect 165580 3136 165586 3148
rect 168374 3136 168380 3148
rect 168432 3136 168438 3188
rect 175090 3136 175096 3188
rect 175148 3176 175154 3188
rect 181438 3176 181444 3188
rect 175148 3148 181444 3176
rect 175148 3136 175154 3148
rect 181438 3136 181444 3148
rect 181496 3136 181502 3188
rect 197262 3136 197268 3188
rect 197320 3176 197326 3188
rect 212166 3176 212172 3188
rect 197320 3148 212172 3176
rect 197320 3136 197326 3148
rect 212166 3136 212172 3148
rect 212224 3136 212230 3188
rect 213822 3136 213828 3188
rect 213880 3176 213886 3188
rect 234614 3176 234620 3188
rect 213880 3148 234620 3176
rect 213880 3136 213886 3148
rect 234614 3136 234620 3148
rect 234672 3136 234678 3188
rect 237282 3136 237288 3188
rect 237340 3176 237346 3188
rect 266538 3176 266544 3188
rect 237340 3148 266544 3176
rect 237340 3136 237346 3148
rect 266538 3136 266544 3148
rect 266596 3136 266602 3188
rect 278682 3136 278688 3188
rect 278740 3176 278746 3188
rect 323302 3176 323308 3188
rect 278740 3148 323308 3176
rect 278740 3136 278746 3148
rect 323302 3136 323308 3148
rect 323360 3136 323366 3188
rect 324314 3136 324320 3188
rect 324372 3176 324378 3188
rect 325602 3176 325608 3188
rect 324372 3148 325608 3176
rect 324372 3136 324378 3148
rect 325602 3136 325608 3148
rect 325660 3136 325666 3188
rect 340782 3136 340788 3188
rect 340840 3176 340846 3188
rect 408402 3176 408408 3188
rect 340840 3148 408408 3176
rect 340840 3136 340846 3148
rect 408402 3136 408408 3148
rect 408460 3136 408466 3188
rect 427722 3136 427728 3188
rect 427780 3176 427786 3188
rect 529014 3176 529020 3188
rect 427780 3148 529020 3176
rect 427780 3136 427786 3148
rect 529014 3136 529020 3148
rect 529072 3136 529078 3188
rect 37240 3080 38240 3108
rect 37240 3068 37246 3080
rect 40678 3068 40684 3120
rect 40736 3108 40742 3120
rect 70486 3108 70492 3120
rect 40736 3080 70492 3108
rect 40736 3068 40742 3080
rect 70486 3068 70492 3080
rect 70544 3068 70550 3120
rect 193122 3068 193128 3120
rect 193180 3108 193186 3120
rect 206186 3108 206192 3120
rect 193180 3080 206192 3108
rect 193180 3068 193186 3080
rect 206186 3068 206192 3080
rect 206244 3068 206250 3120
rect 209682 3068 209688 3120
rect 209740 3108 209746 3120
rect 229830 3108 229836 3120
rect 209740 3080 229836 3108
rect 209740 3068 209746 3080
rect 229830 3068 229836 3080
rect 229888 3068 229894 3120
rect 235902 3068 235908 3120
rect 235960 3108 235966 3120
rect 265342 3108 265348 3120
rect 235960 3080 265348 3108
rect 235960 3068 235966 3080
rect 265342 3068 265348 3080
rect 265400 3068 265406 3120
rect 307665 3111 307723 3117
rect 307665 3077 307677 3111
rect 307711 3108 307723 3111
rect 312630 3108 312636 3120
rect 307711 3080 312636 3108
rect 307711 3077 307723 3080
rect 307665 3071 307723 3077
rect 312630 3068 312636 3080
rect 312688 3068 312694 3120
rect 338022 3068 338028 3120
rect 338080 3108 338086 3120
rect 404814 3108 404820 3120
rect 338080 3080 404820 3108
rect 338080 3068 338086 3080
rect 404814 3068 404820 3080
rect 404872 3068 404878 3120
rect 430482 3068 430488 3120
rect 430540 3108 430546 3120
rect 532510 3108 532516 3120
rect 430540 3080 532516 3108
rect 430540 3068 430546 3080
rect 532510 3068 532516 3080
rect 532568 3068 532574 3120
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 46198 3040 46204 3052
rect 19484 3012 46204 3040
rect 19484 3000 19490 3012
rect 46198 3000 46204 3012
rect 46256 3000 46262 3052
rect 47854 3000 47860 3052
rect 47912 3040 47918 3052
rect 53745 3043 53803 3049
rect 53745 3040 53757 3043
rect 47912 3012 53757 3040
rect 47912 3000 47918 3012
rect 53745 3009 53757 3012
rect 53791 3009 53803 3043
rect 53745 3003 53803 3009
rect 148318 3000 148324 3052
rect 148376 3040 148382 3052
rect 148962 3040 148968 3052
rect 148376 3012 148968 3040
rect 148376 3000 148382 3012
rect 148962 3000 148968 3012
rect 149020 3000 149026 3052
rect 162762 3000 162768 3052
rect 162820 3040 162826 3052
rect 164878 3040 164884 3052
rect 162820 3012 164884 3040
rect 162820 3000 162826 3012
rect 164878 3000 164884 3012
rect 164936 3000 164942 3052
rect 209590 3000 209596 3052
rect 209648 3040 209654 3052
rect 228726 3040 228732 3052
rect 209648 3012 228732 3040
rect 209648 3000 209654 3012
rect 228726 3000 228732 3012
rect 228784 3000 228790 3052
rect 238662 3000 238668 3052
rect 238720 3040 238726 3052
rect 268838 3040 268844 3052
rect 238720 3012 268844 3040
rect 238720 3000 238726 3012
rect 268838 3000 268844 3012
rect 268896 3000 268902 3052
rect 335262 3000 335268 3052
rect 335320 3040 335326 3052
rect 335320 3012 398788 3040
rect 335320 3000 335326 3012
rect 28902 2932 28908 2984
rect 28960 2972 28966 2984
rect 48866 2972 48872 2984
rect 28960 2944 48872 2972
rect 28960 2932 28966 2944
rect 48866 2932 48872 2944
rect 48924 2932 48930 2984
rect 141234 2932 141240 2984
rect 141292 2972 141298 2984
rect 142062 2972 142068 2984
rect 141292 2944 142068 2972
rect 141292 2932 141298 2944
rect 142062 2932 142068 2944
rect 142120 2932 142126 2984
rect 175182 2932 175188 2984
rect 175240 2972 175246 2984
rect 182542 2972 182548 2984
rect 175240 2944 182548 2972
rect 175240 2932 175246 2944
rect 182542 2932 182548 2944
rect 182600 2932 182606 2984
rect 208302 2932 208308 2984
rect 208360 2972 208366 2984
rect 227530 2972 227536 2984
rect 208360 2944 227536 2972
rect 208360 2932 208366 2944
rect 227530 2932 227536 2944
rect 227588 2932 227594 2984
rect 233142 2932 233148 2984
rect 233200 2972 233206 2984
rect 261754 2972 261760 2984
rect 233200 2944 261760 2972
rect 233200 2932 233206 2944
rect 261754 2932 261760 2944
rect 261812 2932 261818 2984
rect 332502 2932 332508 2984
rect 332560 2972 332566 2984
rect 397730 2972 397736 2984
rect 332560 2944 397736 2972
rect 332560 2932 332566 2944
rect 397730 2932 397736 2944
rect 397788 2932 397794 2984
rect 398760 2972 398788 3012
rect 398834 3000 398840 3052
rect 398892 3040 398898 3052
rect 400122 3040 400128 3052
rect 398892 3012 400128 3040
rect 398892 3000 398898 3012
rect 400122 3000 400128 3012
rect 400180 3000 400186 3052
rect 422110 3000 422116 3052
rect 422168 3040 422174 3052
rect 521838 3040 521844 3052
rect 422168 3012 521844 3040
rect 422168 3000 422174 3012
rect 521838 3000 521844 3012
rect 521896 3000 521902 3052
rect 560938 3000 560944 3052
rect 560996 3040 561002 3052
rect 563238 3040 563244 3052
rect 560996 3012 563244 3040
rect 560996 3000 561002 3012
rect 563238 3000 563244 3012
rect 563296 3000 563302 3052
rect 401318 2972 401324 2984
rect 398760 2944 401324 2972
rect 401318 2932 401324 2944
rect 401376 2932 401382 2984
rect 424778 2932 424784 2984
rect 424836 2972 424842 2984
rect 525426 2972 525432 2984
rect 424836 2944 525432 2972
rect 424836 2932 424842 2944
rect 525426 2932 525432 2944
rect 525484 2932 525490 2984
rect 35986 2864 35992 2916
rect 36044 2904 36050 2916
rect 55858 2904 55864 2916
rect 36044 2876 55864 2904
rect 36044 2864 36050 2876
rect 55858 2864 55864 2876
rect 55916 2864 55922 2916
rect 202782 2864 202788 2916
rect 202840 2904 202846 2916
rect 219250 2904 219256 2916
rect 202840 2876 219256 2904
rect 202840 2864 202846 2876
rect 219250 2864 219256 2876
rect 219308 2864 219314 2916
rect 229002 2864 229008 2916
rect 229060 2904 229066 2916
rect 255866 2904 255872 2916
rect 229060 2876 255872 2904
rect 229060 2864 229066 2876
rect 255866 2864 255872 2876
rect 255924 2864 255930 2916
rect 329742 2864 329748 2916
rect 329800 2904 329806 2916
rect 394234 2904 394240 2916
rect 329800 2876 394240 2904
rect 329800 2864 329806 2876
rect 394234 2864 394240 2876
rect 394292 2864 394298 2916
rect 420822 2864 420828 2916
rect 420880 2904 420886 2916
rect 518342 2904 518348 2916
rect 420880 2876 518348 2904
rect 420880 2864 420886 2876
rect 518342 2864 518348 2876
rect 518400 2864 518406 2916
rect 43070 2796 43076 2848
rect 43128 2836 43134 2848
rect 62758 2836 62764 2848
rect 43128 2808 62764 2836
rect 43128 2796 43134 2808
rect 62758 2796 62764 2808
rect 62816 2796 62822 2848
rect 198642 2796 198648 2848
rect 198700 2836 198706 2848
rect 213362 2836 213368 2848
rect 198700 2808 213368 2836
rect 198700 2796 198706 2808
rect 213362 2796 213368 2808
rect 213420 2796 213426 2848
rect 226242 2796 226248 2848
rect 226300 2836 226306 2848
rect 251174 2836 251180 2848
rect 226300 2808 251180 2836
rect 226300 2796 226306 2808
rect 251174 2796 251180 2808
rect 251232 2796 251238 2848
rect 321462 2796 321468 2848
rect 321520 2836 321526 2848
rect 383562 2836 383568 2848
rect 321520 2808 383568 2836
rect 321520 2796 321526 2808
rect 383562 2796 383568 2808
rect 383620 2796 383626 2848
rect 383654 2796 383660 2848
rect 383712 2836 383718 2848
rect 468662 2836 468668 2848
rect 383712 2808 468668 2836
rect 383712 2796 383718 2808
rect 468662 2796 468668 2808
rect 468720 2796 468726 2848
<< via1 >>
rect 238668 700952 238720 701004
rect 397460 700952 397512 701004
rect 241428 700884 241480 700936
rect 413652 700884 413704 700936
rect 89168 700816 89220 700868
rect 296720 700816 296772 700868
rect 72976 700748 73028 700800
rect 292580 700748 292632 700800
rect 227628 700680 227680 700732
rect 462320 700680 462372 700732
rect 230388 700612 230440 700664
rect 478512 700612 478564 700664
rect 40500 700544 40552 700596
rect 300860 700544 300912 700596
rect 24308 700476 24360 700528
rect 307760 700476 307812 700528
rect 8116 700408 8168 700460
rect 303620 700408 303672 700460
rect 215208 700340 215260 700392
rect 527180 700340 527232 700392
rect 219348 700272 219400 700324
rect 543464 700272 543516 700324
rect 137836 700204 137888 700256
rect 281540 700204 281592 700256
rect 154120 700136 154172 700188
rect 285680 700136 285732 700188
rect 252468 700068 252520 700120
rect 348792 700068 348844 700120
rect 249708 700000 249760 700052
rect 332508 700000 332560 700052
rect 202788 699932 202840 699984
rect 270500 699932 270552 699984
rect 218980 699864 219032 699916
rect 274640 699864 274692 699916
rect 264888 699796 264940 699848
rect 283840 699796 283892 699848
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 260748 699660 260800 699712
rect 267648 699660 267700 699712
rect 204168 696940 204220 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 311900 683204 311952 683256
rect 208308 683136 208360 683188
rect 580172 683136 580224 683188
rect 3424 670760 3476 670812
rect 318800 670760 318852 670812
rect 201408 670692 201460 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 314660 656888 314712 656940
rect 193128 643084 193180 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 322940 632068 322992 632120
rect 197268 630640 197320 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 329840 618264 329892 618316
rect 190368 616836 190420 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 325700 605820 325752 605872
rect 182088 590656 182140 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 333980 579640 334032 579692
rect 186228 576852 186280 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 340880 565836 340932 565888
rect 177948 563048 178000 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 338120 553392 338172 553444
rect 170956 536800 171008 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 345020 527144 345072 527196
rect 175188 524424 175240 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 351920 514768 351972 514820
rect 166908 510620 166960 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 349160 500964 349212 501016
rect 160008 484372 160060 484424
rect 580172 484372 580224 484424
rect 3424 474716 3476 474768
rect 356244 474716 356296 474768
rect 22836 472132 22888 472184
rect 386420 472132 386472 472184
rect 129648 472064 129700 472116
rect 512644 472064 512696 472116
rect 85120 471996 85172 472048
rect 511264 471996 511316 472048
rect 159548 471928 159600 471980
rect 160008 471928 160060 471980
rect 174452 471928 174504 471980
rect 175188 471928 175240 471980
rect 185676 471928 185728 471980
rect 186228 471928 186280 471980
rect 189356 471928 189408 471980
rect 190368 471928 190420 471980
rect 196808 471928 196860 471980
rect 197268 471928 197320 471980
rect 200580 471928 200632 471980
rect 201408 471928 201460 471980
rect 226616 471928 226668 471980
rect 227628 471928 227680 471980
rect 248972 471928 249024 471980
rect 249708 471928 249760 471980
rect 260104 471928 260156 471980
rect 260748 471928 260800 471980
rect 263876 471928 263928 471980
rect 264888 471928 264940 471980
rect 235908 471860 235960 471912
rect 266912 471860 266964 471912
rect 256424 471792 256476 471844
rect 299480 471792 299532 471844
rect 171048 471724 171100 471776
rect 278136 471724 278188 471776
rect 81348 471656 81400 471708
rect 106188 471588 106240 471640
rect 148416 471520 148468 471572
rect 223396 471520 223448 471572
rect 234068 471656 234120 471708
rect 234988 471520 235040 471572
rect 237840 471656 237892 471708
rect 238668 471656 238720 471708
rect 245292 471656 245344 471708
rect 364340 471656 364392 471708
rect 289268 471588 289320 471640
rect 429200 471520 429252 471572
rect 222936 471452 222988 471504
rect 494060 471452 494112 471504
rect 140688 471384 140740 471436
rect 467380 471384 467432 471436
rect 211712 471316 211764 471368
rect 558920 471316 558972 471368
rect 118608 471248 118660 471300
rect 467288 471248 467340 471300
rect 107476 471180 107528 471232
rect 467196 471180 467248 471232
rect 96252 471112 96304 471164
rect 467104 471112 467156 471164
rect 29736 471044 29788 471096
rect 408500 471044 408552 471096
rect 32404 470976 32456 471028
rect 419632 470976 419684 471028
rect 33784 470908 33836 470960
rect 430856 470908 430908 470960
rect 92388 470840 92440 470892
rect 497464 470840 497516 470892
rect 35164 470772 35216 470824
rect 441988 470772 442040 470824
rect 36544 470704 36596 470756
rect 453212 470704 453264 470756
rect 163320 470636 163372 470688
rect 580172 470636 580224 470688
rect 40684 470568 40736 470620
rect 464344 470568 464396 470620
rect 155868 470364 155920 470416
rect 468484 470364 468536 470416
rect 39396 470296 39448 470348
rect 389824 470296 389876 470348
rect 133512 470228 133564 470280
rect 486424 470228 486476 470280
rect 223396 470160 223448 470212
rect 580448 470160 580500 470212
rect 3608 470092 3660 470144
rect 367468 470092 367520 470144
rect 111156 470024 111208 470076
rect 483664 470024 483716 470076
rect 15844 469956 15896 470008
rect 393596 469956 393648 470008
rect 88800 469888 88852 469940
rect 479524 469888 479576 469940
rect 18604 469820 18656 469872
rect 412180 469820 412232 469872
rect 103244 469752 103296 469804
rect 500224 469752 500276 469804
rect 17224 469684 17276 469736
rect 415952 469684 416004 469736
rect 65984 469616 66036 469668
rect 472624 469616 472676 469668
rect 21364 469548 21416 469600
rect 434720 469548 434772 469600
rect 70216 469480 70268 469532
rect 493324 469480 493376 469532
rect 7564 469412 7616 469464
rect 438308 469412 438360 469464
rect 29644 469344 29696 469396
rect 461124 469344 461176 469396
rect 58992 469276 59044 469328
rect 490564 469276 490616 469328
rect 11704 469208 11756 469260
rect 456892 469208 456944 469260
rect 152096 469047 152148 469056
rect 152096 469013 152105 469047
rect 152105 469013 152139 469047
rect 152139 469013 152148 469047
rect 152096 469004 152148 469013
rect 234988 469004 235040 469056
rect 580264 469004 580316 469056
rect 15936 468936 15988 468988
rect 360200 468936 360252 468988
rect 144736 468868 144788 468920
rect 489184 468868 489236 468920
rect 17316 468800 17368 468852
rect 371562 468800 371614 468852
rect 122380 468732 122432 468784
rect 485044 468732 485096 468784
rect 4896 468664 4948 468716
rect 378692 468664 378744 468716
rect 7656 468596 7708 468648
rect 382372 468596 382424 468648
rect 100024 468528 100076 468580
rect 482284 468528 482336 468580
rect 14464 468460 14516 468512
rect 401048 468460 401100 468512
rect 114928 468392 114980 468444
rect 501604 468392 501656 468444
rect 77668 468324 77720 468376
rect 475384 468324 475436 468376
rect 25504 468256 25556 468308
rect 423588 468256 423640 468308
rect 3516 468188 3568 468240
rect 404728 468188 404780 468240
rect 39304 468120 39356 468172
rect 449440 468120 449492 468172
rect 55128 468052 55180 468104
rect 471244 468052 471296 468104
rect 4804 467984 4856 468036
rect 427084 467984 427136 468036
rect 22744 467916 22796 467968
rect 445760 467984 445812 468036
rect 580356 467848 580408 467900
rect 3424 463632 3476 463684
rect 13820 463632 13872 463684
rect 468484 458124 468536 458176
rect 580172 458124 580224 458176
rect 3332 449828 3384 449880
rect 15936 449828 15988 449880
rect 2964 411204 3016 411256
rect 40776 411204 40828 411256
rect 489184 405628 489236 405680
rect 579620 405628 579672 405680
rect 3240 398760 3292 398812
rect 17316 398760 17368 398812
rect 504364 379448 504416 379500
rect 580172 379448 580224 379500
rect 2780 371356 2832 371408
rect 4896 371356 4948 371408
rect 467380 365644 467432 365696
rect 580172 365644 580224 365696
rect 3332 358708 3384 358760
rect 22836 358708 22888 358760
rect 486424 353200 486476 353252
rect 580172 353200 580224 353252
rect 3148 346332 3200 346384
rect 7656 346332 7708 346384
rect 502984 325592 503036 325644
rect 579896 325592 579948 325644
rect 3516 320084 3568 320136
rect 39396 320084 39448 320136
rect 512644 313216 512696 313268
rect 580172 313216 580224 313268
rect 3516 306280 3568 306332
rect 35256 306280 35308 306332
rect 485044 299412 485096 299464
rect 579620 299412 579672 299464
rect 3056 293904 3108 293956
rect 15844 293904 15896 293956
rect 501604 273164 501656 273216
rect 579896 273164 579948 273216
rect 3516 267656 3568 267708
rect 14464 267656 14516 267708
rect 467288 259360 467340 259412
rect 579804 259360 579856 259412
rect 3148 255212 3200 255264
rect 29736 255212 29788 255264
rect 483664 245556 483716 245608
rect 580172 245556 580224 245608
rect 500224 233180 500276 233232
rect 580172 233180 580224 233232
rect 467196 219376 467248 219428
rect 579896 219376 579948 219428
rect 3332 215228 3384 215280
rect 18604 215228 18656 215280
rect 482284 206932 482336 206984
rect 580172 206932 580224 206984
rect 3424 202784 3476 202836
rect 32404 202784 32456 202836
rect 497464 193128 497516 193180
rect 580172 193128 580224 193180
rect 3424 188980 3476 189032
rect 17224 188980 17276 189032
rect 467104 179324 467156 179376
rect 579988 179324 580040 179376
rect 479524 166948 479576 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 25504 164160 25556 164212
rect 3424 150356 3476 150408
rect 33784 150356 33836 150408
rect 511264 139340 511316 139392
rect 580172 139340 580224 139392
rect 2780 137096 2832 137148
rect 4804 137096 4856 137148
rect 475384 126896 475436 126948
rect 580172 126896 580224 126948
rect 493324 113092 493376 113144
rect 579804 113092 579856 113144
rect 3424 111732 3476 111784
rect 21364 111732 21416 111784
rect 508504 100648 508556 100700
rect 580172 100648 580224 100700
rect 3424 97928 3476 97980
rect 35164 97928 35216 97980
rect 472624 86912 472676 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 7564 85484 7616 85536
rect 490564 73108 490616 73160
rect 580172 73108 580224 73160
rect 3424 71680 3476 71732
rect 22744 71680 22796 71732
rect 507124 60664 507176 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 36544 59304 36596 59356
rect 471244 46860 471296 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 39304 45500 39356 45552
rect 56600 41828 56652 41880
rect 57842 41828 57894 41880
rect 70492 41828 70544 41880
rect 71642 41828 71694 41880
rect 26148 39992 26200 40044
rect 60372 39992 60424 40044
rect 67548 39992 67600 40044
rect 90548 39992 90600 40044
rect 95056 39992 95108 40044
rect 111156 39992 111208 40044
rect 111616 39992 111668 40044
rect 122380 39992 122432 40044
rect 128268 39992 128320 40044
rect 134432 39992 134484 40044
rect 142068 39992 142120 40044
rect 144736 39992 144788 40044
rect 266268 39992 266320 40044
rect 297272 39992 297324 40044
rect 299204 39992 299256 40044
rect 301596 39992 301648 40044
rect 322204 39992 322256 40044
rect 327448 39992 327500 40044
rect 342904 39992 342956 40044
rect 393780 39992 393832 40044
rect 481640 39992 481692 40044
rect 28908 39924 28960 39976
rect 62120 39924 62172 39976
rect 64788 39924 64840 39976
rect 88800 39924 88852 39976
rect 89628 39924 89680 39976
rect 106924 39924 106976 39976
rect 108948 39924 109000 39976
rect 120632 39924 120684 39976
rect 140688 39924 140740 39976
rect 143908 39924 143960 39976
rect 255136 39924 255188 39976
rect 24768 39856 24820 39908
rect 59544 39856 59596 39908
rect 62028 39856 62080 39908
rect 86224 39856 86276 39908
rect 86868 39856 86920 39908
rect 104256 39856 104308 39908
rect 107568 39856 107620 39908
rect 119804 39856 119856 39908
rect 126888 39856 126940 39908
rect 133604 39856 133656 39908
rect 137928 39856 137980 39908
rect 142160 39856 142212 39908
rect 268016 39924 268068 39976
rect 304264 39924 304316 39976
rect 319720 39924 319772 39976
rect 343824 39924 343876 39976
rect 352564 39924 352616 39976
rect 391204 39924 391256 39976
rect 478880 39924 478932 39976
rect 269672 39856 269724 39908
rect 23388 39788 23440 39840
rect 58624 39788 58676 39840
rect 60648 39788 60700 39840
rect 85396 39788 85448 39840
rect 91008 39788 91060 39840
rect 107752 39788 107804 39840
rect 110328 39788 110380 39840
rect 121552 39788 121604 39840
rect 122748 39788 122800 39840
rect 131120 39788 131172 39840
rect 244740 39788 244792 39840
rect 262864 39788 262916 39840
rect 275744 39788 275796 39840
rect 318064 39856 318116 39908
rect 325700 39856 325752 39908
rect 359556 39856 359608 39908
rect 486424 39856 486476 39908
rect 281816 39788 281868 39840
rect 327724 39788 327776 39840
rect 336004 39788 336056 39840
rect 348976 39788 349028 39840
rect 363512 39788 363564 39840
rect 369676 39788 369728 39840
rect 381544 39788 381596 39840
rect 398932 39788 398984 39840
rect 489920 39788 489972 39840
rect 16488 39720 16540 39772
rect 53472 39720 53524 39772
rect 63408 39720 63460 39772
rect 87972 39720 88024 39772
rect 88248 39720 88300 39772
rect 106004 39720 106056 39772
rect 111708 39720 111760 39772
rect 123208 39720 123260 39772
rect 125508 39720 125560 39772
rect 132684 39720 132736 39772
rect 257712 39720 257764 39772
rect 276572 39720 276624 39772
rect 280068 39720 280120 39772
rect 325700 39720 325752 39772
rect 326620 39720 326672 39772
rect 359464 39720 359516 39772
rect 361856 39720 361908 39772
rect 377312 39720 377364 39772
rect 402336 39720 402388 39772
rect 493324 39720 493376 39772
rect 19248 39652 19300 39704
rect 55220 39652 55272 39704
rect 57888 39652 57940 39704
rect 83648 39652 83700 39704
rect 85488 39652 85540 39704
rect 103520 39652 103572 39704
rect 104808 39652 104860 39704
rect 118056 39652 118108 39704
rect 119988 39652 120040 39704
rect 128452 39652 128504 39704
rect 242164 39652 242216 39704
rect 251824 39652 251876 39704
rect 252560 39652 252612 39704
rect 273904 39652 273956 39704
rect 283564 39652 283616 39704
rect 331220 39652 331272 39704
rect 333520 39652 333572 39704
rect 349712 39652 349764 39704
rect 351552 39652 351604 39704
rect 396724 39652 396776 39704
rect 404084 39652 404136 39704
rect 496820 39652 496872 39704
rect 15108 39584 15160 39636
rect 52644 39584 52696 39636
rect 53748 39584 53800 39636
rect 81072 39584 81124 39636
rect 84108 39584 84160 39636
rect 102600 39584 102652 39636
rect 103336 39584 103388 39636
rect 116400 39584 116452 39636
rect 118608 39584 118660 39636
rect 127532 39584 127584 39636
rect 129648 39584 129700 39636
rect 136180 39584 136232 39636
rect 247316 39584 247368 39636
rect 248972 39584 249024 39636
rect 262772 39584 262824 39636
rect 287704 39584 287756 39636
rect 289544 39584 289596 39636
rect 338764 39584 338816 39636
rect 346400 39584 346452 39636
rect 395344 39584 395396 39636
rect 397184 39584 397236 39636
rect 13728 39516 13780 39568
rect 51724 39516 51776 39568
rect 56508 39516 56560 39568
rect 82820 39516 82872 39568
rect 86776 39516 86828 39568
rect 105176 39516 105228 39568
rect 106188 39516 106240 39568
rect 118976 39516 119028 39568
rect 121368 39516 121420 39568
rect 130108 39516 130160 39568
rect 132408 39516 132460 39568
rect 138020 39516 138072 39568
rect 224132 39516 224184 39568
rect 244924 39516 244976 39568
rect 256792 39516 256844 39568
rect 293960 39516 294012 39568
rect 307668 39516 307720 39568
rect 356612 39516 356664 39568
rect 364524 39516 364576 39568
rect 413284 39516 413336 39568
rect 6828 39448 6880 39500
rect 46572 39448 46624 39500
rect 53656 39448 53708 39500
rect 80152 39448 80204 39500
rect 81348 39448 81400 39500
rect 100852 39448 100904 39500
rect 103428 39448 103480 39500
rect 117320 39448 117372 39500
rect 119896 39448 119948 39500
rect 129280 39448 129332 39500
rect 131028 39448 131080 39500
rect 137008 39448 137060 39500
rect 218980 39448 219032 39500
rect 224224 39448 224276 39500
rect 237012 39448 237064 39500
rect 267096 39448 267148 39500
rect 273168 39448 273220 39500
rect 282184 39448 282236 39500
rect 293868 39448 293920 39500
rect 345020 39448 345072 39500
rect 359280 39448 359332 39500
rect 411904 39448 411956 39500
rect 9588 39380 9640 39432
rect 48320 39380 48372 39432
rect 49608 39380 49660 39432
rect 77576 39380 77628 39432
rect 78496 39380 78548 39432
rect 98276 39380 98328 39432
rect 99288 39380 99340 39432
rect 113732 39380 113784 39432
rect 115848 39380 115900 39432
rect 125876 39380 125928 39432
rect 229284 39380 229336 39432
rect 255872 39380 255924 39432
rect 267188 39380 267240 39432
rect 307760 39380 307812 39432
rect 315396 39380 315448 39432
rect 370412 39380 370464 39432
rect 379980 39380 380032 39432
rect 388444 39380 388496 39432
rect 409236 39380 409288 39432
rect 503720 39584 503772 39636
rect 414388 39516 414440 39568
rect 510620 39516 510672 39568
rect 512644 39448 512696 39500
rect 4068 39312 4120 39364
rect 44916 39312 44968 39364
rect 45468 39312 45520 39364
rect 75000 39312 75052 39364
rect 75828 39312 75880 39364
rect 96620 39312 96672 39364
rect 97908 39312 97960 39364
rect 112904 39312 112956 39364
rect 113088 39312 113140 39364
rect 124220 39312 124272 39364
rect 128176 39312 128228 39364
rect 135260 39312 135312 39364
rect 216312 39312 216364 39364
rect 238024 39312 238076 39364
rect 246488 39312 246540 39364
rect 280252 39312 280304 39364
rect 282644 39312 282696 39364
rect 329932 39312 329984 39364
rect 31668 39244 31720 39296
rect 64696 39244 64748 39296
rect 70308 39244 70360 39296
rect 93124 39244 93176 39296
rect 95148 39244 95200 39296
rect 110420 39244 110472 39296
rect 117228 39244 117280 39296
rect 126704 39244 126756 39296
rect 258540 39244 258592 39296
rect 268384 39244 268436 39296
rect 289084 39244 289136 39296
rect 294696 39244 294748 39296
rect 307024 39244 307076 39296
rect 311992 39244 312044 39296
rect 324964 39244 325016 39296
rect 330852 39244 330904 39296
rect 393964 39312 394016 39364
rect 416136 39312 416188 39364
rect 423864 39312 423916 39364
rect 522304 39380 522356 39432
rect 434260 39312 434312 39364
rect 437296 39312 437348 39364
rect 441988 39312 442040 39364
rect 444196 39312 444248 39364
rect 462688 39312 462740 39364
rect 574744 39312 574796 39364
rect 387708 39244 387760 39296
rect 473360 39244 473412 39296
rect 33048 39176 33100 39228
rect 65524 39176 65576 39228
rect 71688 39176 71740 39228
rect 93952 39176 94004 39228
rect 96528 39176 96580 39228
rect 112076 39176 112128 39228
rect 114468 39176 114520 39228
rect 124956 39176 125008 39228
rect 405004 39176 405056 39228
rect 489184 39176 489236 39228
rect 38568 39108 38620 39160
rect 69848 39108 69900 39160
rect 74448 39108 74500 39160
rect 95700 39108 95752 39160
rect 100668 39108 100720 39160
rect 114652 39108 114704 39160
rect 392032 39108 392084 39160
rect 475384 39108 475436 39160
rect 35808 39040 35860 39092
rect 67272 39040 67324 39092
rect 68928 39040 68980 39092
rect 91100 39040 91152 39092
rect 92388 39040 92440 39092
rect 108580 39040 108632 39092
rect 136548 39040 136600 39092
rect 141332 39040 141384 39092
rect 239588 39040 239640 39092
rect 242164 39040 242216 39092
rect 410156 39040 410208 39092
rect 467104 39040 467156 39092
rect 39948 38972 40000 39024
rect 70676 38972 70728 39024
rect 73068 38972 73120 39024
rect 94872 38972 94924 39024
rect 102048 38972 102100 39024
rect 115480 38972 115532 39024
rect 139308 38972 139360 39024
rect 143080 38972 143132 39024
rect 143448 38972 143500 39024
rect 145656 38972 145708 39024
rect 146208 38972 146260 39024
rect 148232 38972 148284 39024
rect 148968 38972 149020 39024
rect 149980 38972 150032 39024
rect 151820 38972 151872 39024
rect 152556 38972 152608 39024
rect 157800 38972 157852 39024
rect 158536 38972 158588 39024
rect 159548 38972 159600 39024
rect 160008 38972 160060 39024
rect 162124 38972 162176 39024
rect 162768 38972 162820 39024
rect 162952 38972 163004 39024
rect 165712 38972 165764 39024
rect 166356 38972 166408 39024
rect 166908 38972 166960 39024
rect 167276 38972 167328 39024
rect 168288 38972 168340 39024
rect 169024 38972 169076 39024
rect 169668 38972 169720 39024
rect 169852 38972 169904 39024
rect 170956 38972 171008 39024
rect 171600 38972 171652 39024
rect 172336 38972 172388 39024
rect 173256 38972 173308 39024
rect 173808 38972 173860 39024
rect 175832 38972 175884 39024
rect 176568 38972 176620 39024
rect 178500 38972 178552 39024
rect 179328 38972 179380 39024
rect 180156 38972 180208 39024
rect 180708 38972 180760 39024
rect 181076 38972 181128 39024
rect 182088 38972 182140 39024
rect 182732 38972 182784 39024
rect 183468 38972 183520 39024
rect 183652 38972 183704 39024
rect 184848 38972 184900 39024
rect 185308 38972 185360 39024
rect 186136 38972 186188 39024
rect 187056 38972 187108 39024
rect 187608 38972 187660 39024
rect 187976 38972 188028 39024
rect 188896 38972 188948 39024
rect 189632 38972 189684 39024
rect 190368 38972 190420 39024
rect 190552 38972 190604 39024
rect 191656 38972 191708 39024
rect 192208 38972 192260 39024
rect 193128 38972 193180 39024
rect 193956 38972 194008 39024
rect 194508 38972 194560 39024
rect 194784 38972 194836 39024
rect 195796 38972 195848 39024
rect 196532 38972 196584 39024
rect 197268 38972 197320 39024
rect 197360 38972 197412 39024
rect 198648 38972 198700 39024
rect 199108 38972 199160 39024
rect 200028 38972 200080 39024
rect 200856 38972 200908 39024
rect 201408 38972 201460 39024
rect 201684 38972 201736 39024
rect 202788 38972 202840 39024
rect 203432 38972 203484 39024
rect 204168 38972 204220 39024
rect 206008 38972 206060 39024
rect 206836 38972 206888 39024
rect 207756 38972 207808 39024
rect 208308 38972 208360 39024
rect 208584 38972 208636 39024
rect 209596 38972 209648 39024
rect 210332 38972 210384 39024
rect 211068 38972 211120 39024
rect 211160 38972 211212 39024
rect 212356 38972 212408 39024
rect 212908 38972 212960 39024
rect 213828 38972 213880 39024
rect 214656 38972 214708 39024
rect 215208 38972 215260 39024
rect 215484 38972 215536 39024
rect 216588 38972 216640 39024
rect 217232 38972 217284 39024
rect 217968 38972 218020 39024
rect 218060 38972 218112 39024
rect 219348 38972 219400 39024
rect 219808 38972 219860 39024
rect 220728 38972 220780 39024
rect 224960 38972 225012 39024
rect 226248 38972 226300 39024
rect 226708 38972 226760 39024
rect 227536 38972 227588 39024
rect 228364 38972 228416 39024
rect 229008 38972 229060 39024
rect 231032 38972 231084 39024
rect 231768 38972 231820 39024
rect 232688 38972 232740 39024
rect 233148 38972 233200 39024
rect 235264 38972 235316 39024
rect 235908 38972 235960 39024
rect 236184 38972 236236 39024
rect 237288 38972 237340 39024
rect 237840 38972 237892 39024
rect 238668 38972 238720 39024
rect 238760 38972 238812 39024
rect 240048 38972 240100 39024
rect 240508 38972 240560 39024
rect 241428 38972 241480 39024
rect 243084 38972 243136 39024
rect 244188 38972 244240 39024
rect 245660 38972 245712 39024
rect 246948 38972 247000 39024
rect 249064 38972 249116 39024
rect 249708 38972 249760 39024
rect 249984 38972 250036 39024
rect 250996 38972 251048 39024
rect 251640 38972 251692 39024
rect 252468 38972 252520 39024
rect 253388 38972 253440 39024
rect 253848 38972 253900 39024
rect 254216 38972 254268 39024
rect 255228 38972 255280 39024
rect 255964 38972 256016 39024
rect 256608 38972 256660 39024
rect 260288 38972 260340 39024
rect 260748 38972 260800 39024
rect 261116 38972 261168 39024
rect 262956 38972 263008 39024
rect 263692 38972 263744 39024
rect 264796 38972 264848 39024
rect 265440 38972 265492 39024
rect 267004 38972 267056 39024
rect 269764 38972 269816 39024
rect 270408 38972 270460 39024
rect 270592 38972 270644 39024
rect 271788 38972 271840 39024
rect 272340 38972 272392 39024
rect 273168 38972 273220 39024
rect 274088 38972 274140 39024
rect 274548 38972 274600 39024
rect 274916 38972 274968 39024
rect 275928 38972 275980 39024
rect 276664 38972 276716 39024
rect 277308 38972 277360 39024
rect 277492 38972 277544 39024
rect 278688 38972 278740 39024
rect 279240 38972 279292 39024
rect 280804 38972 280856 39024
rect 280988 38972 281040 39024
rect 281448 38972 281500 39024
rect 286140 38972 286192 39024
rect 286968 38972 287020 39024
rect 288716 38972 288768 39024
rect 289728 38972 289780 39024
rect 290372 38972 290424 39024
rect 291108 38972 291160 39024
rect 291292 38972 291344 39024
rect 292488 38972 292540 39024
rect 293040 38972 293092 39024
rect 293868 38972 293920 39024
rect 295616 38972 295668 39024
rect 296628 38972 296680 39024
rect 298192 38972 298244 39024
rect 299388 38972 299440 39024
rect 299848 38972 299900 39024
rect 300676 38972 300728 39024
rect 302516 38972 302568 39024
rect 303436 38972 303488 39024
rect 305092 38972 305144 39024
rect 306196 38972 306248 39024
rect 306748 38972 306800 39024
rect 307668 38972 307720 39024
rect 309324 38972 309376 39024
rect 310428 38972 310480 39024
rect 311072 38972 311124 39024
rect 311808 38972 311860 39024
rect 313648 38972 313700 39024
rect 314568 38972 314620 39024
rect 316224 38972 316276 39024
rect 317328 38972 317380 39024
rect 317972 38972 318024 39024
rect 318708 38972 318760 39024
rect 318800 38972 318852 39024
rect 320088 38972 320140 39024
rect 320548 38972 320600 39024
rect 321376 38972 321428 39024
rect 323124 38972 323176 39024
rect 324136 38972 324188 39024
rect 324872 38972 324924 39024
rect 325608 38972 325660 39024
rect 329196 38972 329248 39024
rect 329748 38972 329800 39024
rect 330024 38972 330076 39024
rect 331128 38972 331180 39024
rect 331772 38972 331824 39024
rect 332508 38972 332560 39024
rect 332600 38972 332652 39024
rect 333888 38972 333940 39024
rect 334348 38972 334400 39024
rect 335268 38972 335320 39024
rect 336096 38972 336148 39024
rect 336648 38972 336700 39024
rect 336924 38972 336976 39024
rect 338028 38972 338080 39024
rect 338672 38972 338724 39024
rect 339408 38972 339460 39024
rect 339500 38972 339552 39024
rect 340788 38972 340840 39024
rect 341248 38972 341300 39024
rect 342076 38972 342128 39024
rect 342996 38972 343048 39024
rect 343548 38972 343600 39024
rect 345572 38972 345624 39024
rect 346308 38972 346360 39024
rect 347228 38972 347280 39024
rect 347688 38972 347740 39024
rect 348148 38972 348200 39024
rect 349068 38972 349120 39024
rect 349804 38972 349856 39024
rect 350448 38972 350500 39024
rect 350724 38972 350776 39024
rect 351828 38972 351880 39024
rect 352380 38972 352432 39024
rect 353208 38972 353260 39024
rect 353300 38972 353352 39024
rect 354588 38972 354640 39024
rect 355048 38972 355100 39024
rect 355968 38972 356020 39024
rect 356704 38972 356756 39024
rect 357348 38972 357400 39024
rect 357624 38972 357676 39024
rect 358728 38972 358780 39024
rect 360200 38972 360252 39024
rect 361488 38972 361540 39024
rect 363604 38972 363656 39024
rect 364248 38972 364300 39024
rect 366180 38972 366232 39024
rect 367008 38972 367060 39024
rect 367928 38972 367980 39024
rect 368388 38972 368440 39024
rect 368756 38972 368808 39024
rect 369768 38972 369820 39024
rect 370504 38972 370556 39024
rect 371148 38972 371200 39024
rect 373080 38972 373132 39024
rect 373908 38972 373960 39024
rect 374000 38972 374052 39024
rect 375288 38972 375340 39024
rect 375656 38972 375708 39024
rect 376668 38972 376720 39024
rect 377404 38972 377456 39024
rect 378048 38972 378100 39024
rect 382556 38972 382608 39024
rect 383476 38972 383528 39024
rect 384304 38972 384356 39024
rect 384948 38972 385000 39024
rect 388628 38972 388680 39024
rect 389088 38972 389140 39024
rect 389456 38972 389508 39024
rect 390468 38972 390520 39024
rect 395528 38972 395580 39024
rect 395988 38972 396040 39024
rect 396356 38972 396408 39024
rect 397368 38972 397420 39024
rect 398104 38972 398156 39024
rect 398748 38972 398800 39024
rect 400680 38972 400732 39024
rect 401508 38972 401560 39024
rect 403256 38972 403308 39024
rect 404268 38972 404320 39024
rect 405832 38972 405884 39024
rect 407028 38972 407080 39024
rect 417056 38972 417108 39024
rect 417976 38972 418028 39024
rect 418712 38972 418764 39024
rect 419448 38972 419500 39024
rect 419632 38972 419684 39024
rect 420828 38972 420880 39024
rect 423036 38972 423088 39024
rect 423588 38972 423640 39024
rect 425612 38972 425664 39024
rect 426348 38972 426400 39024
rect 428188 38972 428240 39024
rect 429108 38972 429160 39024
rect 429936 38972 429988 39024
rect 430488 38972 430540 39024
rect 430764 38972 430816 39024
rect 431868 38972 431920 39024
rect 432512 38972 432564 39024
rect 433248 38972 433300 39024
rect 433340 38972 433392 39024
rect 434628 38972 434680 39024
rect 435088 38972 435140 39024
rect 436008 38972 436060 39024
rect 436836 38972 436888 39024
rect 437388 38972 437440 39024
rect 437664 38972 437716 39024
rect 438768 38972 438820 39024
rect 440240 38972 440292 39024
rect 441528 38972 441580 39024
rect 443736 38972 443788 39024
rect 444288 38972 444340 39024
rect 446312 38972 446364 39024
rect 447048 38972 447100 39024
rect 448888 38972 448940 39024
rect 449808 38972 449860 39024
rect 450636 38972 450688 39024
rect 451188 38972 451240 39024
rect 451464 38972 451516 39024
rect 452476 38972 452528 39024
rect 453212 38972 453264 39024
rect 453948 38972 454000 39024
rect 454040 38972 454092 39024
rect 455328 38972 455380 39024
rect 455788 38972 455840 39024
rect 456708 38972 456760 39024
rect 457536 38972 457588 39024
rect 458088 38972 458140 39024
rect 458364 38972 458416 39024
rect 459468 38972 459520 39024
rect 460940 38972 460992 39024
rect 462228 38972 462280 39024
rect 465264 38972 465316 39024
rect 466276 38972 466328 39024
rect 42708 38904 42760 38956
rect 72424 38904 72476 38956
rect 77208 38904 77260 38956
rect 97448 38904 97500 38956
rect 137284 38904 137336 38956
rect 140504 38904 140556 38956
rect 144828 38904 144880 38956
rect 146484 38904 146536 38956
rect 147588 38904 147640 38956
rect 149060 38904 149112 38956
rect 154580 38904 154632 38956
rect 155132 38904 155184 38956
rect 160376 38904 160428 38956
rect 161388 38904 161440 38956
rect 176752 38904 176804 38956
rect 177856 38904 177908 38956
rect 222384 38904 222436 38956
rect 223488 38904 223540 38956
rect 231860 38904 231912 38956
rect 233056 38904 233108 38956
rect 284392 38904 284444 38956
rect 285496 38904 285548 38956
rect 308496 38904 308548 38956
rect 309048 38904 309100 38956
rect 322296 38904 322348 38956
rect 322848 38904 322900 38956
rect 367100 38904 367152 38956
rect 368296 38904 368348 38956
rect 371332 38904 371384 38956
rect 372528 38904 372580 38956
rect 378232 38904 378284 38956
rect 379428 38904 379480 38956
rect 426532 38904 426584 38956
rect 429844 38904 429896 38956
rect 464344 38904 464396 38956
rect 464988 38904 465040 38956
rect 43444 38836 43496 38888
rect 49148 38836 49200 38888
rect 50988 38836 51040 38888
rect 78404 38836 78456 38888
rect 79968 38836 80020 38888
rect 100024 38836 100076 38888
rect 133788 38836 133840 38888
rect 138756 38836 138808 38888
rect 304172 38836 304224 38888
rect 304908 38836 304960 38888
rect 381728 38836 381780 38888
rect 382188 38836 382240 38888
rect 48964 38768 49016 38820
rect 62948 38768 63000 38820
rect 64144 38768 64196 38820
rect 75920 38768 75972 38820
rect 78588 38768 78640 38820
rect 99104 38768 99156 38820
rect 135168 38768 135220 38820
rect 139584 38768 139636 38820
rect 164700 38768 164752 38820
rect 165528 38768 165580 38820
rect 168104 38768 168156 38820
rect 169024 38768 169076 38820
rect 174176 38768 174228 38820
rect 175096 38768 175148 38820
rect 204260 38768 204312 38820
rect 205456 38768 205508 38820
rect 221556 38768 221608 38820
rect 228364 38768 228416 38820
rect 233608 38768 233660 38820
rect 234528 38768 234580 38820
rect 287796 38768 287848 38820
rect 288348 38768 288400 38820
rect 386880 38768 386932 38820
rect 387708 38768 387760 38820
rect 55864 38700 55916 38752
rect 68100 38700 68152 38752
rect 82728 38700 82780 38752
rect 101680 38700 101732 38752
rect 144736 38700 144788 38752
rect 147404 38700 147456 38752
rect 439412 38700 439464 38752
rect 440148 38700 440200 38752
rect 46204 38632 46256 38684
rect 56048 38632 56100 38684
rect 62764 38632 62816 38684
rect 73252 38632 73304 38684
rect 93768 38632 93820 38684
rect 109500 38632 109552 38684
rect 124128 38632 124180 38684
rect 131856 38632 131908 38684
rect 385132 38360 385184 38412
rect 470600 38360 470652 38412
rect 407580 38292 407632 38344
rect 500960 38292 501012 38344
rect 412732 38224 412784 38276
rect 507860 38224 507912 38276
rect 421288 38156 421340 38208
rect 520280 38156 520332 38208
rect 437296 38088 437348 38140
rect 538220 38088 538272 38140
rect 444196 38020 444248 38072
rect 547880 38020 547932 38072
rect 444564 37952 444616 38004
rect 551284 37952 551336 38004
rect 299204 37884 299256 37936
rect 349160 37884 349212 37936
rect 349712 37884 349764 37936
rect 398840 37884 398892 37936
rect 452292 37884 452344 37936
rect 560944 37884 560996 37936
rect 406660 36864 406712 36916
rect 499580 36864 499632 36916
rect 411812 36796 411864 36848
rect 506480 36796 506532 36848
rect 447140 36728 447192 36780
rect 556252 36728 556304 36780
rect 449716 36660 449768 36712
rect 558184 36660 558236 36712
rect 454868 36592 454920 36644
rect 565820 36592 565872 36644
rect 460112 36524 460164 36576
rect 572720 36524 572772 36576
rect 397368 35232 397420 35284
rect 485780 35232 485832 35284
rect 417976 35164 418028 35216
rect 514760 35164 514812 35216
rect 378048 33736 378100 33788
rect 459560 33736 459612 33788
rect 2872 33056 2924 33108
rect 11704 33056 11756 33108
rect 383476 31016 383528 31068
rect 466460 31016 466512 31068
rect 339408 29588 339460 29640
rect 407212 29588 407264 29640
rect 375196 28228 375248 28280
rect 456892 28228 456944 28280
rect 372436 26868 372488 26920
rect 452660 26868 452712 26920
rect 357348 25508 357400 25560
rect 432052 25508 432104 25560
rect 342076 24080 342128 24132
rect 409880 24080 409932 24132
rect 328368 22720 328420 22772
rect 391940 22720 391992 22772
rect 401416 22720 401468 22772
rect 492680 22720 492732 22772
rect 280804 21360 280856 21412
rect 324320 21360 324372 21412
rect 325608 21360 325660 21412
rect 387800 21360 387852 21412
rect 388444 21360 388496 21412
rect 463700 21360 463752 21412
rect 3424 20612 3476 20664
rect 40684 20612 40736 20664
rect 336004 18572 336056 18624
rect 380900 18572 380952 18624
rect 381544 18572 381596 18624
rect 448520 18572 448572 18624
rect 286876 17280 286928 17332
rect 335360 17280 335412 17332
rect 317236 17212 317288 17264
rect 376760 17212 376812 17264
rect 377404 17212 377456 17264
rect 438860 17212 438912 17264
rect 289728 15920 289780 15972
rect 338672 15920 338724 15972
rect 336648 15852 336700 15904
rect 403624 15852 403676 15904
rect 307668 14424 307720 14476
rect 363512 14424 363564 14476
rect 363604 14424 363656 14476
rect 420920 14424 420972 14476
rect 299296 13064 299348 13116
rect 352564 13064 352616 13116
rect 414296 13064 414348 13116
rect 352840 12996 352892 13048
rect 304908 11704 304960 11756
rect 359280 11704 359332 11756
rect 368296 11704 368348 11756
rect 445760 11704 445812 11756
rect 233056 10276 233108 10328
rect 260656 10276 260708 10328
rect 278596 10276 278648 10328
rect 324412 10276 324464 10328
rect 324964 10276 325016 10328
rect 370136 10276 370188 10328
rect 458088 10276 458140 10328
rect 569224 10276 569276 10328
rect 264796 8984 264848 9036
rect 304356 8984 304408 9036
rect 390376 8984 390428 9036
rect 478144 8984 478196 9036
rect 296536 8916 296588 8968
rect 349252 8916 349304 8968
rect 359556 8916 359608 8968
rect 389456 8916 389508 8968
rect 411168 8916 411220 8968
rect 506480 8916 506532 8968
rect 338764 8236 338816 8288
rect 339868 8236 339920 8288
rect 411904 8236 411956 8288
rect 435548 8236 435600 8288
rect 441344 8236 441396 8288
rect 441528 8236 441580 8288
rect 413284 8168 413336 8220
rect 442632 8168 442684 8220
rect 394608 8100 394660 8152
rect 484032 8100 484084 8152
rect 400128 8032 400180 8084
rect 491116 8032 491168 8084
rect 413836 7964 413888 8016
rect 510068 7964 510120 8016
rect 322204 7896 322256 7948
rect 356336 7896 356388 7948
rect 419448 7896 419500 7948
rect 517152 7896 517204 7948
rect 310336 7828 310388 7880
rect 368204 7828 368256 7880
rect 429844 7828 429896 7880
rect 527824 7828 527876 7880
rect 318708 7760 318760 7812
rect 378876 7760 378928 7812
rect 431776 7760 431828 7812
rect 534908 7760 534960 7812
rect 321376 7692 321428 7744
rect 382372 7692 382424 7744
rect 395344 7692 395396 7744
rect 417884 7692 417936 7744
rect 429016 7692 429068 7744
rect 531320 7692 531372 7744
rect 249064 7624 249116 7676
rect 281908 7624 281960 7676
rect 282184 7624 282236 7676
rect 317236 7624 317288 7676
rect 324136 7624 324188 7676
rect 385960 7624 386012 7676
rect 396724 7624 396776 7676
rect 424876 7624 424928 7676
rect 437388 7624 437440 7676
rect 541992 7624 542044 7676
rect 228364 7556 228416 7608
rect 246396 7556 246448 7608
rect 277308 7556 277360 7608
rect 322112 7556 322164 7608
rect 354496 7556 354548 7608
rect 428464 7556 428516 7608
rect 440148 7556 440200 7608
rect 545488 7556 545540 7608
rect 370504 6876 370556 6928
rect 375288 6876 375340 6928
rect 3424 6808 3476 6860
rect 29644 6808 29696 6860
rect 379336 6808 379388 6860
rect 462780 6808 462832 6860
rect 467196 6808 467248 6860
rect 505376 6808 505428 6860
rect 384948 6740 385000 6792
rect 469864 6740 469916 6792
rect 390468 6672 390520 6724
rect 476948 6672 477000 6724
rect 292396 6604 292448 6656
rect 343364 6604 343416 6656
rect 356704 6604 356756 6656
rect 364616 6604 364668 6656
rect 387708 6604 387760 6656
rect 473452 6604 473504 6656
rect 300676 6536 300728 6588
rect 354036 6536 354088 6588
rect 359372 6536 359424 6588
rect 390652 6536 390704 6588
rect 395988 6536 396040 6588
rect 485228 6536 485280 6588
rect 306196 6468 306248 6520
rect 361120 6468 361172 6520
rect 393228 6468 393280 6520
rect 481732 6468 481784 6520
rect 310428 6400 310480 6452
rect 366916 6400 366968 6452
rect 401508 6400 401560 6452
rect 492312 6400 492364 6452
rect 313188 6332 313240 6384
rect 371700 6332 371752 6384
rect 398748 6332 398800 6384
rect 488816 6332 488868 6384
rect 489184 6332 489236 6384
rect 498200 6332 498252 6384
rect 262956 6264 263008 6316
rect 300676 6264 300728 6316
rect 314476 6264 314528 6316
rect 374092 6264 374144 6316
rect 404268 6264 404320 6316
rect 495900 6264 495952 6316
rect 269028 6196 269080 6248
rect 311440 6196 311492 6248
rect 322848 6196 322900 6248
rect 384764 6196 384816 6248
rect 407028 6196 407080 6248
rect 499396 6196 499448 6248
rect 274548 6128 274600 6180
rect 318524 6128 318576 6180
rect 324228 6128 324280 6180
rect 387156 6128 387208 6180
rect 408316 6128 408368 6180
rect 502984 6128 503036 6180
rect 382188 6060 382240 6112
rect 466276 6060 466328 6112
rect 342904 5992 342956 6044
rect 391848 5992 391900 6044
rect 393964 5516 394016 5568
rect 396540 5516 396592 5568
rect 475384 5516 475436 5568
rect 480536 5516 480588 5568
rect 486424 5516 486476 5568
rect 487620 5516 487672 5568
rect 493324 5516 493376 5568
rect 494704 5516 494756 5568
rect 512644 5516 512696 5568
rect 513564 5516 513616 5568
rect 269764 5448 269816 5500
rect 292580 5448 292632 5500
rect 354588 5448 354640 5500
rect 427268 5448 427320 5500
rect 435916 5448 435968 5500
rect 540796 5448 540848 5500
rect 268384 5380 268436 5432
rect 297272 5380 297324 5432
rect 351828 5380 351880 5432
rect 423772 5380 423824 5432
rect 438676 5380 438728 5432
rect 544384 5380 544436 5432
rect 256608 5312 256660 5364
rect 293684 5312 293736 5364
rect 304264 5312 304316 5364
rect 310244 5312 310296 5364
rect 355876 5312 355928 5364
rect 430856 5312 430908 5364
rect 444288 5312 444340 5364
rect 551468 5312 551520 5364
rect 267004 5244 267056 5296
rect 306748 5244 306800 5296
rect 307024 5244 307076 5296
rect 346952 5244 347004 5296
rect 358636 5244 358688 5296
rect 434444 5244 434496 5296
rect 441436 5244 441488 5296
rect 547880 5244 547932 5296
rect 271788 5176 271840 5228
rect 313832 5176 313884 5228
rect 364248 5176 364300 5228
rect 441528 5176 441580 5228
rect 449808 5176 449860 5228
rect 558552 5176 558604 5228
rect 271696 5108 271748 5160
rect 315028 5108 315080 5160
rect 361396 5108 361448 5160
rect 437940 5108 437992 5160
rect 447048 5108 447100 5160
rect 554964 5108 555016 5160
rect 242164 5040 242216 5092
rect 271236 5040 271288 5092
rect 281448 5040 281500 5092
rect 328000 5040 328052 5092
rect 367008 5040 367060 5092
rect 445024 5040 445076 5092
rect 452476 5040 452528 5092
rect 562048 5040 562100 5092
rect 234436 4972 234488 5024
rect 264152 4972 264204 5024
rect 267096 4972 267148 5024
rect 267740 4972 267792 5024
rect 286968 4972 287020 5024
rect 335084 4972 335136 5024
rect 372528 4972 372580 5024
rect 452108 4972 452160 5024
rect 455328 4972 455380 5024
rect 565636 4972 565688 5024
rect 224224 4904 224276 4956
rect 242900 4904 242952 4956
rect 250996 4904 251048 4956
rect 285404 4904 285456 4956
rect 285496 4904 285548 4956
rect 332692 4904 332744 4956
rect 369768 4904 369820 4956
rect 448612 4904 448664 4956
rect 456616 4904 456668 4956
rect 569132 4904 569184 4956
rect 213736 4836 213788 4888
rect 235816 4836 235868 4888
rect 238024 4836 238076 4888
rect 239312 4836 239364 4888
rect 253848 4836 253900 4888
rect 290188 4836 290240 4888
rect 292488 4836 292540 4888
rect 342168 4836 342220 4888
rect 375196 4836 375248 4888
rect 455696 4836 455748 4888
rect 462136 4836 462188 4888
rect 576308 4836 576360 4888
rect 227536 4768 227588 4820
rect 253480 4768 253532 4820
rect 260748 4768 260800 4820
rect 299664 4768 299716 4820
rect 303436 4768 303488 4820
rect 357532 4768 357584 4820
rect 376576 4768 376628 4820
rect 459192 4768 459244 4820
rect 459376 4768 459428 4820
rect 572720 4768 572772 4820
rect 251824 4700 251876 4752
rect 274824 4700 274876 4752
rect 289084 4700 289136 4752
rect 276664 4632 276716 4684
rect 296076 4632 296128 4684
rect 349068 4700 349120 4752
rect 420184 4700 420236 4752
rect 434628 4700 434680 4752
rect 537208 4700 537260 4752
rect 307944 4632 307996 4684
rect 346308 4632 346360 4684
rect 416688 4632 416740 4684
rect 431868 4632 431920 4684
rect 533712 4632 533764 4684
rect 273904 4564 273956 4616
rect 288992 4564 289044 4616
rect 343548 4564 343600 4616
rect 413100 4564 413152 4616
rect 429108 4564 429160 4616
rect 530124 4564 530176 4616
rect 262864 4496 262916 4548
rect 278320 4496 278372 4548
rect 287704 4496 287756 4548
rect 303160 4496 303212 4548
rect 337936 4496 337988 4548
rect 406016 4496 406068 4548
rect 423588 4496 423640 4548
rect 523040 4496 523092 4548
rect 340696 4428 340748 4480
rect 409604 4428 409656 4480
rect 426348 4428 426400 4480
rect 526628 4428 526680 4480
rect 244924 4360 244976 4412
rect 249984 4360 250036 4412
rect 335176 4360 335228 4412
rect 402520 4360 402572 4412
rect 420736 4360 420788 4412
rect 519544 4360 519596 4412
rect 333888 4292 333940 4344
rect 398932 4292 398984 4344
rect 418068 4292 418120 4344
rect 515956 4292 516008 4344
rect 331128 4224 331180 4276
rect 395344 4224 395396 4276
rect 415308 4224 415360 4276
rect 512460 4224 512512 4276
rect 255964 4156 256016 4208
rect 257068 4156 257120 4208
rect 318064 4156 318116 4208
rect 320916 4156 320968 4208
rect 327724 4156 327776 4208
rect 329196 4156 329248 4208
rect 522304 4156 522356 4208
rect 524236 4156 524288 4208
rect 26516 4088 26568 4140
rect 60740 4088 60792 4140
rect 168288 4088 168340 4140
rect 171968 4088 172020 4140
rect 186136 4088 186188 4140
rect 196808 4088 196860 4140
rect 204168 4088 204220 4140
rect 221556 4088 221608 4140
rect 223488 4088 223540 4140
rect 247592 4088 247644 4140
rect 248328 4088 248380 4140
rect 283104 4088 283156 4140
rect 291108 4088 291160 4140
rect 340972 4088 341024 4140
rect 347688 4088 347740 4140
rect 350448 4088 350500 4140
rect 422576 4088 422628 4140
rect 424784 4088 424836 4140
rect 424968 4088 425020 4140
rect 441344 4088 441396 4140
rect 546684 4088 546736 4140
rect 574744 4088 574796 4140
rect 577412 4088 577464 4140
rect 17040 3952 17092 4004
rect 53840 3952 53892 4004
rect 20628 3884 20680 3936
rect 182088 4020 182140 4072
rect 190828 4020 190880 4072
rect 191656 4020 191708 4072
rect 203892 4020 203944 4072
rect 205548 4020 205600 4072
rect 223948 4020 224000 4072
rect 226156 4020 226208 4072
rect 252376 4020 252428 4072
rect 252468 4020 252520 4072
rect 287796 4020 287848 4072
rect 299388 4020 299440 4072
rect 351644 4020 351696 4072
rect 353208 4020 353260 4072
rect 426164 4020 426216 4072
rect 442908 4020 442960 4072
rect 550272 4020 550324 4072
rect 81440 3952 81492 4004
rect 161296 3952 161348 4004
rect 163688 3952 163740 4004
rect 169024 3952 169076 4004
rect 173164 3952 173216 4004
rect 179328 3952 179380 4004
rect 187332 3952 187384 4004
rect 190368 3952 190420 4004
rect 202604 3952 202656 4004
rect 202696 3952 202748 4004
rect 220452 3952 220504 4004
rect 220636 3952 220688 4004
rect 245200 3952 245252 4004
rect 249708 3952 249760 4004
rect 284300 3952 284352 4004
rect 296628 3952 296680 4004
rect 348056 3952 348108 4004
rect 358636 3952 358688 4004
rect 11152 3816 11204 3868
rect 49700 3816 49752 3868
rect 56600 3884 56652 3936
rect 69112 3884 69164 3936
rect 91192 3884 91244 3936
rect 177948 3884 178000 3936
rect 186136 3884 186188 3936
rect 188896 3884 188948 3936
rect 200304 3884 200356 3936
rect 205456 3884 205508 3936
rect 222752 3884 222804 3936
rect 223396 3884 223448 3936
rect 248788 3884 248840 3936
rect 251088 3884 251140 3936
rect 286600 3884 286652 3936
rect 303528 3884 303580 3936
rect 358728 3884 358780 3936
rect 429660 3952 429712 4004
rect 448428 3952 448480 4004
rect 557356 3952 557408 4004
rect 433248 3884 433300 3936
rect 445576 3884 445628 3936
rect 553768 3884 553820 3936
rect 12348 3748 12400 3800
rect 7656 3680 7708 3732
rect 2872 3612 2924 3664
rect 42892 3612 42944 3664
rect 64144 3816 64196 3868
rect 65524 3816 65576 3868
rect 89720 3816 89772 3868
rect 180708 3816 180760 3868
rect 189724 3816 189776 3868
rect 191748 3816 191800 3868
rect 205088 3816 205140 3868
rect 206836 3816 206888 3868
rect 225144 3816 225196 3868
rect 227628 3816 227680 3868
rect 254676 3816 254728 3868
rect 255228 3816 255280 3868
rect 291384 3816 291436 3868
rect 300768 3816 300820 3868
rect 355232 3816 355284 3868
rect 355968 3816 356020 3868
rect 361488 3816 361540 3868
rect 436744 3816 436796 3868
rect 451188 3816 451240 3868
rect 560852 3816 560904 3868
rect 56048 3748 56100 3800
rect 56508 3748 56560 3800
rect 61936 3748 61988 3800
rect 87052 3748 87104 3800
rect 183468 3748 183520 3800
rect 193220 3748 193272 3800
rect 194508 3748 194560 3800
rect 208584 3748 208636 3800
rect 211068 3748 211120 3800
rect 231032 3748 231084 3800
rect 231768 3748 231820 3800
rect 259460 3748 259512 3800
rect 262128 3748 262180 3800
rect 301964 3748 302016 3800
rect 306288 3748 306340 3800
rect 362316 3748 362368 3800
rect 362868 3748 362920 3800
rect 440332 3748 440384 3800
rect 453948 3748 454000 3800
rect 564440 3748 564492 3800
rect 56692 3680 56744 3732
rect 58440 3680 58492 3732
rect 84292 3680 84344 3732
rect 179236 3680 179288 3732
rect 188528 3680 188580 3732
rect 188988 3680 189040 3732
rect 201500 3680 201552 3732
rect 206928 3680 206980 3732
rect 226340 3680 226392 3732
rect 230388 3680 230440 3732
rect 258264 3680 258316 3732
rect 259368 3680 259420 3732
rect 298468 3680 298520 3732
rect 311808 3680 311860 3732
rect 369400 3680 369452 3732
rect 371148 3680 371200 3732
rect 450912 3680 450964 3732
rect 456708 3680 456760 3732
rect 568028 3680 568080 3732
rect 49792 3612 49844 3664
rect 54944 3612 54996 3664
rect 5264 3544 5316 3596
rect 45652 3544 45704 3596
rect 51356 3544 51408 3596
rect 78680 3612 78732 3664
rect 85672 3612 85724 3664
rect 86776 3612 86828 3664
rect 170956 3612 171008 3664
rect 175464 3612 175516 3664
rect 176568 3612 176620 3664
rect 183744 3612 183796 3664
rect 184756 3612 184808 3664
rect 195612 3612 195664 3664
rect 195796 3612 195848 3664
rect 209780 3612 209832 3664
rect 212356 3612 212408 3664
rect 232228 3612 232280 3664
rect 234528 3612 234580 3664
rect 262956 3612 263008 3664
rect 264888 3612 264940 3664
rect 305552 3612 305604 3664
rect 308956 3612 309008 3664
rect 365812 3612 365864 3664
rect 368388 3612 368440 3664
rect 447416 3612 447468 3664
rect 448520 3612 448572 3664
rect 449808 3612 449860 3664
rect 459468 3612 459520 3664
rect 571524 3612 571576 3664
rect 1676 3476 1728 3528
rect 572 3408 624 3460
rect 41512 3408 41564 3460
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 46940 3476 46992 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 52552 3476 52604 3528
rect 53656 3476 53708 3528
rect 76104 3544 76156 3596
rect 93952 3544 94004 3596
rect 95056 3544 95108 3596
rect 161388 3544 161440 3596
rect 162492 3544 162544 3596
rect 165436 3544 165488 3596
rect 169576 3544 169628 3596
rect 172336 3544 172388 3596
rect 177856 3544 177908 3596
rect 181996 3544 182048 3596
rect 192024 3544 192076 3596
rect 193036 3544 193088 3596
rect 207388 3544 207440 3596
rect 212448 3544 212500 3596
rect 233424 3544 233476 3596
rect 241336 3544 241388 3596
rect 273628 3544 273680 3596
rect 275928 3544 275980 3596
rect 319720 3544 319772 3596
rect 320088 3544 320140 3596
rect 379980 3544 380032 3596
rect 380808 3544 380860 3596
rect 465172 3544 465224 3596
rect 466184 3544 466236 3596
rect 582196 3544 582248 3596
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 77392 3476 77444 3528
rect 78496 3476 78548 3528
rect 80888 3476 80940 3528
rect 81348 3476 81400 3528
rect 82084 3476 82136 3528
rect 82728 3476 82780 3528
rect 83280 3476 83332 3528
rect 84108 3476 84160 3528
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 89168 3476 89220 3528
rect 89628 3476 89680 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 92388 3476 92440 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 101036 3476 101088 3528
rect 102048 3476 102100 3528
rect 102232 3476 102284 3528
rect 103244 3476 103296 3528
rect 105728 3476 105780 3528
rect 106188 3476 106240 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 109316 3476 109368 3528
rect 110328 3476 110380 3528
rect 110512 3476 110564 3528
rect 111524 3476 111576 3528
rect 114008 3476 114060 3528
rect 114468 3476 114520 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 116400 3476 116452 3528
rect 117228 3476 117280 3528
rect 117596 3476 117648 3528
rect 118608 3476 118660 3528
rect 118792 3476 118844 3528
rect 119988 3476 120040 3528
rect 122288 3476 122340 3528
rect 122748 3476 122800 3528
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 125876 3476 125928 3528
rect 126888 3476 126940 3528
rect 126980 3476 127032 3528
rect 128268 3476 128320 3528
rect 130568 3476 130620 3528
rect 131028 3476 131080 3528
rect 132960 3476 133012 3528
rect 133788 3476 133840 3528
rect 134156 3476 134208 3528
rect 135168 3476 135220 3528
rect 135260 3476 135312 3528
rect 137284 3476 137336 3528
rect 140044 3476 140096 3528
rect 140688 3476 140740 3528
rect 142436 3476 142488 3528
rect 143448 3476 143500 3528
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 149520 3476 149572 3528
rect 150440 3476 150492 3528
rect 153292 3476 153344 3528
rect 154212 3476 154264 3528
rect 155960 3476 156012 3528
rect 156604 3476 156656 3528
rect 157248 3476 157300 3528
rect 157800 3476 157852 3528
rect 158444 3476 158496 3528
rect 158904 3476 158956 3528
rect 160008 3476 160060 3528
rect 161296 3476 161348 3528
rect 164148 3476 164200 3528
rect 167184 3476 167236 3528
rect 169668 3476 169720 3528
rect 174268 3476 174320 3528
rect 187608 3476 187660 3528
rect 199108 3476 199160 3528
rect 199936 3476 199988 3528
rect 216864 3476 216916 3528
rect 217968 3476 218020 3528
rect 240508 3476 240560 3528
rect 241428 3476 241480 3528
rect 272432 3476 272484 3528
rect 273168 3476 273220 3528
rect 316224 3476 316276 3528
rect 317420 3476 317472 3528
rect 376484 3476 376536 3528
rect 376668 3476 376720 3528
rect 458088 3476 458140 3528
rect 462228 3476 462280 3528
rect 575112 3476 575164 3528
rect 42892 3408 42944 3460
rect 44272 3408 44324 3460
rect 8760 3340 8812 3392
rect 9588 3340 9640 3392
rect 15936 3340 15988 3392
rect 16488 3340 16540 3392
rect 18236 3340 18288 3392
rect 19248 3340 19300 3392
rect 24216 3340 24268 3392
rect 24768 3340 24820 3392
rect 25320 3340 25372 3392
rect 26148 3340 26200 3392
rect 27712 3340 27764 3392
rect 28908 3340 28960 3392
rect 32404 3340 32456 3392
rect 33048 3340 33100 3392
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 9956 3272 10008 3324
rect 43444 3272 43496 3324
rect 46664 3272 46716 3324
rect 57244 3340 57296 3392
rect 57888 3340 57940 3392
rect 59636 3340 59688 3392
rect 60648 3340 60700 3392
rect 60832 3340 60884 3392
rect 62028 3340 62080 3392
rect 64328 3340 64380 3392
rect 64788 3340 64840 3392
rect 66720 3408 66772 3460
rect 67548 3408 67600 3460
rect 67916 3408 67968 3460
rect 68928 3408 68980 3460
rect 72608 3408 72660 3460
rect 73068 3408 73120 3460
rect 73804 3408 73856 3460
rect 74448 3408 74500 3460
rect 131764 3408 131816 3460
rect 132408 3408 132460 3460
rect 158536 3408 158588 3460
rect 160100 3408 160152 3460
rect 166908 3408 166960 3460
rect 170772 3408 170824 3460
rect 171048 3408 171100 3460
rect 176660 3408 176712 3460
rect 177764 3408 177816 3460
rect 184940 3408 184992 3460
rect 186228 3408 186280 3460
rect 197912 3408 197964 3460
rect 198556 3408 198608 3460
rect 214472 3408 214524 3460
rect 215208 3408 215260 3460
rect 237012 3408 237064 3460
rect 240048 3408 240100 3460
rect 270040 3408 270092 3460
rect 270408 3408 270460 3460
rect 307760 3408 307812 3460
rect 309048 3408 309100 3460
rect 314568 3408 314620 3460
rect 372896 3408 372948 3460
rect 373908 3408 373960 3460
rect 454500 3408 454552 3460
rect 463608 3408 463660 3460
rect 578608 3408 578660 3460
rect 73436 3340 73488 3392
rect 173808 3340 173860 3392
rect 180248 3340 180300 3392
rect 184848 3340 184900 3392
rect 194416 3340 194468 3392
rect 201408 3340 201460 3392
rect 218060 3340 218112 3392
rect 219348 3340 219400 3392
rect 241704 3340 241756 3392
rect 244004 3340 244056 3392
rect 277124 3340 277176 3392
rect 293868 3340 293920 3392
rect 344560 3340 344612 3392
rect 344928 3340 344980 3392
rect 415492 3340 415544 3392
rect 438768 3340 438820 3392
rect 543188 3340 543240 3392
rect 551284 3340 551336 3392
rect 552664 3340 552716 3392
rect 558184 3340 558236 3392
rect 559748 3340 559800 3392
rect 63592 3272 63644 3324
rect 138848 3272 138900 3324
rect 139308 3272 139360 3324
rect 200028 3272 200080 3324
rect 215668 3272 215720 3324
rect 220728 3272 220780 3324
rect 244096 3272 244148 3324
rect 246948 3272 247000 3324
rect 279516 3272 279568 3324
rect 288348 3272 288400 3324
rect 337476 3272 337528 3324
rect 349160 3272 349212 3324
rect 350448 3272 350500 3324
rect 418988 3272 419040 3324
rect 436008 3272 436060 3324
rect 539600 3272 539652 3324
rect 21824 3204 21876 3256
rect 33600 3204 33652 3256
rect 66352 3204 66404 3256
rect 172428 3204 172480 3256
rect 179052 3204 179104 3256
rect 195888 3204 195940 3256
rect 210976 3204 211028 3256
rect 216588 3204 216640 3256
rect 238116 3204 238168 3256
rect 244188 3204 244240 3256
rect 276020 3204 276072 3256
rect 285588 3204 285640 3256
rect 333888 3204 333940 3256
rect 342076 3204 342128 3256
rect 411904 3204 411956 3256
rect 433156 3204 433208 3256
rect 536104 3204 536156 3256
rect 569224 3204 569276 3256
rect 570328 3204 570380 3256
rect 30104 3136 30156 3188
rect 37188 3068 37240 3120
rect 69204 3136 69256 3188
rect 165528 3136 165580 3188
rect 168380 3136 168432 3188
rect 175096 3136 175148 3188
rect 181444 3136 181496 3188
rect 197268 3136 197320 3188
rect 212172 3136 212224 3188
rect 213828 3136 213880 3188
rect 234620 3136 234672 3188
rect 237288 3136 237340 3188
rect 266544 3136 266596 3188
rect 278688 3136 278740 3188
rect 323308 3136 323360 3188
rect 324320 3136 324372 3188
rect 325608 3136 325660 3188
rect 340788 3136 340840 3188
rect 408408 3136 408460 3188
rect 427728 3136 427780 3188
rect 529020 3136 529072 3188
rect 40684 3068 40736 3120
rect 70492 3068 70544 3120
rect 193128 3068 193180 3120
rect 206192 3068 206244 3120
rect 209688 3068 209740 3120
rect 229836 3068 229888 3120
rect 235908 3068 235960 3120
rect 265348 3068 265400 3120
rect 312636 3068 312688 3120
rect 338028 3068 338080 3120
rect 404820 3068 404872 3120
rect 430488 3068 430540 3120
rect 532516 3068 532568 3120
rect 19432 3000 19484 3052
rect 46204 3000 46256 3052
rect 47860 3000 47912 3052
rect 148324 3000 148376 3052
rect 148968 3000 149020 3052
rect 162768 3000 162820 3052
rect 164884 3000 164936 3052
rect 209596 3000 209648 3052
rect 228732 3000 228784 3052
rect 238668 3000 238720 3052
rect 268844 3000 268896 3052
rect 335268 3000 335320 3052
rect 28908 2932 28960 2984
rect 48872 2932 48924 2984
rect 141240 2932 141292 2984
rect 142068 2932 142120 2984
rect 175188 2932 175240 2984
rect 182548 2932 182600 2984
rect 208308 2932 208360 2984
rect 227536 2932 227588 2984
rect 233148 2932 233200 2984
rect 261760 2932 261812 2984
rect 332508 2932 332560 2984
rect 397736 2932 397788 2984
rect 398840 3000 398892 3052
rect 400128 3000 400180 3052
rect 422116 3000 422168 3052
rect 521844 3000 521896 3052
rect 560944 3000 560996 3052
rect 563244 3000 563296 3052
rect 401324 2932 401376 2984
rect 424784 2932 424836 2984
rect 525432 2932 525484 2984
rect 35992 2864 36044 2916
rect 55864 2864 55916 2916
rect 202788 2864 202840 2916
rect 219256 2864 219308 2916
rect 229008 2864 229060 2916
rect 255872 2864 255924 2916
rect 329748 2864 329800 2916
rect 394240 2864 394292 2916
rect 420828 2864 420880 2916
rect 518348 2864 518400 2916
rect 43076 2796 43128 2848
rect 62764 2796 62816 2848
rect 198648 2796 198700 2848
rect 213368 2796 213420 2848
rect 226248 2796 226300 2848
rect 251180 2796 251232 2848
rect 321468 2796 321520 2848
rect 383568 2796 383620 2848
rect 383660 2796 383712 2848
rect 468668 2796 468720 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 8128 700466 8156 703520
rect 24320 700534 24348 703520
rect 40512 700602 40540 703520
rect 72988 700806 73016 703520
rect 89180 700874 89208 703520
rect 89168 700868 89220 700874
rect 89168 700810 89220 700816
rect 72976 700800 73028 700806
rect 72976 700742 73028 700748
rect 40500 700596 40552 700602
rect 40500 700538 40552 700544
rect 24308 700528 24360 700534
rect 24308 700470 24360 700476
rect 8116 700460 8168 700466
rect 8116 700402 8168 700408
rect 105464 699718 105492 703520
rect 137848 700262 137876 703520
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 154132 700194 154160 703520
rect 154120 700188 154172 700194
rect 154120 700130 154172 700136
rect 170324 699718 170352 703520
rect 202800 699990 202828 703520
rect 215208 700392 215260 700398
rect 215208 700334 215260 700340
rect 202788 699984 202840 699990
rect 202788 699926 202840 699932
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 670818 3464 671191
rect 3424 670812 3476 670818
rect 3424 670754 3476 670760
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 22836 472184 22888 472190
rect 22836 472126 22888 472132
rect 3608 470144 3660 470150
rect 3608 470086 3660 470092
rect 3516 468240 3568 468246
rect 3516 468182 3568 468188
rect 3424 463684 3476 463690
rect 3424 463626 3476 463632
rect 3436 462641 3464 463626
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 3528 462482 3556 468182
rect 3436 462454 3556 462482
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3240 398812 3292 398818
rect 3240 398754 3292 398760
rect 3252 397497 3280 398754
rect 3238 397488 3294 397497
rect 3238 397423 3294 397432
rect 2780 371408 2832 371414
rect 2778 371376 2780 371385
rect 2832 371376 2834 371385
rect 2778 371311 2834 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3436 241097 3464 462454
rect 3620 451274 3648 470086
rect 15844 470008 15896 470014
rect 15844 469950 15896 469956
rect 7564 469464 7616 469470
rect 7564 469406 7616 469412
rect 4896 468716 4948 468722
rect 4896 468658 4948 468664
rect 4804 468036 4856 468042
rect 4804 467978 4856 467984
rect 3528 451246 3648 451274
rect 3528 423609 3556 451246
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3516 320136 3568 320142
rect 3516 320078 3568 320084
rect 3528 319297 3556 320078
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 4816 137154 4844 467978
rect 4908 371414 4936 468658
rect 4896 371408 4948 371414
rect 4896 371350 4948 371356
rect 2780 137148 2832 137154
rect 2780 137090 2832 137096
rect 4804 137148 4856 137154
rect 4804 137090 4856 137096
rect 2792 136785 2820 137090
rect 2778 136776 2834 136785
rect 2778 136711 2834 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 7576 85542 7604 469406
rect 11704 469260 11756 469266
rect 11704 469202 11756 469208
rect 7656 468648 7708 468654
rect 7656 468590 7708 468596
rect 7668 346390 7696 468590
rect 7656 346384 7708 346390
rect 7656 346326 7708 346332
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 7564 85536 7616 85542
rect 7564 85478 7616 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 6828 39500 6880 39506
rect 6828 39442 6880 39448
rect 4068 39364 4120 39370
rect 4068 39306 4120 39312
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 2884 480 2912 3606
rect 4080 480 4108 39306
rect 6840 6914 6868 39442
rect 9588 39432 9640 39438
rect 9588 39374 9640 39380
rect 6472 6886 6868 6914
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5276 480 5304 3538
rect 6472 480 6500 6886
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7668 480 7696 3674
rect 9600 3398 9628 39374
rect 11716 33114 11744 469202
rect 14464 468512 14516 468518
rect 14464 468454 14516 468460
rect 13818 467800 13874 467809
rect 13818 467735 13874 467744
rect 13832 463690 13860 467735
rect 13820 463684 13872 463690
rect 13820 463626 13872 463632
rect 14476 267714 14504 468454
rect 15856 293962 15884 469950
rect 18604 469872 18656 469878
rect 18604 469814 18656 469820
rect 17224 469736 17276 469742
rect 17224 469678 17276 469684
rect 15936 468988 15988 468994
rect 15936 468930 15988 468936
rect 15948 449886 15976 468930
rect 15936 449880 15988 449886
rect 15936 449822 15988 449828
rect 15844 293956 15896 293962
rect 15844 293898 15896 293904
rect 14464 267708 14516 267714
rect 14464 267650 14516 267656
rect 17236 189038 17264 469678
rect 17316 468852 17368 468858
rect 17316 468794 17368 468800
rect 17328 398818 17356 468794
rect 17316 398812 17368 398818
rect 17316 398754 17368 398760
rect 18616 215286 18644 469814
rect 21364 469600 21416 469606
rect 21364 469542 21416 469548
rect 18604 215280 18656 215286
rect 18604 215222 18656 215228
rect 17224 189032 17276 189038
rect 17224 188974 17276 188980
rect 21376 111790 21404 469542
rect 22744 467968 22796 467974
rect 22744 467910 22796 467916
rect 21364 111784 21416 111790
rect 21364 111726 21416 111732
rect 22756 71738 22784 467910
rect 22848 358766 22876 472126
rect 85120 472048 85172 472054
rect 85120 471990 85172 471996
rect 81348 471708 81400 471714
rect 81348 471650 81400 471656
rect 29736 471096 29788 471102
rect 29736 471038 29788 471044
rect 29644 469396 29696 469402
rect 29644 469338 29696 469344
rect 25504 468308 25556 468314
rect 25504 468250 25556 468256
rect 22836 358760 22888 358766
rect 22836 358702 22888 358708
rect 25516 164218 25544 468250
rect 25504 164212 25556 164218
rect 25504 164154 25556 164160
rect 22744 71732 22796 71738
rect 22744 71674 22796 71680
rect 26148 40044 26200 40050
rect 26148 39986 26200 39992
rect 24768 39908 24820 39914
rect 24768 39850 24820 39856
rect 23388 39840 23440 39846
rect 23388 39782 23440 39788
rect 16488 39772 16540 39778
rect 16488 39714 16540 39720
rect 15108 39636 15160 39642
rect 15108 39578 15160 39584
rect 13728 39568 13780 39574
rect 13728 39510 13780 39516
rect 11704 33108 11756 33114
rect 11704 33050 11756 33056
rect 13740 6914 13768 39510
rect 15120 6914 15148 39578
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 11152 3868 11204 3874
rect 11152 3810 11204 3816
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 8772 480 8800 3334
rect 9956 3324 10008 3330
rect 9956 3266 10008 3272
rect 9968 480 9996 3266
rect 11164 480 11192 3810
rect 12348 3800 12400 3806
rect 12348 3742 12400 3748
rect 12360 480 12388 3742
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3398 16528 39714
rect 19248 39704 19300 39710
rect 19248 39646 19300 39652
rect 17040 4004 17092 4010
rect 17040 3946 17092 3952
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 15948 480 15976 3334
rect 17052 480 17080 3946
rect 19260 3398 19288 39646
rect 23400 6914 23428 39782
rect 23032 6886 23428 6914
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 18248 480 18276 3334
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 480 19472 2994
rect 20640 480 20668 3878
rect 21824 3256 21876 3262
rect 21824 3198 21876 3204
rect 21836 480 21864 3198
rect 23032 480 23060 6886
rect 24780 3398 24808 39850
rect 26160 3398 26188 39986
rect 28908 39976 28960 39982
rect 28908 39918 28960 39924
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 24228 480 24256 3334
rect 25332 480 25360 3334
rect 26528 480 26556 4082
rect 28920 3398 28948 39918
rect 29656 6866 29684 469338
rect 29748 255270 29776 471038
rect 32404 471028 32456 471034
rect 32404 470970 32456 470976
rect 29736 255264 29788 255270
rect 29736 255206 29788 255212
rect 32416 202842 32444 470970
rect 33784 470960 33836 470966
rect 33784 470902 33836 470908
rect 32404 202836 32456 202842
rect 32404 202778 32456 202784
rect 33796 150414 33824 470902
rect 35164 470824 35216 470830
rect 35164 470766 35216 470772
rect 33784 150408 33836 150414
rect 33784 150350 33836 150356
rect 35176 97986 35204 470766
rect 36544 470756 36596 470762
rect 36544 470698 36596 470704
rect 35254 467664 35310 467673
rect 35254 467599 35310 467608
rect 35268 306338 35296 467599
rect 35256 306332 35308 306338
rect 35256 306274 35308 306280
rect 35164 97980 35216 97986
rect 35164 97922 35216 97928
rect 36556 59362 36584 470698
rect 40684 470620 40736 470626
rect 40684 470562 40736 470568
rect 39396 470348 39448 470354
rect 39396 470290 39448 470296
rect 39304 468172 39356 468178
rect 39304 468114 39356 468120
rect 36544 59356 36596 59362
rect 36544 59298 36596 59304
rect 39316 45558 39344 468114
rect 39408 320142 39436 470290
rect 39396 320136 39448 320142
rect 39396 320078 39448 320084
rect 39304 45552 39356 45558
rect 39304 45494 39356 45500
rect 31668 39296 31720 39302
rect 31668 39238 31720 39244
rect 31680 6914 31708 39238
rect 33048 39228 33100 39234
rect 33048 39170 33100 39176
rect 31312 6886 31708 6914
rect 29644 6860 29696 6866
rect 29644 6802 29696 6808
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27724 480 27752 3334
rect 30104 3188 30156 3194
rect 30104 3130 30156 3136
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 28920 480 28948 2926
rect 30116 480 30144 3130
rect 31312 480 31340 6886
rect 33060 3398 33088 39170
rect 38568 39160 38620 39166
rect 38568 39102 38620 39108
rect 35808 39092 35860 39098
rect 35808 39034 35860 39040
rect 35820 3398 35848 39034
rect 38580 6914 38608 39102
rect 39948 39024 40000 39030
rect 39948 38966 40000 38972
rect 39960 6914 39988 38966
rect 40696 20670 40724 470562
rect 65984 469668 66036 469674
rect 65984 469610 66036 469616
rect 58992 469328 59044 469334
rect 58992 469270 59044 469276
rect 59004 468602 59032 469270
rect 58696 468574 59032 468602
rect 65996 468330 66024 469610
rect 70216 469532 70268 469538
rect 70216 469474 70268 469480
rect 70228 468602 70256 469474
rect 81360 468602 81388 471650
rect 85132 468602 85160 471990
rect 106200 471646 106228 699654
rect 170956 536852 171008 536858
rect 170956 536794 171008 536800
rect 166908 510672 166960 510678
rect 166908 510614 166960 510620
rect 160008 484424 160060 484430
rect 160008 484366 160060 484372
rect 129648 472116 129700 472122
rect 129648 472058 129700 472064
rect 106188 471640 106240 471646
rect 106188 471582 106240 471588
rect 118608 471300 118660 471306
rect 118608 471242 118660 471248
rect 107476 471232 107528 471238
rect 107476 471174 107528 471180
rect 96252 471164 96304 471170
rect 96252 471106 96304 471112
rect 92388 470892 92440 470898
rect 92388 470834 92440 470840
rect 88800 469940 88852 469946
rect 88800 469882 88852 469888
rect 88812 468602 88840 469882
rect 92400 468602 92428 470834
rect 96264 468602 96292 471106
rect 103244 469804 103296 469810
rect 103244 469746 103296 469752
rect 69920 468574 70256 468602
rect 81052 468574 81388 468602
rect 84824 468574 85160 468602
rect 88504 468574 88840 468602
rect 92276 468574 92428 468602
rect 95956 468574 96292 468602
rect 99728 468586 100064 468602
rect 99728 468580 100076 468586
rect 99728 468574 100024 468580
rect 100024 468522 100076 468528
rect 77668 468376 77720 468382
rect 65996 468302 66148 468330
rect 77372 468324 77668 468330
rect 77372 468318 77720 468324
rect 103256 468330 103284 469746
rect 107488 468602 107516 471174
rect 111156 470076 111208 470082
rect 111156 470018 111208 470024
rect 111168 468602 111196 470018
rect 118620 468602 118648 471242
rect 122380 468784 122432 468790
rect 122380 468726 122432 468732
rect 122392 468602 122420 468726
rect 129660 468602 129688 472058
rect 160020 471986 160048 484366
rect 159548 471980 159600 471986
rect 159548 471922 159600 471928
rect 160008 471980 160060 471986
rect 160008 471922 160060 471928
rect 148416 471572 148468 471578
rect 148416 471514 148468 471520
rect 140688 471436 140740 471442
rect 140688 471378 140740 471384
rect 133512 470280 133564 470286
rect 133512 470222 133564 470228
rect 133524 468602 133552 470222
rect 140700 468874 140728 471378
rect 107180 468574 107516 468602
rect 110860 468574 111196 468602
rect 118312 468574 118648 468602
rect 122084 468574 122420 468602
rect 129536 468574 129688 468602
rect 133216 468574 133552 468602
rect 140654 468846 140728 468874
rect 144736 468920 144788 468926
rect 144736 468862 144788 468868
rect 140654 468588 140682 468846
rect 144748 468602 144776 468862
rect 148428 468602 148456 471514
rect 155868 470416 155920 470422
rect 155868 470358 155920 470364
rect 152096 469056 152148 469062
rect 152096 468998 152148 469004
rect 152108 468602 152136 468998
rect 155880 468602 155908 470358
rect 159560 468602 159588 471922
rect 163320 470688 163372 470694
rect 163320 470630 163372 470636
rect 163332 468602 163360 470630
rect 166920 468602 166948 510614
rect 170968 470594 170996 536794
rect 171060 471782 171088 699654
rect 204168 696992 204220 696998
rect 204168 696934 204220 696940
rect 201408 670744 201460 670750
rect 201408 670686 201460 670692
rect 193128 643136 193180 643142
rect 193128 643078 193180 643084
rect 190368 616888 190420 616894
rect 190368 616830 190420 616836
rect 182088 590708 182140 590714
rect 182088 590650 182140 590656
rect 177948 563100 178000 563106
rect 177948 563042 178000 563048
rect 175188 524476 175240 524482
rect 175188 524418 175240 524424
rect 175200 471986 175228 524418
rect 174452 471980 174504 471986
rect 174452 471922 174504 471928
rect 175188 471980 175240 471986
rect 175188 471922 175240 471928
rect 171048 471776 171100 471782
rect 171048 471718 171100 471724
rect 170876 470566 170996 470594
rect 170876 468602 170904 470566
rect 174464 468602 174492 471922
rect 177960 468874 177988 563042
rect 182100 470594 182128 590650
rect 186228 576904 186280 576910
rect 186228 576846 186280 576852
rect 186240 471986 186268 576846
rect 190380 471986 190408 616830
rect 185676 471980 185728 471986
rect 185676 471922 185728 471928
rect 186228 471980 186280 471986
rect 186228 471922 186280 471928
rect 189356 471980 189408 471986
rect 189356 471922 189408 471928
rect 190368 471980 190420 471986
rect 190368 471922 190420 471928
rect 144440 468574 144776 468602
rect 148120 468574 148456 468602
rect 151800 468574 152136 468602
rect 155572 468574 155908 468602
rect 159252 468574 159588 468602
rect 163024 468574 163360 468602
rect 166704 468574 166948 468602
rect 170476 468574 170904 468602
rect 174156 468574 174492 468602
rect 177914 468846 177988 468874
rect 182008 470566 182128 470594
rect 177914 468588 177942 468846
rect 182008 468602 182036 470566
rect 185688 468602 185716 471922
rect 189368 468602 189396 471922
rect 193140 468602 193168 643078
rect 197268 630692 197320 630698
rect 197268 630634 197320 630640
rect 197280 471986 197308 630634
rect 201420 471986 201448 670686
rect 196808 471980 196860 471986
rect 196808 471922 196860 471928
rect 197268 471980 197320 471986
rect 197268 471922 197320 471928
rect 200580 471980 200632 471986
rect 200580 471922 200632 471928
rect 201408 471980 201460 471986
rect 201408 471922 201460 471928
rect 196820 468602 196848 471922
rect 200592 468602 200620 471922
rect 204180 468602 204208 696934
rect 208308 683188 208360 683194
rect 208308 683130 208360 683136
rect 208320 470594 208348 683130
rect 211712 471368 211764 471374
rect 211712 471310 211764 471316
rect 208136 470566 208348 470594
rect 208136 468602 208164 470566
rect 211724 468602 211752 471310
rect 215220 468874 215248 700334
rect 218992 699922 219020 703520
rect 227628 700732 227680 700738
rect 227628 700674 227680 700680
rect 219348 700324 219400 700330
rect 219348 700266 219400 700272
rect 218980 699916 219032 699922
rect 218980 699858 219032 699864
rect 219360 470594 219388 700266
rect 227640 471986 227668 700674
rect 230388 700664 230440 700670
rect 230388 700606 230440 700612
rect 226616 471980 226668 471986
rect 226616 471922 226668 471928
rect 227628 471980 227680 471986
rect 227628 471922 227680 471928
rect 223396 471572 223448 471578
rect 223396 471514 223448 471520
rect 222936 471504 222988 471510
rect 222936 471446 222988 471452
rect 181608 468574 182036 468602
rect 185380 468574 185716 468602
rect 189060 468574 189396 468602
rect 192832 468574 193168 468602
rect 196512 468574 196848 468602
rect 200284 468574 200620 468602
rect 203964 468574 204208 468602
rect 207736 468574 208164 468602
rect 211416 468574 211752 468602
rect 215174 468846 215248 468874
rect 219268 470566 219388 470594
rect 215174 468588 215202 468846
rect 219268 468602 219296 470566
rect 222948 468602 222976 471446
rect 223408 470218 223436 471514
rect 223396 470212 223448 470218
rect 223396 470154 223448 470160
rect 226628 468602 226656 471922
rect 230400 468602 230428 700606
rect 235184 699718 235212 703520
rect 238668 701004 238720 701010
rect 238668 700946 238720 700952
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 235920 471918 235948 699654
rect 235908 471912 235960 471918
rect 235908 471854 235960 471860
rect 238680 471714 238708 700946
rect 241428 700936 241480 700942
rect 241428 700878 241480 700884
rect 234068 471708 234120 471714
rect 234068 471650 234120 471656
rect 237840 471708 237892 471714
rect 237840 471650 237892 471656
rect 238668 471708 238720 471714
rect 238668 471650 238720 471656
rect 234080 468602 234108 471650
rect 234988 471572 235040 471578
rect 234988 471514 235040 471520
rect 235000 469062 235028 471514
rect 234988 469056 235040 469062
rect 234988 468998 235040 469004
rect 237852 468602 237880 471650
rect 241440 468602 241468 700878
rect 252468 700120 252520 700126
rect 252468 700062 252520 700068
rect 249708 700052 249760 700058
rect 249708 699994 249760 700000
rect 249720 471986 249748 699994
rect 248972 471980 249024 471986
rect 248972 471922 249024 471928
rect 249708 471980 249760 471986
rect 249708 471922 249760 471928
rect 245292 471708 245344 471714
rect 245292 471650 245344 471656
rect 245304 468602 245332 471650
rect 248984 468602 249012 471922
rect 252480 468874 252508 700062
rect 264888 699848 264940 699854
rect 264888 699790 264940 699796
rect 260748 699712 260800 699718
rect 260748 699654 260800 699660
rect 260760 471986 260788 699654
rect 264900 471986 264928 699790
rect 267660 699718 267688 703520
rect 281540 700256 281592 700262
rect 281540 700198 281592 700204
rect 270500 699984 270552 699990
rect 270500 699926 270552 699932
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 270512 480254 270540 699926
rect 274640 699916 274692 699922
rect 274640 699858 274692 699864
rect 270512 480226 270632 480254
rect 260104 471980 260156 471986
rect 260104 471922 260156 471928
rect 260748 471980 260800 471986
rect 260748 471922 260800 471928
rect 263876 471980 263928 471986
rect 263876 471922 263928 471928
rect 264888 471980 264940 471986
rect 264888 471922 264940 471928
rect 256424 471844 256476 471850
rect 256424 471786 256476 471792
rect 218868 468574 219296 468602
rect 222640 468574 222976 468602
rect 226320 468574 226656 468602
rect 230092 468574 230428 468602
rect 233772 468574 234108 468602
rect 237544 468574 237880 468602
rect 241224 468574 241468 468602
rect 244996 468574 245332 468602
rect 248676 468574 249012 468602
rect 252434 468846 252508 468874
rect 252434 468588 252462 468846
rect 256436 468602 256464 471786
rect 260116 468602 260144 471922
rect 263888 468602 263916 471922
rect 266912 471912 266964 471918
rect 266912 471854 266964 471860
rect 256128 468574 256464 468602
rect 259808 468574 260144 468602
rect 263580 468574 263916 468602
rect 266924 468602 266952 471854
rect 270604 468602 270632 480226
rect 274652 468874 274680 699858
rect 281552 480254 281580 700198
rect 283852 699854 283880 703520
rect 296720 700868 296772 700874
rect 296720 700810 296772 700816
rect 292580 700800 292632 700806
rect 292580 700742 292632 700748
rect 285680 700188 285732 700194
rect 285680 700130 285732 700136
rect 283840 699848 283892 699854
rect 283840 699790 283892 699796
rect 281552 480226 281764 480254
rect 278136 471776 278188 471782
rect 278136 471718 278188 471724
rect 274652 468846 274726 468874
rect 266924 468574 267260 468602
rect 270604 468574 271032 468602
rect 274698 468588 274726 468846
rect 278148 468602 278176 471718
rect 281736 468602 281764 480226
rect 285692 468602 285720 700130
rect 292592 480254 292620 700742
rect 292592 480226 292988 480254
rect 289268 471640 289320 471646
rect 289268 471582 289320 471588
rect 289280 468602 289308 471582
rect 292960 468602 292988 480226
rect 296732 468602 296760 700810
rect 299492 471850 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 300860 700596 300912 700602
rect 300860 700538 300912 700544
rect 299480 471844 299532 471850
rect 299480 471786 299532 471792
rect 300872 468874 300900 700538
rect 307760 700528 307812 700534
rect 307760 700470 307812 700476
rect 303620 700460 303672 700466
rect 303620 700402 303672 700408
rect 303632 480254 303660 700402
rect 307772 480254 307800 700470
rect 332520 700058 332548 703520
rect 348804 700126 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700120 348844 700126
rect 348792 700062 348844 700068
rect 332508 700052 332560 700058
rect 332508 699994 332560 700000
rect 311900 683256 311952 683262
rect 311900 683198 311952 683204
rect 303632 480226 304120 480254
rect 307772 480226 307892 480254
rect 300826 468846 300900 468874
rect 278148 468574 278484 468602
rect 281736 468574 282164 468602
rect 285692 468574 285936 468602
rect 289280 468574 289616 468602
rect 292960 468574 293388 468602
rect 296732 468574 297068 468602
rect 300826 468588 300854 468846
rect 304092 468602 304120 480226
rect 307864 468602 307892 480226
rect 311912 468874 311940 683198
rect 318800 670812 318852 670818
rect 318800 670754 318852 670760
rect 314660 656940 314712 656946
rect 314660 656882 314712 656888
rect 314672 480254 314700 656882
rect 318812 480254 318840 670754
rect 322940 632120 322992 632126
rect 322940 632062 322992 632068
rect 314672 480226 315344 480254
rect 318812 480226 319024 480254
rect 311912 468846 311986 468874
rect 304092 468574 304520 468602
rect 307864 468574 308292 468602
rect 311958 468588 311986 468846
rect 315316 468602 315344 480226
rect 318996 468602 319024 480226
rect 322952 468602 322980 632062
rect 329840 618316 329892 618322
rect 329840 618258 329892 618264
rect 325700 605872 325752 605878
rect 325700 605814 325752 605820
rect 325712 480254 325740 605814
rect 329852 480254 329880 618258
rect 333980 579692 334032 579698
rect 333980 579634 334032 579640
rect 325712 480226 326476 480254
rect 329852 480226 330248 480254
rect 326448 468602 326476 480226
rect 330220 468602 330248 480226
rect 333992 468602 334020 579634
rect 340880 565888 340932 565894
rect 340880 565830 340932 565836
rect 338120 553444 338172 553450
rect 338120 553386 338172 553392
rect 338132 468874 338160 553386
rect 340892 480254 340920 565830
rect 345020 527196 345072 527202
rect 345020 527138 345072 527144
rect 345032 480254 345060 527138
rect 351920 514820 351972 514826
rect 351920 514762 351972 514768
rect 349160 501016 349212 501022
rect 349160 500958 349212 500964
rect 340892 480226 341380 480254
rect 345032 480226 345152 480254
rect 338086 468846 338160 468874
rect 315316 468574 315744 468602
rect 318996 468574 319424 468602
rect 322952 468574 323196 468602
rect 326448 468574 326876 468602
rect 330220 468574 330648 468602
rect 333992 468574 334328 468602
rect 338086 468588 338114 468846
rect 341352 468602 341380 480226
rect 345124 468602 345152 480226
rect 349172 468874 349200 500958
rect 351932 480254 351960 514762
rect 351932 480226 352604 480254
rect 349172 468846 349246 468874
rect 341352 468574 341780 468602
rect 345124 468574 345552 468602
rect 349218 468588 349246 468846
rect 352576 468602 352604 480226
rect 356244 474768 356296 474774
rect 356244 474710 356296 474716
rect 356256 468602 356284 474710
rect 364352 471714 364380 702406
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 413664 700942 413692 703520
rect 413652 700936 413704 700942
rect 413652 700878 413704 700884
rect 386420 472184 386472 472190
rect 386420 472126 386472 472132
rect 364340 471708 364392 471714
rect 364340 471650 364392 471656
rect 367468 470144 367520 470150
rect 367468 470086 367520 470092
rect 360200 468988 360252 468994
rect 360200 468930 360252 468936
rect 360212 468602 360240 468930
rect 367480 468602 367508 470086
rect 386432 468874 386460 472126
rect 429212 471578 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700738 462360 703520
rect 462320 700732 462372 700738
rect 462320 700674 462372 700680
rect 478524 700670 478552 703520
rect 478512 700664 478564 700670
rect 478512 700606 478564 700612
rect 429200 471572 429252 471578
rect 429200 471514 429252 471520
rect 494072 471510 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 512644 472116 512696 472122
rect 512644 472058 512696 472064
rect 511264 472048 511316 472054
rect 511264 471990 511316 471996
rect 494060 471504 494112 471510
rect 494060 471446 494112 471452
rect 467380 471436 467432 471442
rect 467380 471378 467432 471384
rect 467288 471300 467340 471306
rect 467288 471242 467340 471248
rect 467196 471232 467248 471238
rect 467196 471174 467248 471180
rect 467104 471164 467156 471170
rect 467104 471106 467156 471112
rect 408500 471096 408552 471102
rect 408500 471038 408552 471044
rect 389824 470348 389876 470354
rect 389824 470290 389876 470296
rect 371562 468852 371614 468858
rect 386432 468846 386506 468874
rect 371562 468794 371614 468800
rect 352576 468574 353004 468602
rect 356256 468574 356684 468602
rect 360212 468574 360456 468602
rect 367480 468574 367816 468602
rect 371574 468588 371602 468794
rect 378692 468716 378744 468722
rect 378692 468658 378744 468664
rect 378704 468602 378732 468658
rect 382372 468648 382424 468654
rect 378704 468574 379040 468602
rect 382424 468596 382720 468602
rect 382372 468590 382720 468596
rect 382384 468574 382720 468590
rect 386478 468588 386506 468846
rect 389836 468602 389864 470290
rect 393596 470008 393648 470014
rect 393596 469950 393648 469956
rect 393608 468602 393636 469950
rect 408512 468602 408540 471038
rect 419632 471028 419684 471034
rect 419632 470970 419684 470976
rect 412180 469872 412232 469878
rect 412180 469814 412232 469820
rect 412192 468602 412220 469814
rect 415952 469736 416004 469742
rect 415952 469678 416004 469684
rect 415964 468602 415992 469678
rect 419644 468602 419672 470970
rect 430856 470960 430908 470966
rect 430856 470902 430908 470908
rect 430868 468602 430896 470902
rect 441988 470824 442040 470830
rect 441988 470766 442040 470772
rect 434720 469600 434772 469606
rect 434720 469542 434772 469548
rect 434732 468602 434760 469542
rect 438308 469464 438360 469470
rect 438308 469406 438360 469412
rect 438320 468602 438348 469406
rect 442000 468602 442028 470766
rect 453212 470756 453264 470762
rect 453212 470698 453264 470704
rect 453224 468602 453252 470698
rect 464344 470620 464396 470626
rect 464344 470562 464396 470568
rect 461124 469396 461176 469402
rect 461124 469338 461176 469344
rect 456892 469260 456944 469266
rect 456892 469202 456944 469208
rect 456904 468602 456932 469202
rect 389836 468574 390172 468602
rect 393608 468574 393944 468602
rect 408512 468574 408848 468602
rect 412192 468574 412528 468602
rect 415964 468574 416300 468602
rect 419644 468574 419980 468602
rect 430868 468574 431204 468602
rect 434732 468574 434884 468602
rect 438320 468574 438656 468602
rect 442000 468574 442336 468602
rect 453224 468574 453560 468602
rect 456904 468574 457240 468602
rect 401048 468512 401100 468518
rect 114632 468450 114968 468466
rect 401100 468460 401396 468466
rect 401048 468454 401396 468460
rect 114632 468444 114980 468450
rect 114632 468438 114928 468444
rect 401060 468438 401396 468454
rect 114928 468386 114980 468392
rect 461136 468330 461164 469338
rect 464356 468602 464384 470562
rect 464356 468574 464692 468602
rect 77372 468302 77708 468318
rect 103256 468302 103408 468330
rect 423600 468314 423752 468330
rect 423588 468308 423752 468314
rect 423640 468302 423752 468308
rect 461012 468302 461164 468330
rect 423588 468250 423640 468256
rect 404728 468240 404780 468246
rect 404780 468188 405076 468194
rect 404728 468182 405076 468188
rect 404740 468166 405076 468182
rect 449452 468178 449788 468194
rect 449440 468172 449788 468178
rect 449492 468166 449788 468172
rect 449440 468114 449492 468120
rect 55128 468104 55180 468110
rect 43994 468072 44050 468081
rect 43884 468030 43994 468058
rect 47858 468072 47914 468081
rect 47564 468030 47858 468058
rect 43994 468007 44050 468016
rect 51538 468072 51594 468081
rect 51244 468030 51538 468058
rect 47858 468007 47914 468016
rect 55016 468052 55128 468058
rect 62762 468072 62818 468081
rect 55016 468046 55180 468052
rect 55016 468030 55168 468046
rect 62468 468030 62762 468058
rect 51538 468007 51594 468016
rect 73802 468072 73858 468081
rect 73600 468030 73802 468058
rect 62762 468007 62818 468016
rect 126058 468072 126114 468081
rect 125764 468030 126058 468058
rect 73802 468007 73858 468016
rect 137282 468072 137338 468081
rect 136988 468030 137282 468058
rect 126058 468007 126114 468016
rect 137282 468007 137338 468016
rect 363878 468072 363934 468081
rect 374918 468072 374974 468081
rect 363934 468030 364136 468058
rect 363878 468007 363934 468016
rect 397458 468072 397514 468081
rect 374974 468030 375268 468058
rect 374918 468007 374974 468016
rect 397514 468030 397624 468058
rect 427096 468042 427432 468058
rect 445772 468042 446108 468058
rect 427084 468036 427432 468042
rect 397458 468007 397514 468016
rect 427136 468030 427432 468036
rect 445760 468036 446108 468042
rect 427084 467978 427136 467984
rect 445812 468030 446108 468036
rect 445760 467978 445812 467984
rect 40774 466984 40830 466993
rect 40774 466919 40830 466928
rect 40788 411262 40816 466919
rect 40776 411256 40828 411262
rect 40776 411198 40828 411204
rect 467116 179382 467144 471106
rect 467208 219434 467236 471174
rect 467300 259418 467328 471242
rect 467392 365702 467420 471378
rect 497464 470892 497516 470898
rect 497464 470834 497516 470840
rect 468484 470416 468536 470422
rect 468484 470358 468536 470364
rect 468496 458182 468524 470358
rect 486424 470280 486476 470286
rect 486424 470222 486476 470228
rect 483664 470076 483716 470082
rect 483664 470018 483716 470024
rect 479524 469940 479576 469946
rect 479524 469882 479576 469888
rect 472624 469668 472676 469674
rect 472624 469610 472676 469616
rect 471244 468104 471296 468110
rect 471244 468046 471296 468052
rect 468484 458176 468536 458182
rect 468484 458118 468536 458124
rect 467380 365696 467432 365702
rect 467380 365638 467432 365644
rect 467288 259412 467340 259418
rect 467288 259354 467340 259360
rect 467196 219428 467248 219434
rect 467196 219370 467248 219376
rect 467104 179376 467156 179382
rect 467104 179318 467156 179324
rect 471256 46918 471284 468046
rect 472636 86970 472664 469610
rect 475384 468376 475436 468382
rect 475384 468318 475436 468324
rect 475396 126954 475424 468318
rect 479536 167006 479564 469882
rect 482284 468580 482336 468586
rect 482284 468522 482336 468528
rect 482296 206990 482324 468522
rect 483676 245614 483704 470018
rect 485044 468784 485096 468790
rect 485044 468726 485096 468732
rect 485056 299470 485084 468726
rect 486436 353258 486464 470222
rect 493324 469532 493376 469538
rect 493324 469474 493376 469480
rect 490564 469328 490616 469334
rect 490564 469270 490616 469276
rect 489184 468920 489236 468926
rect 489184 468862 489236 468868
rect 489196 405686 489224 468862
rect 489184 405680 489236 405686
rect 489184 405622 489236 405628
rect 486424 353252 486476 353258
rect 486424 353194 486476 353200
rect 485044 299464 485096 299470
rect 485044 299406 485096 299412
rect 483664 245608 483716 245614
rect 483664 245550 483716 245556
rect 482284 206984 482336 206990
rect 482284 206926 482336 206932
rect 479524 167000 479576 167006
rect 479524 166942 479576 166948
rect 475384 126948 475436 126954
rect 475384 126890 475436 126896
rect 472624 86964 472676 86970
rect 472624 86906 472676 86912
rect 490576 73166 490604 469270
rect 493336 113150 493364 469474
rect 497476 193186 497504 470834
rect 500224 469804 500276 469810
rect 500224 469746 500276 469752
rect 500236 233238 500264 469746
rect 501604 468444 501656 468450
rect 501604 468386 501656 468392
rect 501616 273222 501644 468386
rect 504362 467528 504418 467537
rect 504362 467463 504418 467472
rect 502982 467392 503038 467401
rect 502982 467327 503038 467336
rect 502996 325650 503024 467327
rect 504376 379506 504404 467463
rect 508502 467256 508558 467265
rect 508502 467191 508558 467200
rect 507122 467120 507178 467129
rect 507122 467055 507178 467064
rect 504364 379500 504416 379506
rect 504364 379442 504416 379448
rect 502984 325644 503036 325650
rect 502984 325586 503036 325592
rect 501604 273216 501656 273222
rect 501604 273158 501656 273164
rect 500224 233232 500276 233238
rect 500224 233174 500276 233180
rect 497464 193180 497516 193186
rect 497464 193122 497516 193128
rect 493324 113144 493376 113150
rect 493324 113086 493376 113092
rect 490564 73160 490616 73166
rect 490564 73102 490616 73108
rect 507136 60722 507164 467055
rect 508516 100706 508544 467191
rect 511276 139398 511304 471990
rect 512656 313274 512684 472058
rect 558932 471374 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 558920 471368 558972 471374
rect 558920 471310 558972 471316
rect 580184 470694 580212 471407
rect 580172 470688 580224 470694
rect 580172 470630 580224 470636
rect 580448 470212 580500 470218
rect 580448 470154 580500 470160
rect 580264 469056 580316 469062
rect 580264 468998 580316 469004
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 579620 405680 579672 405686
rect 579620 405622 579672 405628
rect 579632 404977 579660 405622
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 512644 313268 512696 313274
rect 512644 313210 512696 313216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 579896 219428 579948 219434
rect 579896 219370 579948 219376
rect 579908 219065 579936 219370
rect 579894 219056 579950 219065
rect 579894 218991 579950 219000
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 579988 179376 580040 179382
rect 579988 179318 580040 179324
rect 580000 179217 580028 179318
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580276 152697 580304 468998
rect 580356 467900 580408 467906
rect 580356 467842 580408 467848
rect 580368 418305 580396 467842
rect 580460 431633 580488 470154
rect 580446 431624 580502 431633
rect 580446 431559 580502 431568
rect 580354 418296 580410 418305
rect 580354 418231 580410 418240
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 511264 139392 511316 139398
rect 580172 139392 580224 139398
rect 511264 139334 511316 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 508504 100700 508556 100706
rect 508504 100642 508556 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 507124 60716 507176 60722
rect 507124 60658 507176 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 471244 46912 471296 46918
rect 471244 46854 471296 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 41524 42078 42412 42106
rect 40684 20664 40736 20670
rect 40684 20606 40736 20612
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 32416 480 32444 3334
rect 33600 3256 33652 3262
rect 33600 3198 33652 3204
rect 33612 480 33640 3198
rect 34808 480 34836 3334
rect 37188 3120 37240 3126
rect 37188 3062 37240 3068
rect 35992 2916 36044 2922
rect 35992 2858 36044 2864
rect 36004 480 36032 2858
rect 37200 480 37228 3062
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41524 3466 41552 42078
rect 43226 41834 43254 42092
rect 44054 41834 44082 42092
rect 44974 41834 45002 42092
rect 45802 41834 45830 42092
rect 46630 41834 46658 42092
rect 47550 41834 47578 42092
rect 48378 41834 48406 42092
rect 49206 41834 49234 42092
rect 50126 41834 50154 42092
rect 50954 41834 50982 42092
rect 51782 41834 51810 42092
rect 52702 41834 52730 42092
rect 53530 41834 53558 42092
rect 54450 41834 54478 42092
rect 55278 41834 55306 42092
rect 56106 41834 56134 42092
rect 42812 41806 43254 41834
rect 43364 41806 44082 41834
rect 44928 41806 45002 41834
rect 45664 41806 45830 41834
rect 46584 41806 46658 41834
rect 46952 41806 47578 41834
rect 48332 41806 48406 41834
rect 49160 41806 49234 41834
rect 49712 41806 50154 41834
rect 50356 41806 50982 41834
rect 51736 41806 51810 41834
rect 52656 41806 52730 41834
rect 53484 41806 53558 41834
rect 53852 41806 54478 41834
rect 55232 41806 55306 41834
rect 56060 41806 56134 41834
rect 56600 41880 56652 41886
rect 57026 41834 57054 42092
rect 57854 41886 57882 42092
rect 56600 41822 56652 41828
rect 42708 38956 42760 38962
rect 42708 38898 42760 38904
rect 42720 3534 42748 38898
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 42812 3482 42840 41806
rect 43364 26234 43392 41806
rect 44928 39370 44956 41806
rect 44916 39364 44968 39370
rect 44916 39306 44968 39312
rect 45468 39364 45520 39370
rect 45468 39306 45520 39312
rect 43444 38888 43496 38894
rect 43444 38830 43496 38836
rect 42904 26206 43392 26234
rect 42904 3670 42932 26206
rect 42892 3664 42944 3670
rect 42892 3606 42944 3612
rect 41512 3460 41564 3466
rect 41512 3402 41564 3408
rect 40684 3120 40736 3126
rect 40684 3062 40736 3068
rect 40696 480 40724 3062
rect 41892 480 41920 3470
rect 42812 3466 42932 3482
rect 42812 3460 42944 3466
rect 42812 3454 42892 3460
rect 42892 3402 42944 3408
rect 43456 3330 43484 38830
rect 44272 3460 44324 3466
rect 44272 3402 44324 3408
rect 43444 3324 43496 3330
rect 43444 3266 43496 3272
rect 43076 2848 43128 2854
rect 43076 2790 43128 2796
rect 43088 480 43116 2790
rect 44284 480 44312 3402
rect 45480 480 45508 39306
rect 45664 3602 45692 41806
rect 46584 39506 46612 41806
rect 46572 39500 46624 39506
rect 46572 39442 46624 39448
rect 46204 38684 46256 38690
rect 46204 38626 46256 38632
rect 45652 3596 45704 3602
rect 45652 3538 45704 3544
rect 46216 3058 46244 38626
rect 46952 3534 46980 41806
rect 48332 39438 48360 41806
rect 48320 39432 48372 39438
rect 48320 39374 48372 39380
rect 49160 38894 49188 41806
rect 49608 39432 49660 39438
rect 49608 39374 49660 39380
rect 49148 38888 49200 38894
rect 49148 38830 49200 38836
rect 48964 38820 49016 38826
rect 48964 38762 49016 38768
rect 48976 6914 49004 38762
rect 48884 6886 49004 6914
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 46664 3324 46716 3330
rect 46664 3266 46716 3272
rect 46204 3052 46256 3058
rect 46204 2994 46256 3000
rect 46676 480 46704 3266
rect 47860 3052 47912 3058
rect 47860 2994 47912 3000
rect 47872 480 47900 2994
rect 48884 2990 48912 6886
rect 49620 3534 49648 39374
rect 49712 3874 49740 41806
rect 50356 26234 50384 41806
rect 51736 39574 51764 41806
rect 52656 39642 52684 41806
rect 53484 39778 53512 41806
rect 53472 39772 53524 39778
rect 53472 39714 53524 39720
rect 52644 39636 52696 39642
rect 52644 39578 52696 39584
rect 53748 39636 53800 39642
rect 53748 39578 53800 39584
rect 51724 39568 51776 39574
rect 51724 39510 51776 39516
rect 53656 39500 53708 39506
rect 53656 39442 53708 39448
rect 50988 38888 51040 38894
rect 50988 38830 51040 38836
rect 49804 26206 50384 26234
rect 49700 3868 49752 3874
rect 49700 3810 49752 3816
rect 49804 3670 49832 26206
rect 49792 3664 49844 3670
rect 49792 3606 49844 3612
rect 51000 3534 51028 38830
rect 51356 3596 51408 3602
rect 51356 3538 51408 3544
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 48872 2984 48924 2990
rect 48872 2926 48924 2932
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51368 480 51396 3538
rect 53668 3534 53696 39442
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 53656 3528 53708 3534
rect 53656 3470 53708 3476
rect 52564 480 52592 3470
rect 53760 480 53788 39578
rect 53852 4010 53880 41806
rect 55232 39710 55260 41806
rect 55220 39704 55272 39710
rect 55220 39646 55272 39652
rect 55864 38752 55916 38758
rect 55864 38694 55916 38700
rect 53840 4004 53892 4010
rect 53840 3946 53892 3952
rect 54944 3664 54996 3670
rect 54944 3606 54996 3612
rect 54956 480 54984 3606
rect 55876 2922 55904 38694
rect 56060 38690 56088 41806
rect 56508 39568 56560 39574
rect 56508 39510 56560 39516
rect 56048 38684 56100 38690
rect 56048 38626 56100 38632
rect 56520 3806 56548 39510
rect 56612 3942 56640 41822
rect 56704 41806 57054 41834
rect 57842 41880 57894 41886
rect 58682 41834 58710 42092
rect 59602 41834 59630 42092
rect 60430 41834 60458 42092
rect 61258 41834 61286 42092
rect 62178 41834 62206 42092
rect 63006 41834 63034 42092
rect 63926 41834 63954 42092
rect 64754 41834 64782 42092
rect 65582 41834 65610 42092
rect 66502 41834 66530 42092
rect 67330 41834 67358 42092
rect 68158 41834 68186 42092
rect 57842 41822 57894 41828
rect 58636 41806 58710 41834
rect 59556 41806 59630 41834
rect 60384 41806 60458 41834
rect 60752 41806 61286 41834
rect 62132 41806 62206 41834
rect 62960 41806 63034 41834
rect 63604 41806 63954 41834
rect 64708 41806 64782 41834
rect 65536 41806 65610 41834
rect 66364 41806 66530 41834
rect 67284 41806 67358 41834
rect 68112 41806 68186 41834
rect 69078 41834 69106 42092
rect 69906 41834 69934 42092
rect 69078 41806 69244 41834
rect 56600 3936 56652 3942
rect 56600 3878 56652 3884
rect 56048 3800 56100 3806
rect 56048 3742 56100 3748
rect 56508 3800 56560 3806
rect 56508 3742 56560 3748
rect 55864 2916 55916 2922
rect 55864 2858 55916 2864
rect 56060 480 56088 3742
rect 56704 3738 56732 41806
rect 58636 39846 58664 41806
rect 59556 39914 59584 41806
rect 60384 40050 60412 41806
rect 60372 40044 60424 40050
rect 60372 39986 60424 39992
rect 59544 39908 59596 39914
rect 59544 39850 59596 39856
rect 58624 39840 58676 39846
rect 58624 39782 58676 39788
rect 60648 39840 60700 39846
rect 60648 39782 60700 39788
rect 57888 39704 57940 39710
rect 57888 39646 57940 39652
rect 56692 3732 56744 3738
rect 56692 3674 56744 3680
rect 57900 3398 57928 39646
rect 58440 3732 58492 3738
rect 58440 3674 58492 3680
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 57888 3392 57940 3398
rect 57888 3334 57940 3340
rect 57256 480 57284 3334
rect 58452 480 58480 3674
rect 60660 3398 60688 39782
rect 60752 4146 60780 41806
rect 62132 39982 62160 41806
rect 62120 39976 62172 39982
rect 62120 39918 62172 39924
rect 62028 39908 62080 39914
rect 62028 39850 62080 39856
rect 60740 4140 60792 4146
rect 60740 4082 60792 4088
rect 61936 3800 61988 3806
rect 61936 3742 61988 3748
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60832 3392 60884 3398
rect 60832 3334 60884 3340
rect 59648 480 59676 3334
rect 60844 480 60872 3334
rect 61948 1986 61976 3742
rect 62040 3398 62068 39850
rect 62960 38826 62988 41806
rect 63408 39772 63460 39778
rect 63408 39714 63460 39720
rect 62948 38820 63000 38826
rect 62948 38762 63000 38768
rect 62764 38684 62816 38690
rect 62764 38626 62816 38632
rect 62028 3392 62080 3398
rect 62028 3334 62080 3340
rect 62776 2854 62804 38626
rect 63420 6914 63448 39714
rect 63236 6886 63448 6914
rect 62764 2848 62816 2854
rect 62764 2790 62816 2796
rect 61948 1958 62068 1986
rect 62040 480 62068 1958
rect 63236 480 63264 6886
rect 63604 3330 63632 41806
rect 64708 39302 64736 41806
rect 64788 39976 64840 39982
rect 64788 39918 64840 39924
rect 64696 39296 64748 39302
rect 64696 39238 64748 39244
rect 64144 38820 64196 38826
rect 64144 38762 64196 38768
rect 64156 3874 64184 38762
rect 64144 3868 64196 3874
rect 64144 3810 64196 3816
rect 64800 3398 64828 39918
rect 65536 39234 65564 41806
rect 65524 39228 65576 39234
rect 65524 39170 65576 39176
rect 65524 3868 65576 3874
rect 65524 3810 65576 3816
rect 64328 3392 64380 3398
rect 64328 3334 64380 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 63592 3324 63644 3330
rect 63592 3266 63644 3272
rect 64340 480 64368 3334
rect 65536 480 65564 3810
rect 66364 3262 66392 41806
rect 67284 39098 67312 41806
rect 67548 40044 67600 40050
rect 67548 39986 67600 39992
rect 67272 39092 67324 39098
rect 67272 39034 67324 39040
rect 67560 3466 67588 39986
rect 68112 38758 68140 41806
rect 68928 39092 68980 39098
rect 68928 39034 68980 39040
rect 68100 38752 68152 38758
rect 68100 38694 68152 38700
rect 68940 3466 68968 39034
rect 69112 3936 69164 3942
rect 69112 3878 69164 3884
rect 66720 3460 66772 3466
rect 66720 3402 66772 3408
rect 67548 3460 67600 3466
rect 67548 3402 67600 3408
rect 67916 3460 67968 3466
rect 67916 3402 67968 3408
rect 68928 3460 68980 3466
rect 68928 3402 68980 3408
rect 66352 3256 66404 3262
rect 66352 3198 66404 3204
rect 66732 480 66760 3402
rect 67928 480 67956 3402
rect 69124 480 69152 3878
rect 69216 3194 69244 41806
rect 69860 41806 69934 41834
rect 70492 41880 70544 41886
rect 70734 41834 70762 42092
rect 71654 41886 71682 42092
rect 70492 41822 70544 41828
rect 69860 39166 69888 41806
rect 70308 39296 70360 39302
rect 70308 39238 70360 39244
rect 69848 39160 69900 39166
rect 69848 39102 69900 39108
rect 69204 3188 69256 3194
rect 69204 3130 69256 3136
rect 70320 480 70348 39238
rect 70504 3126 70532 41822
rect 70688 41806 70762 41834
rect 71642 41880 71694 41886
rect 72482 41834 72510 42092
rect 73310 41834 73338 42092
rect 74230 41834 74258 42092
rect 75058 41834 75086 42092
rect 75978 41834 76006 42092
rect 76806 41834 76834 42092
rect 77634 41834 77662 42092
rect 78554 41834 78582 42092
rect 79382 41834 79410 42092
rect 80210 41834 80238 42092
rect 81130 41834 81158 42092
rect 81958 41834 81986 42092
rect 71642 41822 71694 41828
rect 72436 41806 72510 41834
rect 73264 41806 73338 41834
rect 73448 41806 74258 41834
rect 75012 41806 75086 41834
rect 75932 41806 76006 41834
rect 76116 41806 76834 41834
rect 77588 41806 77662 41834
rect 78416 41806 78582 41834
rect 78692 41806 79410 41834
rect 80164 41806 80238 41834
rect 81084 41806 81158 41834
rect 81452 41806 81986 41834
rect 82786 41834 82814 42092
rect 83706 41834 83734 42092
rect 84534 41834 84562 42092
rect 85454 41834 85482 42092
rect 86282 41834 86310 42092
rect 87110 41834 87138 42092
rect 88030 41834 88058 42092
rect 88858 41834 88886 42092
rect 82786 41806 82860 41834
rect 70688 39030 70716 41806
rect 71688 39228 71740 39234
rect 71688 39170 71740 39176
rect 70676 39024 70728 39030
rect 70676 38966 70728 38972
rect 71700 6914 71728 39170
rect 72436 38962 72464 41806
rect 73068 39024 73120 39030
rect 73068 38966 73120 38972
rect 72424 38956 72476 38962
rect 72424 38898 72476 38904
rect 71516 6886 71728 6914
rect 70492 3120 70544 3126
rect 70492 3062 70544 3068
rect 71516 480 71544 6886
rect 73080 3466 73108 38966
rect 73264 38690 73292 41806
rect 73252 38684 73304 38690
rect 73252 38626 73304 38632
rect 72608 3460 72660 3466
rect 72608 3402 72660 3408
rect 73068 3460 73120 3466
rect 73068 3402 73120 3408
rect 72620 480 72648 3402
rect 73448 3398 73476 41806
rect 75012 39370 75040 41806
rect 75000 39364 75052 39370
rect 75000 39306 75052 39312
rect 75828 39364 75880 39370
rect 75828 39306 75880 39312
rect 74448 39160 74500 39166
rect 74448 39102 74500 39108
rect 74460 3466 74488 39102
rect 75840 3534 75868 39306
rect 75932 38826 75960 41806
rect 75920 38820 75972 38826
rect 75920 38762 75972 38768
rect 76116 3602 76144 41806
rect 77588 39438 77616 41806
rect 77576 39432 77628 39438
rect 77576 39374 77628 39380
rect 77208 38956 77260 38962
rect 77208 38898 77260 38904
rect 76104 3596 76156 3602
rect 76104 3538 76156 3544
rect 77220 3534 77248 38898
rect 78416 38894 78444 41806
rect 78496 39432 78548 39438
rect 78496 39374 78548 39380
rect 78404 38888 78456 38894
rect 78404 38830 78456 38836
rect 78508 3534 78536 39374
rect 78588 38820 78640 38826
rect 78588 38762 78640 38768
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 77392 3528 77444 3534
rect 77392 3470 77444 3476
rect 78496 3528 78548 3534
rect 78496 3470 78548 3476
rect 73804 3460 73856 3466
rect 73804 3402 73856 3408
rect 74448 3460 74500 3466
rect 74448 3402 74500 3408
rect 73436 3392 73488 3398
rect 73436 3334 73488 3340
rect 73816 480 73844 3402
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77404 480 77432 3470
rect 78600 480 78628 38762
rect 78692 3670 78720 41806
rect 80164 39506 80192 41806
rect 81084 39642 81112 41806
rect 81072 39636 81124 39642
rect 81072 39578 81124 39584
rect 80152 39500 80204 39506
rect 80152 39442 80204 39448
rect 81348 39500 81400 39506
rect 81348 39442 81400 39448
rect 79968 38888 80020 38894
rect 79968 38830 80020 38836
rect 79980 6914 80008 38830
rect 79704 6886 80008 6914
rect 78680 3664 78732 3670
rect 78680 3606 78732 3612
rect 79704 480 79732 6886
rect 81360 3534 81388 39442
rect 81452 4010 81480 41806
rect 82832 39574 82860 41806
rect 83660 41806 83734 41834
rect 84304 41806 84562 41834
rect 85408 41806 85482 41834
rect 86236 41806 86310 41834
rect 87064 41806 87138 41834
rect 87984 41806 88058 41834
rect 88812 41806 88886 41834
rect 89686 41834 89714 42092
rect 90606 41834 90634 42092
rect 91434 41970 91462 42092
rect 89686 41806 89760 41834
rect 83660 39710 83688 41806
rect 83648 39704 83700 39710
rect 83648 39646 83700 39652
rect 84108 39636 84160 39642
rect 84108 39578 84160 39584
rect 82820 39568 82872 39574
rect 82820 39510 82872 39516
rect 82728 38752 82780 38758
rect 82728 38694 82780 38700
rect 81440 4004 81492 4010
rect 81440 3946 81492 3952
rect 82740 3534 82768 38694
rect 84120 3534 84148 39578
rect 84304 3738 84332 41806
rect 85408 39846 85436 41806
rect 86236 39914 86264 41806
rect 86224 39908 86276 39914
rect 86224 39850 86276 39856
rect 86868 39908 86920 39914
rect 86868 39850 86920 39856
rect 85396 39840 85448 39846
rect 85396 39782 85448 39788
rect 85488 39704 85540 39710
rect 85488 39646 85540 39652
rect 84292 3732 84344 3738
rect 84292 3674 84344 3680
rect 85500 3534 85528 39646
rect 86776 39568 86828 39574
rect 86776 39510 86828 39516
rect 86788 16574 86816 39510
rect 86696 16546 86816 16574
rect 85672 3664 85724 3670
rect 85672 3606 85724 3612
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81348 3528 81400 3534
rect 81348 3470 81400 3476
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 82728 3528 82780 3534
rect 82728 3470 82780 3476
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 84108 3528 84160 3534
rect 84108 3470 84160 3476
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 80900 480 80928 3470
rect 82096 480 82124 3470
rect 83292 480 83320 3470
rect 84488 480 84516 3470
rect 85684 480 85712 3606
rect 86696 3516 86724 16546
rect 86880 6914 86908 39850
rect 86788 6886 86908 6914
rect 86788 3670 86816 6886
rect 87064 3806 87092 41806
rect 87984 39778 88012 41806
rect 88812 39982 88840 41806
rect 88800 39976 88852 39982
rect 88800 39918 88852 39924
rect 89628 39976 89680 39982
rect 89628 39918 89680 39924
rect 87972 39772 88024 39778
rect 87972 39714 88024 39720
rect 88248 39772 88300 39778
rect 88248 39714 88300 39720
rect 88260 6914 88288 39714
rect 87984 6886 88288 6914
rect 87052 3800 87104 3806
rect 87052 3742 87104 3748
rect 86776 3664 86828 3670
rect 86776 3606 86828 3612
rect 86696 3488 86908 3516
rect 86880 480 86908 3488
rect 87984 480 88012 6886
rect 89640 3534 89668 39918
rect 89732 3874 89760 41806
rect 90560 41806 90634 41834
rect 91112 41942 91462 41970
rect 90560 40050 90588 41806
rect 90548 40044 90600 40050
rect 90548 39986 90600 39992
rect 91008 39840 91060 39846
rect 91008 39782 91060 39788
rect 89720 3868 89772 3874
rect 89720 3810 89772 3816
rect 91020 3534 91048 39782
rect 91112 39098 91140 41942
rect 92262 41834 92290 42092
rect 93182 41834 93210 42092
rect 94010 41834 94038 42092
rect 94930 41834 94958 42092
rect 95758 41834 95786 42092
rect 91204 41806 92290 41834
rect 93136 41806 93210 41834
rect 93964 41806 94038 41834
rect 94884 41806 94958 41834
rect 95712 41806 95786 41834
rect 96586 41834 96614 42092
rect 97506 41834 97534 42092
rect 98334 41834 98362 42092
rect 99162 41834 99190 42092
rect 100082 41834 100110 42092
rect 100910 41834 100938 42092
rect 101738 41834 101766 42092
rect 102658 41834 102686 42092
rect 96586 41806 96660 41834
rect 91100 39092 91152 39098
rect 91100 39034 91152 39040
rect 91204 3942 91232 41806
rect 93136 39302 93164 41806
rect 93124 39296 93176 39302
rect 93124 39238 93176 39244
rect 93964 39234 93992 41806
rect 93952 39228 94004 39234
rect 93952 39170 94004 39176
rect 92388 39092 92440 39098
rect 92388 39034 92440 39040
rect 91192 3936 91244 3942
rect 91192 3878 91244 3884
rect 92400 3534 92428 39034
rect 94884 39030 94912 41806
rect 95056 40044 95108 40050
rect 95056 39986 95108 39992
rect 94872 39024 94924 39030
rect 94872 38966 94924 38972
rect 93768 38684 93820 38690
rect 93768 38626 93820 38632
rect 93780 3534 93808 38626
rect 95068 16574 95096 39986
rect 95148 39296 95200 39302
rect 95148 39238 95200 39244
rect 94976 16546 95096 16574
rect 93952 3596 94004 3602
rect 93952 3538 94004 3544
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 89628 3528 89680 3534
rect 89628 3470 89680 3476
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 92388 3528 92440 3534
rect 92388 3470 92440 3476
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 89180 480 89208 3470
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 92768 480 92796 3470
rect 93964 480 93992 3538
rect 94976 3482 95004 16546
rect 95160 6914 95188 39238
rect 95712 39166 95740 41806
rect 96632 39370 96660 41806
rect 97460 41806 97534 41834
rect 98288 41806 98362 41834
rect 99116 41806 99190 41834
rect 100036 41806 100110 41834
rect 100864 41806 100938 41834
rect 101692 41806 101766 41834
rect 102612 41806 102686 41834
rect 103486 41834 103514 42092
rect 104314 41834 104342 42092
rect 105234 41834 105262 42092
rect 106062 41834 106090 42092
rect 106982 41834 107010 42092
rect 107810 41834 107838 42092
rect 108638 41834 108666 42092
rect 109558 41834 109586 42092
rect 103486 41806 103560 41834
rect 96620 39364 96672 39370
rect 96620 39306 96672 39312
rect 96528 39228 96580 39234
rect 96528 39170 96580 39176
rect 95700 39160 95752 39166
rect 95700 39102 95752 39108
rect 96540 6914 96568 39170
rect 97460 38962 97488 41806
rect 98288 39438 98316 41806
rect 98276 39432 98328 39438
rect 98276 39374 98328 39380
rect 97908 39364 97960 39370
rect 97908 39306 97960 39312
rect 97448 38956 97500 38962
rect 97448 38898 97500 38904
rect 95068 6886 95188 6914
rect 96264 6886 96568 6914
rect 95068 3602 95096 6886
rect 95056 3596 95108 3602
rect 95056 3538 95108 3544
rect 94976 3454 95188 3482
rect 95160 480 95188 3454
rect 96264 480 96292 6886
rect 97920 3534 97948 39306
rect 99116 38826 99144 41806
rect 99288 39432 99340 39438
rect 99288 39374 99340 39380
rect 99104 38820 99156 38826
rect 99104 38762 99156 38768
rect 99300 3534 99328 39374
rect 100036 38894 100064 41806
rect 100864 39506 100892 41806
rect 100852 39500 100904 39506
rect 100852 39442 100904 39448
rect 100668 39160 100720 39166
rect 100668 39102 100720 39108
rect 100024 38888 100076 38894
rect 100024 38830 100076 38836
rect 100680 3534 100708 39102
rect 101692 38758 101720 41806
rect 102612 39642 102640 41806
rect 103532 39710 103560 41806
rect 104268 41806 104342 41834
rect 105188 41806 105262 41834
rect 106016 41806 106090 41834
rect 106936 41806 107010 41834
rect 107764 41806 107838 41834
rect 108592 41806 108666 41834
rect 109512 41806 109586 41834
rect 110386 41834 110414 42092
rect 111214 41834 111242 42092
rect 112134 41834 112162 42092
rect 112962 41834 112990 42092
rect 113790 41834 113818 42092
rect 114710 41834 114738 42092
rect 115538 41834 115566 42092
rect 116458 41834 116486 42092
rect 110386 41806 110460 41834
rect 104268 39914 104296 41806
rect 104256 39908 104308 39914
rect 104256 39850 104308 39856
rect 103520 39704 103572 39710
rect 103520 39646 103572 39652
rect 104808 39704 104860 39710
rect 104808 39646 104860 39652
rect 102600 39636 102652 39642
rect 102600 39578 102652 39584
rect 103336 39636 103388 39642
rect 103336 39578 103388 39584
rect 102048 39024 102100 39030
rect 102048 38966 102100 38972
rect 101680 38752 101732 38758
rect 101680 38694 101732 38700
rect 102060 3534 102088 38966
rect 103348 16574 103376 39578
rect 103428 39500 103480 39506
rect 103428 39442 103480 39448
rect 103256 16546 103376 16574
rect 103256 3534 103284 16546
rect 103440 6914 103468 39442
rect 104820 6914 104848 39646
rect 105188 39574 105216 41806
rect 106016 39778 106044 41806
rect 106936 39982 106964 41806
rect 106924 39976 106976 39982
rect 106924 39918 106976 39924
rect 107568 39908 107620 39914
rect 107568 39850 107620 39856
rect 106004 39772 106056 39778
rect 106004 39714 106056 39720
rect 105176 39568 105228 39574
rect 105176 39510 105228 39516
rect 106188 39568 106240 39574
rect 106188 39510 106240 39516
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 102232 3528 102284 3534
rect 102232 3470 102284 3476
rect 103244 3528 103296 3534
rect 103244 3470 103296 3476
rect 97460 480 97488 3470
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 101048 480 101076 3470
rect 102244 480 102272 3470
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 106200 3534 106228 39510
rect 107580 3534 107608 39850
rect 107764 39846 107792 41806
rect 107752 39840 107804 39846
rect 107752 39782 107804 39788
rect 108592 39098 108620 41806
rect 108948 39976 109000 39982
rect 108948 39918 109000 39924
rect 108580 39092 108632 39098
rect 108580 39034 108632 39040
rect 108960 3534 108988 39918
rect 109512 38690 109540 41806
rect 110328 39840 110380 39846
rect 110328 39782 110380 39788
rect 109500 38684 109552 38690
rect 109500 38626 109552 38632
rect 110340 3534 110368 39782
rect 110432 39302 110460 41806
rect 111168 41806 111242 41834
rect 112088 41806 112162 41834
rect 112916 41806 112990 41834
rect 113744 41806 113818 41834
rect 114664 41806 114738 41834
rect 115492 41806 115566 41834
rect 116412 41806 116486 41834
rect 117286 41834 117314 42092
rect 118114 41834 118142 42092
rect 119034 41834 119062 42092
rect 119862 41834 119890 42092
rect 120690 41834 120718 42092
rect 121610 41834 121638 42092
rect 122438 41834 122466 42092
rect 123266 41834 123294 42092
rect 117286 41806 117360 41834
rect 111168 40050 111196 41806
rect 111156 40044 111208 40050
rect 111156 39986 111208 39992
rect 111616 40044 111668 40050
rect 111616 39986 111668 39992
rect 110420 39296 110472 39302
rect 110420 39238 110472 39244
rect 111628 16574 111656 39986
rect 111708 39772 111760 39778
rect 111708 39714 111760 39720
rect 111536 16546 111656 16574
rect 111536 3534 111564 16546
rect 111720 6914 111748 39714
rect 112088 39234 112116 41806
rect 112916 39370 112944 41806
rect 113744 39438 113772 41806
rect 113732 39432 113784 39438
rect 113732 39374 113784 39380
rect 112904 39364 112956 39370
rect 112904 39306 112956 39312
rect 113088 39364 113140 39370
rect 113088 39306 113140 39312
rect 112076 39228 112128 39234
rect 112076 39170 112128 39176
rect 113100 6914 113128 39306
rect 114468 39228 114520 39234
rect 114468 39170 114520 39176
rect 111628 6886 111748 6914
rect 112824 6886 113128 6914
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 110328 3528 110380 3534
rect 110328 3470 110380 3476
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 111524 3528 111576 3534
rect 111524 3470 111576 3476
rect 105740 480 105768 3470
rect 106936 480 106964 3470
rect 108132 480 108160 3470
rect 109328 480 109356 3470
rect 110524 480 110552 3470
rect 111628 480 111656 6886
rect 112824 480 112852 6886
rect 114480 3534 114508 39170
rect 114664 39166 114692 41806
rect 114652 39160 114704 39166
rect 114652 39102 114704 39108
rect 115492 39030 115520 41806
rect 116412 39642 116440 41806
rect 116400 39636 116452 39642
rect 116400 39578 116452 39584
rect 117332 39506 117360 41806
rect 118068 41806 118142 41834
rect 118988 41806 119062 41834
rect 119816 41806 119890 41834
rect 120644 41806 120718 41834
rect 121564 41806 121638 41834
rect 122392 41806 122466 41834
rect 123220 41806 123294 41834
rect 124186 41834 124214 42092
rect 125014 41834 125042 42092
rect 125934 41834 125962 42092
rect 126762 41834 126790 42092
rect 127590 41834 127618 42092
rect 128510 41834 128538 42092
rect 129338 41834 129366 42092
rect 130166 41834 130194 42092
rect 124186 41806 124260 41834
rect 118068 39710 118096 41806
rect 118056 39704 118108 39710
rect 118056 39646 118108 39652
rect 118608 39636 118660 39642
rect 118608 39578 118660 39584
rect 117320 39500 117372 39506
rect 117320 39442 117372 39448
rect 115848 39432 115900 39438
rect 115848 39374 115900 39380
rect 115480 39024 115532 39030
rect 115480 38966 115532 38972
rect 115860 3534 115888 39374
rect 117228 39296 117280 39302
rect 117228 39238 117280 39244
rect 117240 3534 117268 39238
rect 118620 3534 118648 39578
rect 118988 39574 119016 41806
rect 119816 39914 119844 41806
rect 120644 39982 120672 41806
rect 120632 39976 120684 39982
rect 120632 39918 120684 39924
rect 119804 39908 119856 39914
rect 119804 39850 119856 39856
rect 121564 39846 121592 41806
rect 122392 40050 122420 41806
rect 122380 40044 122432 40050
rect 122380 39986 122432 39992
rect 121552 39840 121604 39846
rect 121552 39782 121604 39788
rect 122748 39840 122800 39846
rect 122748 39782 122800 39788
rect 119988 39704 120040 39710
rect 119988 39646 120040 39652
rect 118976 39568 119028 39574
rect 118976 39510 119028 39516
rect 119896 39500 119948 39506
rect 119896 39442 119948 39448
rect 114008 3528 114060 3534
rect 114008 3470 114060 3476
rect 114468 3528 114520 3534
rect 114468 3470 114520 3476
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 117228 3528 117280 3534
rect 117228 3470 117280 3476
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 118608 3528 118660 3534
rect 118608 3470 118660 3476
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 114020 480 114048 3470
rect 115216 480 115244 3470
rect 116412 480 116440 3470
rect 117608 480 117636 3470
rect 118804 480 118832 3470
rect 119908 480 119936 39442
rect 120000 3534 120028 39646
rect 121368 39568 121420 39574
rect 121368 39510 121420 39516
rect 121380 6914 121408 39510
rect 121104 6886 121408 6914
rect 119988 3528 120040 3534
rect 119988 3470 120040 3476
rect 121104 480 121132 6886
rect 122760 3534 122788 39782
rect 123220 39778 123248 41806
rect 123208 39772 123260 39778
rect 123208 39714 123260 39720
rect 124232 39370 124260 41806
rect 124968 41806 125042 41834
rect 125888 41806 125962 41834
rect 126716 41806 126790 41834
rect 127544 41806 127618 41834
rect 128464 41806 128538 41834
rect 129292 41806 129366 41834
rect 130120 41806 130194 41834
rect 131086 41834 131114 42092
rect 131914 41834 131942 42092
rect 132742 41834 132770 42092
rect 133662 41834 133690 42092
rect 134490 41834 134518 42092
rect 135318 41834 135346 42092
rect 136238 41834 136266 42092
rect 137066 41834 137094 42092
rect 131086 41806 131160 41834
rect 124220 39364 124272 39370
rect 124220 39306 124272 39312
rect 124968 39234 124996 41806
rect 125508 39772 125560 39778
rect 125508 39714 125560 39720
rect 124956 39228 125008 39234
rect 124956 39170 125008 39176
rect 124128 38684 124180 38690
rect 124128 38626 124180 38632
rect 124140 3534 124168 38626
rect 125520 3534 125548 39714
rect 125888 39438 125916 41806
rect 125876 39432 125928 39438
rect 125876 39374 125928 39380
rect 126716 39302 126744 41806
rect 126888 39908 126940 39914
rect 126888 39850 126940 39856
rect 126704 39296 126756 39302
rect 126704 39238 126756 39244
rect 126900 3534 126928 39850
rect 127544 39642 127572 41806
rect 128268 40044 128320 40050
rect 128268 39986 128320 39992
rect 127532 39636 127584 39642
rect 127532 39578 127584 39584
rect 128176 39364 128228 39370
rect 128176 39306 128228 39312
rect 122288 3528 122340 3534
rect 122288 3470 122340 3476
rect 122748 3528 122800 3534
rect 122748 3470 122800 3476
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 122300 480 122328 3470
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 126992 480 127020 3470
rect 128188 480 128216 39306
rect 128280 3534 128308 39986
rect 128464 39710 128492 41806
rect 128452 39704 128504 39710
rect 128452 39646 128504 39652
rect 129292 39506 129320 41806
rect 129648 39636 129700 39642
rect 129648 39578 129700 39584
rect 129280 39500 129332 39506
rect 129280 39442 129332 39448
rect 129660 6914 129688 39578
rect 130120 39574 130148 41806
rect 131132 39846 131160 41806
rect 131868 41806 131942 41834
rect 132696 41806 132770 41834
rect 133616 41806 133690 41834
rect 134444 41806 134518 41834
rect 135272 41806 135346 41834
rect 136192 41806 136266 41834
rect 137020 41806 137094 41834
rect 137986 41834 138014 42092
rect 138814 41834 138842 42092
rect 139642 41834 139670 42092
rect 140562 41834 140590 42092
rect 141390 41834 141418 42092
rect 142218 41834 142246 42092
rect 143138 41834 143166 42092
rect 143966 41834 143994 42092
rect 144794 41834 144822 42092
rect 145714 41834 145742 42092
rect 146542 41834 146570 42092
rect 147462 41834 147490 42092
rect 148290 41834 148318 42092
rect 149118 41834 149146 42092
rect 150038 41834 150066 42092
rect 150866 41834 150894 42092
rect 151694 41834 151722 42092
rect 152614 41834 152642 42092
rect 153442 41834 153470 42092
rect 154270 41834 154298 42092
rect 155190 41834 155218 42092
rect 156018 41834 156046 42092
rect 137986 41806 138060 41834
rect 131120 39840 131172 39846
rect 131120 39782 131172 39788
rect 130108 39568 130160 39574
rect 130108 39510 130160 39516
rect 131028 39500 131080 39506
rect 131028 39442 131080 39448
rect 129384 6886 129688 6914
rect 128268 3528 128320 3534
rect 128268 3470 128320 3476
rect 129384 480 129412 6886
rect 131040 3534 131068 39442
rect 131868 38690 131896 41806
rect 132696 39778 132724 41806
rect 133616 39914 133644 41806
rect 134444 40050 134472 41806
rect 134432 40044 134484 40050
rect 134432 39986 134484 39992
rect 133604 39908 133656 39914
rect 133604 39850 133656 39856
rect 132684 39772 132736 39778
rect 132684 39714 132736 39720
rect 132408 39568 132460 39574
rect 132408 39510 132460 39516
rect 131856 38684 131908 38690
rect 131856 38626 131908 38632
rect 130568 3528 130620 3534
rect 130568 3470 130620 3476
rect 131028 3528 131080 3534
rect 131028 3470 131080 3476
rect 130580 480 130608 3470
rect 132420 3466 132448 39510
rect 135272 39370 135300 41806
rect 136192 39642 136220 41806
rect 136180 39636 136232 39642
rect 136180 39578 136232 39584
rect 137020 39506 137048 41806
rect 137928 39908 137980 39914
rect 137928 39850 137980 39856
rect 137008 39500 137060 39506
rect 137008 39442 137060 39448
rect 135260 39364 135312 39370
rect 135260 39306 135312 39312
rect 136548 39092 136600 39098
rect 136548 39034 136600 39040
rect 133788 38888 133840 38894
rect 133788 38830 133840 38836
rect 133800 3534 133828 38830
rect 135168 38820 135220 38826
rect 135168 38762 135220 38768
rect 135180 3534 135208 38762
rect 136560 6914 136588 39034
rect 137284 38956 137336 38962
rect 137284 38898 137336 38904
rect 136468 6886 136588 6914
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 134156 3528 134208 3534
rect 134156 3470 134208 3476
rect 135168 3528 135220 3534
rect 135168 3470 135220 3476
rect 135260 3528 135312 3534
rect 135260 3470 135312 3476
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 132408 3460 132460 3466
rect 132408 3402 132460 3408
rect 131776 480 131804 3402
rect 132972 480 133000 3470
rect 134168 480 134196 3470
rect 135272 480 135300 3470
rect 136468 480 136496 6886
rect 137296 3534 137324 38898
rect 137940 6914 137968 39850
rect 138032 39574 138060 41806
rect 138768 41806 138842 41834
rect 139596 41806 139670 41834
rect 140516 41806 140590 41834
rect 141344 41806 141418 41834
rect 142172 41806 142246 41834
rect 143092 41806 143166 41834
rect 143920 41806 143994 41834
rect 144748 41806 144822 41834
rect 145668 41806 145742 41834
rect 146496 41806 146570 41834
rect 147416 41806 147490 41834
rect 148244 41806 148318 41834
rect 149072 41806 149146 41834
rect 149992 41806 150066 41834
rect 150452 41806 150894 41834
rect 151648 41806 151722 41834
rect 152568 41806 152642 41834
rect 153212 41806 153470 41834
rect 153580 41806 154298 41834
rect 155144 41806 155218 41834
rect 155972 41806 156046 41834
rect 156938 41834 156966 42092
rect 157766 41834 157794 42092
rect 158594 41834 158622 42092
rect 159514 41834 159542 42092
rect 160342 41834 160370 42092
rect 161170 41834 161198 42092
rect 162090 41834 162118 42092
rect 162918 41834 162946 42092
rect 163746 41834 163774 42092
rect 164666 41834 164694 42092
rect 165494 41834 165522 42092
rect 156938 41806 157288 41834
rect 157766 41806 157840 41834
rect 158594 41806 158668 41834
rect 159514 41806 159588 41834
rect 160342 41806 160416 41834
rect 161170 41806 161336 41834
rect 162090 41806 162164 41834
rect 162918 41806 162992 41834
rect 163746 41806 164188 41834
rect 164666 41806 164740 41834
rect 138020 39568 138072 39574
rect 138020 39510 138072 39516
rect 138768 38894 138796 41806
rect 139308 39024 139360 39030
rect 139308 38966 139360 38972
rect 138756 38888 138808 38894
rect 138756 38830 138808 38836
rect 137664 6886 137968 6914
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 137664 480 137692 6886
rect 139320 3330 139348 38966
rect 139596 38826 139624 41806
rect 140516 38962 140544 41806
rect 140688 39976 140740 39982
rect 140688 39918 140740 39924
rect 140504 38956 140556 38962
rect 140504 38898 140556 38904
rect 139584 38820 139636 38826
rect 139584 38762 139636 38768
rect 140700 3534 140728 39918
rect 141344 39098 141372 41806
rect 142068 40044 142120 40050
rect 142068 39986 142120 39992
rect 141332 39092 141384 39098
rect 141332 39034 141384 39040
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 140688 3528 140740 3534
rect 140688 3470 140740 3476
rect 138848 3324 138900 3330
rect 138848 3266 138900 3272
rect 139308 3324 139360 3330
rect 139308 3266 139360 3272
rect 138860 480 138888 3266
rect 140056 480 140084 3470
rect 142080 2990 142108 39986
rect 142172 39914 142200 41806
rect 142160 39908 142212 39914
rect 142160 39850 142212 39856
rect 143092 39030 143120 41806
rect 143920 39982 143948 41806
rect 144748 40050 144776 41806
rect 144736 40044 144788 40050
rect 144736 39986 144788 39992
rect 143908 39976 143960 39982
rect 143908 39918 143960 39924
rect 145668 39030 145696 41806
rect 143080 39024 143132 39030
rect 143080 38966 143132 38972
rect 143448 39024 143500 39030
rect 143448 38966 143500 38972
rect 145656 39024 145708 39030
rect 145656 38966 145708 38972
rect 146208 39024 146260 39030
rect 146208 38966 146260 38972
rect 143460 3534 143488 38966
rect 144828 38956 144880 38962
rect 144828 38898 144880 38904
rect 144736 38752 144788 38758
rect 144736 38694 144788 38700
rect 142436 3528 142488 3534
rect 142436 3470 142488 3476
rect 143448 3528 143500 3534
rect 143448 3470 143500 3476
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 141240 2984 141292 2990
rect 141240 2926 141292 2932
rect 142068 2984 142120 2990
rect 142068 2926 142120 2932
rect 141252 480 141280 2926
rect 142448 480 142476 3470
rect 143552 480 143580 3470
rect 144748 480 144776 38694
rect 144840 3534 144868 38898
rect 146220 6914 146248 38966
rect 146496 38962 146524 41806
rect 146484 38956 146536 38962
rect 146484 38898 146536 38904
rect 147416 38758 147444 41806
rect 148244 39030 148272 41806
rect 148232 39024 148284 39030
rect 148232 38966 148284 38972
rect 148968 39024 149020 39030
rect 148968 38966 149020 38972
rect 147588 38956 147640 38962
rect 147588 38898 147640 38904
rect 147404 38752 147456 38758
rect 147404 38694 147456 38700
rect 145944 6886 146248 6914
rect 144828 3528 144880 3534
rect 144828 3470 144880 3476
rect 145944 480 145972 6886
rect 147600 3534 147628 38898
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 147140 480 147168 3470
rect 148980 3058 149008 38966
rect 149072 38962 149100 41806
rect 149992 39030 150020 41806
rect 149980 39024 150032 39030
rect 149980 38966 150032 38972
rect 149060 38956 149112 38962
rect 149060 38898 149112 38904
rect 150452 3534 150480 41806
rect 151648 26234 151676 41806
rect 152568 39030 152596 41806
rect 151820 39024 151872 39030
rect 151820 38966 151872 38972
rect 152556 39024 152608 39030
rect 153212 38978 153240 41806
rect 152556 38966 152608 38972
rect 150544 26206 151676 26234
rect 150544 16574 150572 26206
rect 150544 16546 150664 16574
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 150440 3528 150492 3534
rect 150440 3470 150492 3476
rect 148324 3052 148376 3058
rect 148324 2994 148376 3000
rect 148968 3052 149020 3058
rect 148968 2994 149020 3000
rect 148336 480 148364 2994
rect 149532 480 149560 3470
rect 150636 480 150664 16546
rect 151832 480 151860 38966
rect 153120 38950 153240 38978
rect 153120 6914 153148 38950
rect 153580 26234 153608 41806
rect 155144 38962 155172 41806
rect 154580 38956 154632 38962
rect 154580 38898 154632 38904
rect 155132 38956 155184 38962
rect 155132 38898 155184 38904
rect 153028 6886 153148 6914
rect 153304 26206 153608 26234
rect 153028 480 153056 6886
rect 153304 3534 153332 26206
rect 154592 16574 154620 38898
rect 154592 16546 155448 16574
rect 153292 3528 153344 3534
rect 153292 3470 153344 3476
rect 154212 3528 154264 3534
rect 154212 3470 154264 3476
rect 154224 480 154252 3470
rect 155420 480 155448 16546
rect 155972 3534 156000 41806
rect 157260 3534 157288 41806
rect 157812 39030 157840 41806
rect 157800 39024 157852 39030
rect 157800 38966 157852 38972
rect 158536 39024 158588 39030
rect 158536 38966 158588 38972
rect 158548 16574 158576 38966
rect 158456 16546 158576 16574
rect 158456 3534 158484 16546
rect 158640 6914 158668 41806
rect 159560 39030 159588 41806
rect 159548 39024 159600 39030
rect 159548 38966 159600 38972
rect 160008 39024 160060 39030
rect 160008 38966 160060 38972
rect 158548 6886 158668 6914
rect 155960 3528 156012 3534
rect 155960 3470 156012 3476
rect 156604 3528 156656 3534
rect 156604 3470 156656 3476
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 157800 3528 157852 3534
rect 157800 3470 157852 3476
rect 158444 3528 158496 3534
rect 158444 3470 158496 3476
rect 156616 480 156644 3470
rect 157812 480 157840 3470
rect 158548 3466 158576 6886
rect 160020 3534 160048 38966
rect 160388 38962 160416 41806
rect 160376 38956 160428 38962
rect 160376 38898 160428 38904
rect 161308 4010 161336 41806
rect 162136 39030 162164 41806
rect 162964 39030 162992 41806
rect 162124 39024 162176 39030
rect 162124 38966 162176 38972
rect 162768 39024 162820 39030
rect 162768 38966 162820 38972
rect 162952 39024 163004 39030
rect 162952 38966 163004 38972
rect 161388 38956 161440 38962
rect 161388 38898 161440 38904
rect 161296 4004 161348 4010
rect 161296 3946 161348 3952
rect 161400 3602 161428 38898
rect 161388 3596 161440 3602
rect 161388 3538 161440 3544
rect 162492 3596 162544 3602
rect 162492 3538 162544 3544
rect 158904 3528 158956 3534
rect 158904 3470 158956 3476
rect 160008 3528 160060 3534
rect 160008 3470 160060 3476
rect 161296 3528 161348 3534
rect 161296 3470 161348 3476
rect 158536 3460 158588 3466
rect 158536 3402 158588 3408
rect 158916 480 158944 3470
rect 160100 3460 160152 3466
rect 160100 3402 160152 3408
rect 160112 480 160140 3402
rect 161308 480 161336 3470
rect 162504 480 162532 3538
rect 162780 3058 162808 38966
rect 163688 4004 163740 4010
rect 163688 3946 163740 3952
rect 162768 3052 162820 3058
rect 162768 2994 162820 3000
rect 163700 480 163728 3946
rect 164160 3534 164188 41806
rect 164712 38826 164740 41806
rect 165448 41806 165522 41834
rect 166322 41834 166350 42092
rect 167242 41834 167270 42092
rect 168070 41834 168098 42092
rect 168990 41834 169018 42092
rect 169818 41834 169846 42092
rect 170646 41834 170674 42092
rect 171566 41834 171594 42092
rect 172394 41834 172422 42092
rect 173222 41834 173250 42092
rect 174142 41834 174170 42092
rect 174970 41834 174998 42092
rect 175798 41834 175826 42092
rect 176718 41834 176746 42092
rect 177546 41834 177574 42092
rect 178466 41834 178494 42092
rect 179294 41834 179322 42092
rect 166322 41806 166396 41834
rect 167242 41806 167316 41834
rect 168070 41806 168144 41834
rect 168990 41806 169064 41834
rect 169818 41806 169892 41834
rect 170646 41806 171088 41834
rect 171566 41806 171640 41834
rect 172394 41806 172468 41834
rect 173222 41806 173296 41834
rect 174142 41806 174216 41834
rect 174970 41806 175228 41834
rect 175798 41806 175872 41834
rect 176718 41806 176792 41834
rect 177546 41806 177988 41834
rect 178466 41806 178540 41834
rect 164700 38820 164752 38826
rect 164700 38762 164752 38768
rect 165448 3602 165476 41806
rect 166368 39030 166396 41806
rect 167288 39030 167316 41806
rect 165712 39024 165764 39030
rect 165712 38966 165764 38972
rect 166356 39024 166408 39030
rect 166356 38966 166408 38972
rect 166908 39024 166960 39030
rect 166908 38966 166960 38972
rect 167276 39024 167328 39030
rect 167276 38966 167328 38972
rect 165528 38820 165580 38826
rect 165528 38762 165580 38768
rect 165436 3596 165488 3602
rect 165436 3538 165488 3544
rect 164148 3528 164200 3534
rect 164148 3470 164200 3476
rect 165540 3194 165568 38762
rect 165724 16574 165752 38966
rect 165724 16546 166120 16574
rect 165528 3188 165580 3194
rect 165528 3130 165580 3136
rect 164884 3052 164936 3058
rect 164884 2994 164936 3000
rect 164896 480 164924 2994
rect 166092 480 166120 16546
rect 166920 3466 166948 38966
rect 168116 38826 168144 41806
rect 169036 39030 169064 41806
rect 169864 39030 169892 41806
rect 168288 39024 168340 39030
rect 168288 38966 168340 38972
rect 169024 39024 169076 39030
rect 169024 38966 169076 38972
rect 169668 39024 169720 39030
rect 169668 38966 169720 38972
rect 169852 39024 169904 39030
rect 169852 38966 169904 38972
rect 170956 39024 171008 39030
rect 170956 38966 171008 38972
rect 168104 38820 168156 38826
rect 168104 38762 168156 38768
rect 168300 4146 168328 38966
rect 169024 38820 169076 38826
rect 169024 38762 169076 38768
rect 168288 4140 168340 4146
rect 168288 4082 168340 4088
rect 169036 4010 169064 38762
rect 169024 4004 169076 4010
rect 169024 3946 169076 3952
rect 169576 3596 169628 3602
rect 169576 3538 169628 3544
rect 167184 3528 167236 3534
rect 167184 3470 167236 3476
rect 166908 3460 166960 3466
rect 166908 3402 166960 3408
rect 167196 480 167224 3470
rect 168380 3188 168432 3194
rect 168380 3130 168432 3136
rect 168392 480 168420 3130
rect 169588 480 169616 3538
rect 169680 3534 169708 38966
rect 170968 3670 170996 38966
rect 170956 3664 171008 3670
rect 170956 3606 171008 3612
rect 169668 3528 169720 3534
rect 169668 3470 169720 3476
rect 171060 3466 171088 41806
rect 171612 39030 171640 41806
rect 171600 39024 171652 39030
rect 171600 38966 171652 38972
rect 172336 39024 172388 39030
rect 172336 38966 172388 38972
rect 171968 4140 172020 4146
rect 171968 4082 172020 4088
rect 170772 3460 170824 3466
rect 170772 3402 170824 3408
rect 171048 3460 171100 3466
rect 171048 3402 171100 3408
rect 170784 480 170812 3402
rect 171980 480 172008 4082
rect 172348 3602 172376 38966
rect 172336 3596 172388 3602
rect 172336 3538 172388 3544
rect 172440 3262 172468 41806
rect 173268 39030 173296 41806
rect 173256 39024 173308 39030
rect 173256 38966 173308 38972
rect 173808 39024 173860 39030
rect 173808 38966 173860 38972
rect 173164 4004 173216 4010
rect 173164 3946 173216 3952
rect 172428 3256 172480 3262
rect 172428 3198 172480 3204
rect 173176 480 173204 3946
rect 173820 3398 173848 38966
rect 174188 38826 174216 41806
rect 174176 38820 174228 38826
rect 174176 38762 174228 38768
rect 175096 38820 175148 38826
rect 175096 38762 175148 38768
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 173808 3392 173860 3398
rect 173808 3334 173860 3340
rect 174280 480 174308 3470
rect 175108 3194 175136 38762
rect 175096 3188 175148 3194
rect 175096 3130 175148 3136
rect 175200 2990 175228 41806
rect 175844 39030 175872 41806
rect 175832 39024 175884 39030
rect 175832 38966 175884 38972
rect 176568 39024 176620 39030
rect 176568 38966 176620 38972
rect 176580 3670 176608 38966
rect 176764 38962 176792 41806
rect 176752 38956 176804 38962
rect 176752 38898 176804 38904
rect 177856 38956 177908 38962
rect 177856 38898 177908 38904
rect 177868 6914 177896 38898
rect 177776 6886 177896 6914
rect 175464 3664 175516 3670
rect 175464 3606 175516 3612
rect 176568 3664 176620 3670
rect 176568 3606 176620 3612
rect 175188 2984 175240 2990
rect 175188 2926 175240 2932
rect 175476 480 175504 3606
rect 177776 3466 177804 6886
rect 177960 3942 177988 41806
rect 178512 39030 178540 41806
rect 179248 41806 179322 41834
rect 180122 41834 180150 42092
rect 181042 41834 181070 42092
rect 181870 41834 181898 42092
rect 182698 41834 182726 42092
rect 183618 41834 183646 42092
rect 184446 41834 184474 42092
rect 185274 41834 185302 42092
rect 186194 41834 186222 42092
rect 187022 41834 187050 42092
rect 187942 41834 187970 42092
rect 188770 41834 188798 42092
rect 189598 41834 189626 42092
rect 190518 41834 190546 42092
rect 191346 41834 191374 42092
rect 192174 41834 192202 42092
rect 193094 41834 193122 42092
rect 180122 41806 180196 41834
rect 181042 41806 181116 41834
rect 181870 41806 182036 41834
rect 182698 41806 182772 41834
rect 183618 41806 183692 41834
rect 184446 41806 184796 41834
rect 185274 41806 185348 41834
rect 186194 41806 186268 41834
rect 187022 41806 187096 41834
rect 187942 41806 188016 41834
rect 188770 41806 189028 41834
rect 189598 41806 189672 41834
rect 190518 41806 190592 41834
rect 191346 41806 191788 41834
rect 192174 41806 192248 41834
rect 178500 39024 178552 39030
rect 178500 38966 178552 38972
rect 177948 3936 178000 3942
rect 177948 3878 178000 3884
rect 179248 3738 179276 41806
rect 180168 39030 180196 41806
rect 181088 39030 181116 41806
rect 179328 39024 179380 39030
rect 179328 38966 179380 38972
rect 180156 39024 180208 39030
rect 180156 38966 180208 38972
rect 180708 39024 180760 39030
rect 180708 38966 180760 38972
rect 181076 39024 181128 39030
rect 181076 38966 181128 38972
rect 179340 4010 179368 38966
rect 179328 4004 179380 4010
rect 179328 3946 179380 3952
rect 180720 3874 180748 38966
rect 180708 3868 180760 3874
rect 180708 3810 180760 3816
rect 179236 3732 179288 3738
rect 179236 3674 179288 3680
rect 182008 3602 182036 41806
rect 182744 39030 182772 41806
rect 183664 39030 183692 41806
rect 182088 39024 182140 39030
rect 182088 38966 182140 38972
rect 182732 39024 182784 39030
rect 182732 38966 182784 38972
rect 183468 39024 183520 39030
rect 183468 38966 183520 38972
rect 183652 39024 183704 39030
rect 183652 38966 183704 38972
rect 182100 4078 182128 38966
rect 182088 4072 182140 4078
rect 182088 4014 182140 4020
rect 183480 3806 183508 38966
rect 183468 3800 183520 3806
rect 183468 3742 183520 3748
rect 184768 3670 184796 41806
rect 185320 39030 185348 41806
rect 184848 39024 184900 39030
rect 184848 38966 184900 38972
rect 185308 39024 185360 39030
rect 185308 38966 185360 38972
rect 186136 39024 186188 39030
rect 186136 38966 186188 38972
rect 183744 3664 183796 3670
rect 183744 3606 183796 3612
rect 184756 3664 184808 3670
rect 184756 3606 184808 3612
rect 177856 3596 177908 3602
rect 177856 3538 177908 3544
rect 181996 3596 182048 3602
rect 181996 3538 182048 3544
rect 176660 3460 176712 3466
rect 176660 3402 176712 3408
rect 177764 3460 177816 3466
rect 177764 3402 177816 3408
rect 176672 480 176700 3402
rect 177868 480 177896 3538
rect 180248 3392 180300 3398
rect 180248 3334 180300 3340
rect 179052 3256 179104 3262
rect 179052 3198 179104 3204
rect 179064 480 179092 3198
rect 180260 480 180288 3334
rect 181444 3188 181496 3194
rect 181444 3130 181496 3136
rect 181456 480 181484 3130
rect 182548 2984 182600 2990
rect 182548 2926 182600 2932
rect 182560 480 182588 2926
rect 183756 480 183784 3606
rect 184860 3398 184888 38966
rect 186148 4146 186176 38966
rect 186136 4140 186188 4146
rect 186136 4082 186188 4088
rect 186136 3936 186188 3942
rect 186136 3878 186188 3884
rect 184940 3460 184992 3466
rect 184940 3402 184992 3408
rect 184848 3392 184900 3398
rect 184848 3334 184900 3340
rect 184952 480 184980 3402
rect 186148 480 186176 3878
rect 186240 3466 186268 41806
rect 187068 39030 187096 41806
rect 187988 39030 188016 41806
rect 187056 39024 187108 39030
rect 187056 38966 187108 38972
rect 187608 39024 187660 39030
rect 187608 38966 187660 38972
rect 187976 39024 188028 39030
rect 187976 38966 188028 38972
rect 188896 39024 188948 39030
rect 188896 38966 188948 38972
rect 187332 4004 187384 4010
rect 187332 3946 187384 3952
rect 186228 3460 186280 3466
rect 186228 3402 186280 3408
rect 187344 480 187372 3946
rect 187620 3534 187648 38966
rect 188908 3942 188936 38966
rect 188896 3936 188948 3942
rect 188896 3878 188948 3884
rect 189000 3738 189028 41806
rect 189644 39030 189672 41806
rect 190564 39030 190592 41806
rect 189632 39024 189684 39030
rect 189632 38966 189684 38972
rect 190368 39024 190420 39030
rect 190368 38966 190420 38972
rect 190552 39024 190604 39030
rect 190552 38966 190604 38972
rect 191656 39024 191708 39030
rect 191656 38966 191708 38972
rect 190380 4010 190408 38966
rect 191668 4078 191696 38966
rect 190828 4072 190880 4078
rect 190828 4014 190880 4020
rect 191656 4072 191708 4078
rect 191656 4014 191708 4020
rect 190368 4004 190420 4010
rect 190368 3946 190420 3952
rect 189724 3868 189776 3874
rect 189724 3810 189776 3816
rect 188528 3732 188580 3738
rect 188528 3674 188580 3680
rect 188988 3732 189040 3738
rect 188988 3674 189040 3680
rect 187608 3528 187660 3534
rect 187608 3470 187660 3476
rect 188540 480 188568 3674
rect 189736 480 189764 3810
rect 190840 480 190868 4014
rect 191760 3874 191788 41806
rect 192220 39030 192248 41806
rect 193048 41806 193122 41834
rect 193922 41834 193950 42092
rect 194750 41834 194778 42092
rect 195670 41834 195698 42092
rect 196498 41834 196526 42092
rect 197326 41834 197354 42092
rect 198246 41834 198274 42092
rect 199074 41834 199102 42092
rect 199994 41834 200022 42092
rect 193922 41806 193996 41834
rect 194750 41806 194824 41834
rect 195670 41806 195928 41834
rect 196498 41806 196572 41834
rect 197326 41806 197400 41834
rect 198246 41806 198596 41834
rect 199074 41806 199148 41834
rect 192208 39024 192260 39030
rect 192208 38966 192260 38972
rect 191748 3868 191800 3874
rect 191748 3810 191800 3816
rect 193048 3602 193076 41806
rect 193968 39030 193996 41806
rect 194796 39030 194824 41806
rect 193128 39024 193180 39030
rect 193128 38966 193180 38972
rect 193956 39024 194008 39030
rect 193956 38966 194008 38972
rect 194508 39024 194560 39030
rect 194508 38966 194560 38972
rect 194784 39024 194836 39030
rect 194784 38966 194836 38972
rect 195796 39024 195848 39030
rect 195796 38966 195848 38972
rect 192024 3596 192076 3602
rect 192024 3538 192076 3544
rect 193036 3596 193088 3602
rect 193036 3538 193088 3544
rect 192036 480 192064 3538
rect 193140 3126 193168 38966
rect 194520 3806 194548 38966
rect 193220 3800 193272 3806
rect 193220 3742 193272 3748
rect 194508 3800 194560 3806
rect 194508 3742 194560 3748
rect 193128 3120 193180 3126
rect 193128 3062 193180 3068
rect 193232 480 193260 3742
rect 195808 3670 195836 38966
rect 195612 3664 195664 3670
rect 195612 3606 195664 3612
rect 195796 3664 195848 3670
rect 195796 3606 195848 3612
rect 194416 3392 194468 3398
rect 194416 3334 194468 3340
rect 194428 480 194456 3334
rect 195624 480 195652 3606
rect 195900 3262 195928 41806
rect 196544 39030 196572 41806
rect 197372 39030 197400 41806
rect 196532 39024 196584 39030
rect 196532 38966 196584 38972
rect 197268 39024 197320 39030
rect 197268 38966 197320 38972
rect 197360 39024 197412 39030
rect 197360 38966 197412 38972
rect 196808 4140 196860 4146
rect 196808 4082 196860 4088
rect 195888 3256 195940 3262
rect 195888 3198 195940 3204
rect 196820 480 196848 4082
rect 197280 3194 197308 38966
rect 198568 3466 198596 41806
rect 199120 39030 199148 41806
rect 199948 41806 200022 41834
rect 200822 41834 200850 42092
rect 201650 41834 201678 42092
rect 202570 41834 202598 42092
rect 203398 41834 203426 42092
rect 204226 41834 204254 42092
rect 205146 41834 205174 42092
rect 205974 41834 206002 42092
rect 206802 41834 206830 42092
rect 207722 41834 207750 42092
rect 208550 41834 208578 42092
rect 209470 41834 209498 42092
rect 210298 41834 210326 42092
rect 211126 41834 211154 42092
rect 212046 41834 212074 42092
rect 212874 41834 212902 42092
rect 213702 41834 213730 42092
rect 214622 41834 214650 42092
rect 215450 41834 215478 42092
rect 216278 41834 216306 42092
rect 217198 41834 217226 42092
rect 218026 41834 218054 42092
rect 218946 41834 218974 42092
rect 219774 41834 219802 42092
rect 220602 41834 220630 42092
rect 221522 41834 221550 42092
rect 222350 41834 222378 42092
rect 223178 41834 223206 42092
rect 224098 41834 224126 42092
rect 224926 41834 224954 42092
rect 225754 41834 225782 42092
rect 226674 41834 226702 42092
rect 227502 41834 227530 42092
rect 228330 41834 228358 42092
rect 229250 41834 229278 42092
rect 230078 41834 230106 42092
rect 230998 41834 231026 42092
rect 231826 41834 231854 42092
rect 232654 41834 232682 42092
rect 233574 41834 233602 42092
rect 234402 41834 234430 42092
rect 235230 41834 235258 42092
rect 236150 41834 236178 42092
rect 236978 41834 237006 42092
rect 237806 41834 237834 42092
rect 238726 41834 238754 42092
rect 239554 41834 239582 42092
rect 240474 41834 240502 42092
rect 241302 41834 241330 42092
rect 242130 41834 242158 42092
rect 243050 41834 243078 42092
rect 243878 41834 243906 42092
rect 244706 41834 244734 42092
rect 245626 41834 245654 42092
rect 246454 41834 246482 42092
rect 247282 41834 247310 42092
rect 248202 41834 248230 42092
rect 249030 41834 249058 42092
rect 249950 41834 249978 42092
rect 250778 41834 250806 42092
rect 251606 41834 251634 42092
rect 252526 41834 252554 42092
rect 253354 41834 253382 42092
rect 254182 41834 254210 42092
rect 255102 41834 255130 42092
rect 255930 41834 255958 42092
rect 256758 41834 256786 42092
rect 257678 41834 257706 42092
rect 258506 41834 258534 42092
rect 259334 41834 259362 42092
rect 260254 41834 260282 42092
rect 261082 41834 261110 42092
rect 262002 41834 262030 42092
rect 262830 41834 262858 42092
rect 200822 41806 200896 41834
rect 201650 41806 201724 41834
rect 202570 41806 202736 41834
rect 203398 41806 203472 41834
rect 204226 41806 204300 41834
rect 205146 41806 205588 41834
rect 205974 41806 206048 41834
rect 206802 41806 206968 41834
rect 207722 41806 207796 41834
rect 208550 41806 208624 41834
rect 209470 41806 209728 41834
rect 210298 41806 210372 41834
rect 211126 41806 211200 41834
rect 212046 41806 212488 41834
rect 212874 41806 212948 41834
rect 213702 41806 213776 41834
rect 214622 41806 214696 41834
rect 215450 41806 215524 41834
rect 216278 41806 216352 41834
rect 217198 41806 217272 41834
rect 218026 41806 218100 41834
rect 218946 41806 219020 41834
rect 219774 41806 219848 41834
rect 220602 41806 220676 41834
rect 221522 41806 221596 41834
rect 222350 41806 222424 41834
rect 223178 41806 223436 41834
rect 224098 41806 224172 41834
rect 224926 41806 225000 41834
rect 225754 41806 226196 41834
rect 226674 41806 226748 41834
rect 227502 41806 227668 41834
rect 228330 41806 228404 41834
rect 229250 41806 229324 41834
rect 230078 41806 230428 41834
rect 230998 41806 231072 41834
rect 231826 41806 231900 41834
rect 232654 41806 232728 41834
rect 233574 41806 233648 41834
rect 234402 41806 234476 41834
rect 235230 41806 235304 41834
rect 236150 41806 236224 41834
rect 236978 41806 237052 41834
rect 237806 41806 237880 41834
rect 238726 41806 238800 41834
rect 239554 41806 239628 41834
rect 240474 41806 240548 41834
rect 241302 41806 241376 41834
rect 242130 41806 242204 41834
rect 243050 41806 243124 41834
rect 243878 41806 244136 41834
rect 244706 41806 244780 41834
rect 245626 41806 245700 41834
rect 246454 41806 246528 41834
rect 247282 41806 247356 41834
rect 248202 41806 248368 41834
rect 249030 41806 249104 41834
rect 249950 41806 250024 41834
rect 250778 41806 251128 41834
rect 251606 41806 251680 41834
rect 252526 41806 252600 41834
rect 253354 41806 253428 41834
rect 254182 41806 254256 41834
rect 255102 41806 255176 41834
rect 255930 41806 256004 41834
rect 256758 41806 256832 41834
rect 257678 41806 257752 41834
rect 258506 41806 258580 41834
rect 259334 41806 259408 41834
rect 260254 41806 260328 41834
rect 261082 41806 261156 41834
rect 262002 41806 262168 41834
rect 198648 39024 198700 39030
rect 198648 38966 198700 38972
rect 199108 39024 199160 39030
rect 199108 38966 199160 38972
rect 197912 3460 197964 3466
rect 197912 3402 197964 3408
rect 198556 3460 198608 3466
rect 198556 3402 198608 3408
rect 197268 3188 197320 3194
rect 197268 3130 197320 3136
rect 197924 480 197952 3402
rect 198660 2854 198688 38966
rect 199948 3534 199976 41806
rect 200868 39030 200896 41806
rect 201696 39030 201724 41806
rect 200028 39024 200080 39030
rect 200028 38966 200080 38972
rect 200856 39024 200908 39030
rect 200856 38966 200908 38972
rect 201408 39024 201460 39030
rect 201408 38966 201460 38972
rect 201684 39024 201736 39030
rect 201684 38966 201736 38972
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 199936 3528 199988 3534
rect 199936 3470 199988 3476
rect 198648 2848 198700 2854
rect 198648 2790 198700 2796
rect 199120 480 199148 3470
rect 200040 3330 200068 38966
rect 200304 3936 200356 3942
rect 200304 3878 200356 3884
rect 200028 3324 200080 3330
rect 200028 3266 200080 3272
rect 200316 480 200344 3878
rect 201420 3398 201448 38966
rect 202708 4010 202736 41806
rect 203444 39030 203472 41806
rect 202788 39024 202840 39030
rect 202788 38966 202840 38972
rect 203432 39024 203484 39030
rect 203432 38966 203484 38972
rect 204168 39024 204220 39030
rect 204168 38966 204220 38972
rect 202604 4004 202656 4010
rect 202604 3946 202656 3952
rect 202696 4004 202748 4010
rect 202696 3946 202748 3952
rect 201500 3732 201552 3738
rect 201500 3674 201552 3680
rect 201408 3392 201460 3398
rect 201408 3334 201460 3340
rect 201512 480 201540 3674
rect 202616 1986 202644 3946
rect 202800 2922 202828 38966
rect 204180 4146 204208 38966
rect 204272 38826 204300 41806
rect 204260 38820 204312 38826
rect 204260 38762 204312 38768
rect 205456 38820 205508 38826
rect 205456 38762 205508 38768
rect 204168 4140 204220 4146
rect 204168 4082 204220 4088
rect 203892 4072 203944 4078
rect 203892 4014 203944 4020
rect 202788 2916 202840 2922
rect 202788 2858 202840 2864
rect 202616 1958 202736 1986
rect 202708 480 202736 1958
rect 203904 480 203932 4014
rect 205468 3942 205496 38762
rect 205560 4078 205588 41806
rect 206020 39030 206048 41806
rect 206008 39024 206060 39030
rect 206008 38966 206060 38972
rect 206836 39024 206888 39030
rect 206836 38966 206888 38972
rect 205548 4072 205600 4078
rect 205548 4014 205600 4020
rect 205456 3936 205508 3942
rect 205456 3878 205508 3884
rect 206848 3874 206876 38966
rect 205088 3868 205140 3874
rect 205088 3810 205140 3816
rect 206836 3868 206888 3874
rect 206836 3810 206888 3816
rect 205100 480 205128 3810
rect 206940 3738 206968 41806
rect 207768 39030 207796 41806
rect 208596 39030 208624 41806
rect 207756 39024 207808 39030
rect 207756 38966 207808 38972
rect 208308 39024 208360 39030
rect 208308 38966 208360 38972
rect 208584 39024 208636 39030
rect 208584 38966 208636 38972
rect 209596 39024 209648 39030
rect 209596 38966 209648 38972
rect 206928 3732 206980 3738
rect 206928 3674 206980 3680
rect 207388 3596 207440 3602
rect 207388 3538 207440 3544
rect 206192 3120 206244 3126
rect 206192 3062 206244 3068
rect 206204 480 206232 3062
rect 207400 480 207428 3538
rect 208320 2990 208348 38966
rect 208584 3800 208636 3806
rect 208584 3742 208636 3748
rect 208308 2984 208360 2990
rect 208308 2926 208360 2932
rect 208596 480 208624 3742
rect 209608 3058 209636 38966
rect 209700 3126 209728 41806
rect 210344 39030 210372 41806
rect 211172 39030 211200 41806
rect 210332 39024 210384 39030
rect 210332 38966 210384 38972
rect 211068 39024 211120 39030
rect 211068 38966 211120 38972
rect 211160 39024 211212 39030
rect 211160 38966 211212 38972
rect 212356 39024 212408 39030
rect 212356 38966 212408 38972
rect 211080 3806 211108 38966
rect 211068 3800 211120 3806
rect 211068 3742 211120 3748
rect 212368 3670 212396 38966
rect 209780 3664 209832 3670
rect 209780 3606 209832 3612
rect 212356 3664 212408 3670
rect 212356 3606 212408 3612
rect 209688 3120 209740 3126
rect 209688 3062 209740 3068
rect 209596 3052 209648 3058
rect 209596 2994 209648 3000
rect 209792 480 209820 3606
rect 212460 3602 212488 41806
rect 212920 39030 212948 41806
rect 212908 39024 212960 39030
rect 212908 38966 212960 38972
rect 213748 4894 213776 41806
rect 214668 39030 214696 41806
rect 215496 39030 215524 41806
rect 216324 39370 216352 41806
rect 216312 39364 216364 39370
rect 216312 39306 216364 39312
rect 217244 39030 217272 41806
rect 218072 39030 218100 41806
rect 218992 39506 219020 41806
rect 218980 39500 219032 39506
rect 218980 39442 219032 39448
rect 219820 39030 219848 41806
rect 213828 39024 213880 39030
rect 213828 38966 213880 38972
rect 214656 39024 214708 39030
rect 214656 38966 214708 38972
rect 215208 39024 215260 39030
rect 215208 38966 215260 38972
rect 215484 39024 215536 39030
rect 215484 38966 215536 38972
rect 216588 39024 216640 39030
rect 216588 38966 216640 38972
rect 217232 39024 217284 39030
rect 217232 38966 217284 38972
rect 217968 39024 218020 39030
rect 217968 38966 218020 38972
rect 218060 39024 218112 39030
rect 218060 38966 218112 38972
rect 219348 39024 219400 39030
rect 219348 38966 219400 38972
rect 219808 39024 219860 39030
rect 219808 38966 219860 38972
rect 213736 4888 213788 4894
rect 213736 4830 213788 4836
rect 212448 3596 212500 3602
rect 212448 3538 212500 3544
rect 210976 3256 211028 3262
rect 210976 3198 211028 3204
rect 210988 480 211016 3198
rect 213840 3194 213868 38966
rect 215220 3466 215248 38966
rect 214472 3460 214524 3466
rect 214472 3402 214524 3408
rect 215208 3460 215260 3466
rect 215208 3402 215260 3408
rect 212172 3188 212224 3194
rect 212172 3130 212224 3136
rect 213828 3188 213880 3194
rect 213828 3130 213880 3136
rect 212184 480 212212 3130
rect 213368 2848 213420 2854
rect 213368 2790 213420 2796
rect 213380 480 213408 2790
rect 214484 480 214512 3402
rect 215668 3324 215720 3330
rect 215668 3266 215720 3272
rect 215680 480 215708 3266
rect 216600 3262 216628 38966
rect 217980 3534 218008 38966
rect 216864 3528 216916 3534
rect 216864 3470 216916 3476
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 216588 3256 216640 3262
rect 216588 3198 216640 3204
rect 216876 480 216904 3470
rect 219360 3398 219388 38966
rect 220648 4010 220676 41806
rect 220728 39024 220780 39030
rect 220728 38966 220780 38972
rect 220452 4004 220504 4010
rect 220452 3946 220504 3952
rect 220636 4004 220688 4010
rect 220636 3946 220688 3952
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 219348 3392 219400 3398
rect 219348 3334 219400 3340
rect 218072 480 218100 3334
rect 219256 2916 219308 2922
rect 219256 2858 219308 2864
rect 219268 480 219296 2858
rect 220464 480 220492 3946
rect 220740 3330 220768 38966
rect 221568 38826 221596 41806
rect 222396 38962 222424 41806
rect 222384 38956 222436 38962
rect 222384 38898 222436 38904
rect 221556 38820 221608 38826
rect 221556 38762 221608 38768
rect 221556 4140 221608 4146
rect 221556 4082 221608 4088
rect 220728 3324 220780 3330
rect 220728 3266 220780 3272
rect 221568 480 221596 4082
rect 223408 3942 223436 41806
rect 224144 39574 224172 41806
rect 224132 39568 224184 39574
rect 224132 39510 224184 39516
rect 224224 39500 224276 39506
rect 224224 39442 224276 39448
rect 223488 38956 223540 38962
rect 223488 38898 223540 38904
rect 223500 4146 223528 38898
rect 224236 4962 224264 39442
rect 224972 39030 225000 41806
rect 224960 39024 225012 39030
rect 224960 38966 225012 38972
rect 224224 4956 224276 4962
rect 224224 4898 224276 4904
rect 223488 4140 223540 4146
rect 223488 4082 223540 4088
rect 226168 4078 226196 41806
rect 226720 39030 226748 41806
rect 226248 39024 226300 39030
rect 226248 38966 226300 38972
rect 226708 39024 226760 39030
rect 226708 38966 226760 38972
rect 227536 39024 227588 39030
rect 227536 38966 227588 38972
rect 223948 4072 224000 4078
rect 223948 4014 224000 4020
rect 226156 4072 226208 4078
rect 226156 4014 226208 4020
rect 222752 3936 222804 3942
rect 222752 3878 222804 3884
rect 223396 3936 223448 3942
rect 223396 3878 223448 3884
rect 222764 480 222792 3878
rect 223960 480 223988 4014
rect 225144 3868 225196 3874
rect 225144 3810 225196 3816
rect 225156 480 225184 3810
rect 226260 2854 226288 38966
rect 227548 4826 227576 38966
rect 227536 4820 227588 4826
rect 227536 4762 227588 4768
rect 227640 3874 227668 41806
rect 228376 39030 228404 41806
rect 229296 39438 229324 41806
rect 229284 39432 229336 39438
rect 229284 39374 229336 39380
rect 228364 39024 228416 39030
rect 228364 38966 228416 38972
rect 229008 39024 229060 39030
rect 229008 38966 229060 38972
rect 228364 38820 228416 38826
rect 228364 38762 228416 38768
rect 228376 7614 228404 38762
rect 228364 7608 228416 7614
rect 228364 7550 228416 7556
rect 227628 3868 227680 3874
rect 227628 3810 227680 3816
rect 226340 3732 226392 3738
rect 226340 3674 226392 3680
rect 226248 2848 226300 2854
rect 226248 2790 226300 2796
rect 226352 480 226380 3674
rect 228732 3052 228784 3058
rect 228732 2994 228784 3000
rect 227536 2984 227588 2990
rect 227536 2926 227588 2932
rect 227548 480 227576 2926
rect 228744 480 228772 2994
rect 229020 2922 229048 38966
rect 230400 3738 230428 41806
rect 231044 39030 231072 41806
rect 231032 39024 231084 39030
rect 231032 38966 231084 38972
rect 231768 39024 231820 39030
rect 231768 38966 231820 38972
rect 231780 3806 231808 38966
rect 231872 38962 231900 41806
rect 232700 39030 232728 41806
rect 232688 39024 232740 39030
rect 232688 38966 232740 38972
rect 233148 39024 233200 39030
rect 233148 38966 233200 38972
rect 231860 38956 231912 38962
rect 231860 38898 231912 38904
rect 233056 38956 233108 38962
rect 233056 38898 233108 38904
rect 233068 10334 233096 38898
rect 233056 10328 233108 10334
rect 233056 10270 233108 10276
rect 231032 3800 231084 3806
rect 231032 3742 231084 3748
rect 231768 3800 231820 3806
rect 231768 3742 231820 3748
rect 230388 3732 230440 3738
rect 230388 3674 230440 3680
rect 229836 3120 229888 3126
rect 229836 3062 229888 3068
rect 229008 2916 229060 2922
rect 229008 2858 229060 2864
rect 229848 480 229876 3062
rect 231044 480 231072 3742
rect 232228 3664 232280 3670
rect 232228 3606 232280 3612
rect 232240 480 232268 3606
rect 233160 2990 233188 38966
rect 233620 38826 233648 41806
rect 233608 38820 233660 38826
rect 233608 38762 233660 38768
rect 234448 5030 234476 41806
rect 235276 39030 235304 41806
rect 236196 39030 236224 41806
rect 237024 39506 237052 41806
rect 237012 39500 237064 39506
rect 237012 39442 237064 39448
rect 237852 39030 237880 41806
rect 238024 39364 238076 39370
rect 238024 39306 238076 39312
rect 235264 39024 235316 39030
rect 235264 38966 235316 38972
rect 235908 39024 235960 39030
rect 235908 38966 235960 38972
rect 236184 39024 236236 39030
rect 236184 38966 236236 38972
rect 237288 39024 237340 39030
rect 237288 38966 237340 38972
rect 237840 39024 237892 39030
rect 237840 38966 237892 38972
rect 234528 38820 234580 38826
rect 234528 38762 234580 38768
rect 234436 5024 234488 5030
rect 234436 4966 234488 4972
rect 234540 3670 234568 38762
rect 235816 4888 235868 4894
rect 235816 4830 235868 4836
rect 234528 3664 234580 3670
rect 234528 3606 234580 3612
rect 233424 3596 233476 3602
rect 233424 3538 233476 3544
rect 233148 2984 233200 2990
rect 233148 2926 233200 2932
rect 233436 480 233464 3538
rect 234620 3188 234672 3194
rect 234620 3130 234672 3136
rect 234632 480 234660 3130
rect 235828 480 235856 4830
rect 235920 3126 235948 38966
rect 237012 3460 237064 3466
rect 237012 3402 237064 3408
rect 235908 3120 235960 3126
rect 235908 3062 235960 3068
rect 237024 480 237052 3402
rect 237300 3194 237328 38966
rect 238036 4894 238064 39306
rect 238772 39030 238800 41806
rect 239600 39098 239628 41806
rect 239588 39092 239640 39098
rect 239588 39034 239640 39040
rect 240520 39030 240548 41806
rect 238668 39024 238720 39030
rect 238668 38966 238720 38972
rect 238760 39024 238812 39030
rect 238760 38966 238812 38972
rect 240048 39024 240100 39030
rect 240048 38966 240100 38972
rect 240508 39024 240560 39030
rect 240508 38966 240560 38972
rect 238024 4888 238076 4894
rect 238024 4830 238076 4836
rect 238116 3256 238168 3262
rect 238116 3198 238168 3204
rect 237288 3188 237340 3194
rect 237288 3130 237340 3136
rect 238128 480 238156 3198
rect 238680 3058 238708 38966
rect 239312 4888 239364 4894
rect 239312 4830 239364 4836
rect 238668 3052 238720 3058
rect 238668 2994 238720 3000
rect 239324 480 239352 4830
rect 240060 3466 240088 38966
rect 241348 3602 241376 41806
rect 242176 39710 242204 41806
rect 242164 39704 242216 39710
rect 242164 39646 242216 39652
rect 242164 39092 242216 39098
rect 242164 39034 242216 39040
rect 241428 39024 241480 39030
rect 241428 38966 241480 38972
rect 241336 3596 241388 3602
rect 241336 3538 241388 3544
rect 241440 3534 241468 38966
rect 242176 5098 242204 39034
rect 243096 39030 243124 41806
rect 243084 39024 243136 39030
rect 243084 38966 243136 38972
rect 244108 6914 244136 41806
rect 244752 39846 244780 41806
rect 244740 39840 244792 39846
rect 244740 39782 244792 39788
rect 244924 39568 244976 39574
rect 244924 39510 244976 39516
rect 244188 39024 244240 39030
rect 244188 38966 244240 38972
rect 244016 6886 244136 6914
rect 242164 5092 242216 5098
rect 242164 5034 242216 5040
rect 242900 4956 242952 4962
rect 242900 4898 242952 4904
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 240048 3460 240100 3466
rect 240048 3402 240100 3408
rect 240520 480 240548 3470
rect 241704 3392 241756 3398
rect 241704 3334 241756 3340
rect 241716 480 241744 3334
rect 242912 480 242940 4898
rect 244016 3398 244044 6886
rect 244004 3392 244056 3398
rect 244004 3334 244056 3340
rect 244096 3324 244148 3330
rect 244096 3266 244148 3272
rect 244108 480 244136 3266
rect 244200 3262 244228 38966
rect 244936 4418 244964 39510
rect 245672 39030 245700 41806
rect 246500 39370 246528 41806
rect 247328 39642 247356 41806
rect 247316 39636 247368 39642
rect 247316 39578 247368 39584
rect 246488 39364 246540 39370
rect 246488 39306 246540 39312
rect 245660 39024 245712 39030
rect 245660 38966 245712 38972
rect 246948 39024 247000 39030
rect 246948 38966 247000 38972
rect 246396 7608 246448 7614
rect 246396 7550 246448 7556
rect 244924 4412 244976 4418
rect 244924 4354 244976 4360
rect 245200 4004 245252 4010
rect 245200 3946 245252 3952
rect 244188 3256 244240 3262
rect 244188 3198 244240 3204
rect 245212 480 245240 3946
rect 246408 480 246436 7550
rect 246960 3330 246988 38966
rect 248340 4146 248368 41806
rect 248972 39636 249024 39642
rect 248972 39578 249024 39584
rect 248984 35894 249012 39578
rect 249076 39030 249104 41806
rect 249996 39030 250024 41806
rect 249064 39024 249116 39030
rect 249064 38966 249116 38972
rect 249708 39024 249760 39030
rect 249708 38966 249760 38972
rect 249984 39024 250036 39030
rect 249984 38966 250036 38972
rect 250996 39024 251048 39030
rect 250996 38966 251048 38972
rect 248984 35866 249104 35894
rect 249076 7682 249104 35866
rect 249064 7676 249116 7682
rect 249064 7618 249116 7624
rect 247592 4140 247644 4146
rect 247592 4082 247644 4088
rect 248328 4140 248380 4146
rect 248328 4082 248380 4088
rect 246948 3324 247000 3330
rect 246948 3266 247000 3272
rect 247604 480 247632 4082
rect 249720 4010 249748 38966
rect 251008 4962 251036 38966
rect 250996 4956 251048 4962
rect 250996 4898 251048 4904
rect 249984 4412 250036 4418
rect 249984 4354 250036 4360
rect 249708 4004 249760 4010
rect 249708 3946 249760 3952
rect 248788 3936 248840 3942
rect 248788 3878 248840 3884
rect 248800 480 248828 3878
rect 249996 480 250024 4354
rect 251100 3942 251128 41806
rect 251652 39030 251680 41806
rect 252572 39710 252600 41806
rect 251824 39704 251876 39710
rect 251824 39646 251876 39652
rect 252560 39704 252612 39710
rect 252560 39646 252612 39652
rect 251640 39024 251692 39030
rect 251640 38966 251692 38972
rect 251836 4758 251864 39646
rect 253400 39030 253428 41806
rect 254228 39030 254256 41806
rect 255148 39982 255176 41806
rect 255136 39976 255188 39982
rect 255136 39918 255188 39924
rect 255872 39432 255924 39438
rect 255872 39374 255924 39380
rect 252468 39024 252520 39030
rect 252468 38966 252520 38972
rect 253388 39024 253440 39030
rect 253388 38966 253440 38972
rect 253848 39024 253900 39030
rect 253848 38966 253900 38972
rect 254216 39024 254268 39030
rect 254216 38966 254268 38972
rect 255228 39024 255280 39030
rect 255228 38966 255280 38972
rect 251824 4752 251876 4758
rect 251824 4694 251876 4700
rect 252480 4078 252508 38966
rect 253860 4894 253888 38966
rect 253848 4888 253900 4894
rect 253848 4830 253900 4836
rect 253480 4820 253532 4826
rect 253480 4762 253532 4768
rect 252376 4072 252428 4078
rect 252376 4014 252428 4020
rect 252468 4072 252520 4078
rect 252468 4014 252520 4020
rect 251088 3936 251140 3942
rect 251088 3878 251140 3884
rect 251180 2848 251232 2854
rect 251180 2790 251232 2796
rect 251192 480 251220 2790
rect 252388 480 252416 4014
rect 253492 480 253520 4762
rect 255240 3874 255268 38966
rect 255884 35894 255912 39374
rect 255976 39030 256004 41806
rect 256804 39574 256832 41806
rect 257724 39778 257752 41806
rect 257712 39772 257764 39778
rect 257712 39714 257764 39720
rect 256792 39568 256844 39574
rect 256792 39510 256844 39516
rect 258552 39302 258580 41806
rect 258540 39296 258592 39302
rect 258540 39238 258592 39244
rect 255964 39024 256016 39030
rect 255964 38966 256016 38972
rect 256608 39024 256660 39030
rect 256608 38966 256660 38972
rect 255884 35866 256004 35894
rect 255976 4214 256004 35866
rect 256620 5370 256648 38966
rect 256608 5364 256660 5370
rect 256608 5306 256660 5312
rect 255964 4208 256016 4214
rect 255964 4150 256016 4156
rect 257068 4208 257120 4214
rect 257068 4150 257120 4156
rect 254676 3868 254728 3874
rect 254676 3810 254728 3816
rect 255228 3868 255280 3874
rect 255228 3810 255280 3816
rect 254688 480 254716 3810
rect 255872 2916 255924 2922
rect 255872 2858 255924 2864
rect 255884 480 255912 2858
rect 257080 480 257108 4150
rect 259380 3738 259408 41806
rect 260300 39030 260328 41806
rect 261128 39030 261156 41806
rect 260288 39024 260340 39030
rect 260288 38966 260340 38972
rect 260748 39024 260800 39030
rect 260748 38966 260800 38972
rect 261116 39024 261168 39030
rect 261116 38966 261168 38972
rect 260656 10328 260708 10334
rect 260656 10270 260708 10276
rect 259460 3800 259512 3806
rect 259460 3742 259512 3748
rect 258264 3732 258316 3738
rect 258264 3674 258316 3680
rect 259368 3732 259420 3738
rect 259368 3674 259420 3680
rect 258276 480 258304 3674
rect 259472 480 259500 3742
rect 260668 480 260696 10270
rect 260760 4826 260788 38966
rect 260748 4820 260800 4826
rect 260748 4762 260800 4768
rect 262140 3806 262168 41806
rect 262784 41806 262858 41834
rect 263658 41834 263686 42092
rect 264578 41834 264606 42092
rect 265406 41834 265434 42092
rect 266234 41834 266262 42092
rect 267154 41834 267182 42092
rect 267982 41834 268010 42092
rect 268810 41834 268838 42092
rect 269730 41834 269758 42092
rect 270558 41834 270586 42092
rect 271478 41834 271506 42092
rect 272306 41834 272334 42092
rect 273134 41834 273162 42092
rect 274054 41834 274082 42092
rect 274882 41834 274910 42092
rect 275710 41834 275738 42092
rect 276630 41834 276658 42092
rect 277458 41834 277486 42092
rect 278286 41834 278314 42092
rect 279206 41834 279234 42092
rect 280034 41834 280062 42092
rect 280954 41834 280982 42092
rect 281782 41834 281810 42092
rect 282610 41834 282638 42092
rect 283530 41834 283558 42092
rect 284358 41834 284386 42092
rect 285186 41834 285214 42092
rect 286106 41834 286134 42092
rect 286934 41834 286962 42092
rect 263658 41806 263732 41834
rect 264578 41806 264928 41834
rect 265406 41806 265480 41834
rect 266234 41806 266308 41834
rect 267154 41806 267228 41834
rect 267982 41806 268056 41834
rect 268810 41806 269068 41834
rect 269730 41806 269804 41834
rect 270558 41806 270632 41834
rect 271478 41806 271736 41834
rect 272306 41806 272380 41834
rect 273134 41806 273208 41834
rect 274054 41806 274128 41834
rect 274882 41806 274956 41834
rect 275710 41806 275784 41834
rect 276630 41806 276704 41834
rect 277458 41806 277532 41834
rect 278286 41806 278636 41834
rect 279206 41806 279280 41834
rect 280034 41806 280108 41834
rect 280954 41806 281028 41834
rect 281782 41806 281856 41834
rect 282610 41806 282684 41834
rect 283530 41806 283604 41834
rect 284358 41806 284432 41834
rect 285186 41806 285628 41834
rect 286106 41806 286180 41834
rect 262784 39642 262812 41806
rect 262864 39840 262916 39846
rect 262864 39782 262916 39788
rect 262772 39636 262824 39642
rect 262772 39578 262824 39584
rect 262876 4554 262904 39782
rect 263704 39030 263732 41806
rect 262956 39024 263008 39030
rect 262956 38966 263008 38972
rect 263692 39024 263744 39030
rect 263692 38966 263744 38972
rect 264796 39024 264848 39030
rect 264796 38966 264848 38972
rect 262968 6322 262996 38966
rect 264808 9042 264836 38966
rect 264796 9036 264848 9042
rect 264796 8978 264848 8984
rect 262956 6316 263008 6322
rect 262956 6258 263008 6264
rect 264152 5024 264204 5030
rect 264152 4966 264204 4972
rect 262864 4548 262916 4554
rect 262864 4490 262916 4496
rect 262128 3800 262180 3806
rect 262128 3742 262180 3748
rect 262956 3664 263008 3670
rect 262956 3606 263008 3612
rect 261760 2984 261812 2990
rect 261760 2926 261812 2932
rect 261772 480 261800 2926
rect 262968 480 262996 3606
rect 264164 480 264192 4966
rect 264900 3670 264928 41806
rect 265452 39030 265480 41806
rect 266280 40050 266308 41806
rect 266268 40044 266320 40050
rect 266268 39986 266320 39992
rect 267096 39500 267148 39506
rect 267096 39442 267148 39448
rect 265440 39024 265492 39030
rect 265440 38966 265492 38972
rect 267004 39024 267056 39030
rect 267004 38966 267056 38972
rect 267016 5302 267044 38966
rect 267004 5296 267056 5302
rect 267004 5238 267056 5244
rect 267108 5030 267136 39442
rect 267200 39438 267228 41806
rect 268028 39982 268056 41806
rect 268016 39976 268068 39982
rect 268016 39918 268068 39924
rect 267188 39432 267240 39438
rect 267188 39374 267240 39380
rect 268384 39296 268436 39302
rect 268384 39238 268436 39244
rect 268396 5438 268424 39238
rect 269040 6254 269068 41806
rect 269672 39908 269724 39914
rect 269672 39850 269724 39856
rect 269684 35894 269712 39850
rect 269776 39030 269804 41806
rect 270604 39030 270632 41806
rect 269764 39024 269816 39030
rect 269764 38966 269816 38972
rect 270408 39024 270460 39030
rect 270408 38966 270460 38972
rect 270592 39024 270644 39030
rect 270592 38966 270644 38972
rect 269684 35866 269804 35894
rect 269028 6248 269080 6254
rect 269028 6190 269080 6196
rect 269776 5506 269804 35866
rect 269764 5500 269816 5506
rect 269764 5442 269816 5448
rect 268384 5432 268436 5438
rect 268384 5374 268436 5380
rect 267096 5024 267148 5030
rect 267096 4966 267148 4972
rect 267740 5024 267792 5030
rect 267740 4966 267792 4972
rect 264888 3664 264940 3670
rect 264888 3606 264940 3612
rect 266544 3188 266596 3194
rect 266544 3130 266596 3136
rect 265348 3120 265400 3126
rect 265348 3062 265400 3068
rect 265360 480 265388 3062
rect 266556 480 266584 3130
rect 267752 480 267780 4966
rect 270420 3466 270448 38966
rect 271708 5166 271736 41806
rect 272352 39030 272380 41806
rect 273180 39506 273208 41806
rect 273904 39704 273956 39710
rect 273904 39646 273956 39652
rect 273168 39500 273220 39506
rect 273168 39442 273220 39448
rect 271788 39024 271840 39030
rect 271788 38966 271840 38972
rect 272340 39024 272392 39030
rect 272340 38966 272392 38972
rect 273168 39024 273220 39030
rect 273168 38966 273220 38972
rect 271800 5234 271828 38966
rect 271788 5228 271840 5234
rect 271788 5170 271840 5176
rect 271696 5160 271748 5166
rect 271696 5102 271748 5108
rect 271236 5092 271288 5098
rect 271236 5034 271288 5040
rect 270040 3460 270092 3466
rect 270040 3402 270092 3408
rect 270408 3460 270460 3466
rect 270408 3402 270460 3408
rect 268844 3052 268896 3058
rect 268844 2994 268896 3000
rect 268856 480 268884 2994
rect 270052 480 270080 3402
rect 271248 480 271276 5034
rect 273180 3534 273208 38966
rect 273916 4622 273944 39646
rect 274100 39030 274128 41806
rect 274928 39030 274956 41806
rect 275756 39846 275784 41806
rect 275744 39840 275796 39846
rect 275744 39782 275796 39788
rect 276572 39772 276624 39778
rect 276572 39714 276624 39720
rect 274088 39024 274140 39030
rect 274088 38966 274140 38972
rect 274548 39024 274600 39030
rect 274548 38966 274600 38972
rect 274916 39024 274968 39030
rect 274916 38966 274968 38972
rect 275928 39024 275980 39030
rect 275928 38966 275980 38972
rect 274560 6186 274588 38966
rect 274548 6180 274600 6186
rect 274548 6122 274600 6128
rect 274824 4752 274876 4758
rect 274824 4694 274876 4700
rect 273904 4616 273956 4622
rect 273904 4558 273956 4564
rect 273628 3596 273680 3602
rect 273628 3538 273680 3544
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 273168 3528 273220 3534
rect 273168 3470 273220 3476
rect 272444 480 272472 3470
rect 273640 480 273668 3538
rect 274836 480 274864 4694
rect 275940 3602 275968 38966
rect 276584 35894 276612 39714
rect 276676 39030 276704 41806
rect 277504 39030 277532 41806
rect 276664 39024 276716 39030
rect 276664 38966 276716 38972
rect 277308 39024 277360 39030
rect 277308 38966 277360 38972
rect 277492 39024 277544 39030
rect 277492 38966 277544 38972
rect 276584 35866 276704 35894
rect 276676 4690 276704 35866
rect 277320 7614 277348 38966
rect 278608 10334 278636 41806
rect 279252 39030 279280 41806
rect 280080 39778 280108 41806
rect 280068 39772 280120 39778
rect 280068 39714 280120 39720
rect 280252 39364 280304 39370
rect 280252 39306 280304 39312
rect 278688 39024 278740 39030
rect 278688 38966 278740 38972
rect 279240 39024 279292 39030
rect 279240 38966 279292 38972
rect 278596 10328 278648 10334
rect 278596 10270 278648 10276
rect 277308 7608 277360 7614
rect 277308 7550 277360 7556
rect 276664 4684 276716 4690
rect 276664 4626 276716 4632
rect 278320 4548 278372 4554
rect 278320 4490 278372 4496
rect 275928 3596 275980 3602
rect 275928 3538 275980 3544
rect 277124 3392 277176 3398
rect 277124 3334 277176 3340
rect 276020 3256 276072 3262
rect 276020 3198 276072 3204
rect 276032 480 276060 3198
rect 277136 480 277164 3334
rect 278332 480 278360 4490
rect 278700 3194 278728 38966
rect 280264 16574 280292 39306
rect 281000 39030 281028 41806
rect 281828 39846 281856 41806
rect 281816 39840 281868 39846
rect 281816 39782 281868 39788
rect 282184 39500 282236 39506
rect 282184 39442 282236 39448
rect 280804 39024 280856 39030
rect 280804 38966 280856 38972
rect 280988 39024 281040 39030
rect 280988 38966 281040 38972
rect 281448 39024 281500 39030
rect 281448 38966 281500 38972
rect 280816 21418 280844 38966
rect 280804 21412 280856 21418
rect 280804 21354 280856 21360
rect 280264 16546 280752 16574
rect 279516 3324 279568 3330
rect 279516 3266 279568 3272
rect 278688 3188 278740 3194
rect 278688 3130 278740 3136
rect 279528 480 279556 3266
rect 280724 480 280752 16546
rect 281460 5098 281488 38966
rect 282196 7682 282224 39442
rect 282656 39370 282684 41806
rect 283576 39710 283604 41806
rect 283564 39704 283616 39710
rect 283564 39646 283616 39652
rect 282644 39364 282696 39370
rect 282644 39306 282696 39312
rect 284404 38962 284432 41806
rect 284392 38956 284444 38962
rect 284392 38898 284444 38904
rect 285496 38956 285548 38962
rect 285496 38898 285548 38904
rect 281908 7676 281960 7682
rect 281908 7618 281960 7624
rect 282184 7676 282236 7682
rect 282184 7618 282236 7624
rect 281448 5092 281500 5098
rect 281448 5034 281500 5040
rect 281920 480 281948 7618
rect 285508 4962 285536 38898
rect 285404 4956 285456 4962
rect 285404 4898 285456 4904
rect 285496 4956 285548 4962
rect 285496 4898 285548 4904
rect 283104 4140 283156 4146
rect 283104 4082 283156 4088
rect 283116 480 283144 4082
rect 284300 4004 284352 4010
rect 284300 3946 284352 3952
rect 284312 480 284340 3946
rect 285416 480 285444 4898
rect 285600 3262 285628 41806
rect 286152 39030 286180 41806
rect 286888 41806 286962 41834
rect 287762 41834 287790 42092
rect 288682 41834 288710 42092
rect 289510 41834 289538 42092
rect 290338 41834 290366 42092
rect 291258 41834 291286 42092
rect 292086 41834 292114 42092
rect 293006 41834 293034 42092
rect 293834 41834 293862 42092
rect 294662 41834 294690 42092
rect 295582 41834 295610 42092
rect 296410 41834 296438 42092
rect 297238 41834 297266 42092
rect 298158 41834 298186 42092
rect 298986 41834 299014 42092
rect 299814 41834 299842 42092
rect 300734 41834 300762 42092
rect 301562 41834 301590 42092
rect 302482 41834 302510 42092
rect 303310 41834 303338 42092
rect 304138 41834 304166 42092
rect 305058 41834 305086 42092
rect 305886 41834 305914 42092
rect 306714 41834 306742 42092
rect 307634 41834 307662 42092
rect 308462 41834 308490 42092
rect 309290 41834 309318 42092
rect 310210 41834 310238 42092
rect 311038 41834 311066 42092
rect 311958 41834 311986 42092
rect 312786 41834 312814 42092
rect 313614 41834 313642 42092
rect 314534 41834 314562 42092
rect 287762 41806 287836 41834
rect 288682 41806 288756 41834
rect 289510 41806 289584 41834
rect 290338 41806 290412 41834
rect 291258 41806 291332 41834
rect 292086 41806 292436 41834
rect 293006 41806 293080 41834
rect 293834 41806 293908 41834
rect 294662 41806 294736 41834
rect 295582 41806 295656 41834
rect 296410 41806 296576 41834
rect 297238 41806 297312 41834
rect 298158 41806 298232 41834
rect 298986 41806 299336 41834
rect 299814 41806 299888 41834
rect 300734 41806 300808 41834
rect 301562 41806 301636 41834
rect 302482 41806 302556 41834
rect 303310 41806 303568 41834
rect 304138 41806 304212 41834
rect 305058 41806 305132 41834
rect 305886 41806 306328 41834
rect 306714 41806 306788 41834
rect 307634 41806 307708 41834
rect 308462 41806 308536 41834
rect 309290 41806 309364 41834
rect 310210 41806 310376 41834
rect 311038 41806 311112 41834
rect 311958 41806 312032 41834
rect 312786 41806 313228 41834
rect 313614 41806 313688 41834
rect 286140 39024 286192 39030
rect 286140 38966 286192 38972
rect 286888 17338 286916 41806
rect 287704 39636 287756 39642
rect 287704 39578 287756 39584
rect 286968 39024 287020 39030
rect 286968 38966 287020 38972
rect 286876 17332 286928 17338
rect 286876 17274 286928 17280
rect 286980 5030 287008 38966
rect 286968 5024 287020 5030
rect 286968 4966 287020 4972
rect 287716 4554 287744 39578
rect 287808 38826 287836 41806
rect 288728 39030 288756 41806
rect 289556 39642 289584 41806
rect 289544 39636 289596 39642
rect 289544 39578 289596 39584
rect 289084 39296 289136 39302
rect 289084 39238 289136 39244
rect 288716 39024 288768 39030
rect 288716 38966 288768 38972
rect 287796 38820 287848 38826
rect 287796 38762 287848 38768
rect 288348 38820 288400 38826
rect 288348 38762 288400 38768
rect 287704 4548 287756 4554
rect 287704 4490 287756 4496
rect 287796 4072 287848 4078
rect 287796 4014 287848 4020
rect 286600 3936 286652 3942
rect 286600 3878 286652 3884
rect 285588 3256 285640 3262
rect 285588 3198 285640 3204
rect 286612 480 286640 3878
rect 287808 480 287836 4014
rect 288360 3330 288388 38762
rect 289096 4758 289124 39238
rect 290384 39030 290412 41806
rect 291304 39030 291332 41806
rect 289728 39024 289780 39030
rect 289728 38966 289780 38972
rect 290372 39024 290424 39030
rect 290372 38966 290424 38972
rect 291108 39024 291160 39030
rect 291108 38966 291160 38972
rect 291292 39024 291344 39030
rect 291292 38966 291344 38972
rect 289740 15978 289768 38966
rect 289728 15972 289780 15978
rect 289728 15914 289780 15920
rect 290188 4888 290240 4894
rect 290188 4830 290240 4836
rect 289084 4752 289136 4758
rect 289084 4694 289136 4700
rect 288992 4616 289044 4622
rect 288992 4558 289044 4564
rect 288348 3324 288400 3330
rect 288348 3266 288400 3272
rect 289004 480 289032 4558
rect 290200 480 290228 4830
rect 291120 4146 291148 38966
rect 292408 6662 292436 41806
rect 293052 39030 293080 41806
rect 293880 39506 293908 41806
rect 293960 39568 294012 39574
rect 293960 39510 294012 39516
rect 293868 39500 293920 39506
rect 293868 39442 293920 39448
rect 292488 39024 292540 39030
rect 292488 38966 292540 38972
rect 293040 39024 293092 39030
rect 293040 38966 293092 38972
rect 293868 39024 293920 39030
rect 293868 38966 293920 38972
rect 292396 6656 292448 6662
rect 292396 6598 292448 6604
rect 292500 4894 292528 38966
rect 292580 5500 292632 5506
rect 292580 5442 292632 5448
rect 292488 4888 292540 4894
rect 292488 4830 292540 4836
rect 291108 4140 291160 4146
rect 291108 4082 291160 4088
rect 291384 3868 291436 3874
rect 291384 3810 291436 3816
rect 291396 480 291424 3810
rect 292592 480 292620 5442
rect 293684 5364 293736 5370
rect 293684 5306 293736 5312
rect 293696 480 293724 5306
rect 293880 3398 293908 38966
rect 293972 16574 294000 39510
rect 294708 39302 294736 41806
rect 294696 39296 294748 39302
rect 294696 39238 294748 39244
rect 295628 39030 295656 41806
rect 295616 39024 295668 39030
rect 295616 38966 295668 38972
rect 293972 16546 294920 16574
rect 293868 3392 293920 3398
rect 293868 3334 293920 3340
rect 294892 480 294920 16546
rect 296548 8974 296576 41806
rect 297284 40050 297312 41806
rect 297272 40044 297324 40050
rect 297272 39986 297324 39992
rect 298204 39030 298232 41806
rect 299204 40044 299256 40050
rect 299204 39986 299256 39992
rect 296628 39024 296680 39030
rect 296628 38966 296680 38972
rect 298192 39024 298244 39030
rect 298192 38966 298244 38972
rect 296536 8968 296588 8974
rect 296536 8910 296588 8916
rect 296076 4684 296128 4690
rect 296076 4626 296128 4632
rect 296088 480 296116 4626
rect 296640 4010 296668 38966
rect 299216 37942 299244 39986
rect 299204 37936 299256 37942
rect 299204 37878 299256 37884
rect 299308 13122 299336 41806
rect 299860 39030 299888 41806
rect 299388 39024 299440 39030
rect 299388 38966 299440 38972
rect 299848 39024 299900 39030
rect 299848 38966 299900 38972
rect 300676 39024 300728 39030
rect 300676 38966 300728 38972
rect 299296 13116 299348 13122
rect 299296 13058 299348 13064
rect 297272 5432 297324 5438
rect 297272 5374 297324 5380
rect 296628 4004 296680 4010
rect 296628 3946 296680 3952
rect 297284 480 297312 5374
rect 299400 4078 299428 38966
rect 300688 6594 300716 38966
rect 300676 6588 300728 6594
rect 300676 6530 300728 6536
rect 300676 6316 300728 6322
rect 300676 6258 300728 6264
rect 299664 4820 299716 4826
rect 299664 4762 299716 4768
rect 299388 4072 299440 4078
rect 299388 4014 299440 4020
rect 298468 3732 298520 3738
rect 298468 3674 298520 3680
rect 298480 480 298508 3674
rect 299676 480 299704 4762
rect 300688 3210 300716 6258
rect 300780 3874 300808 41806
rect 301608 40050 301636 41806
rect 301596 40044 301648 40050
rect 301596 39986 301648 39992
rect 302528 39030 302556 41806
rect 302516 39024 302568 39030
rect 302516 38966 302568 38972
rect 303436 39024 303488 39030
rect 303436 38966 303488 38972
rect 303448 4826 303476 38966
rect 303436 4820 303488 4826
rect 303436 4762 303488 4768
rect 303160 4548 303212 4554
rect 303160 4490 303212 4496
rect 300768 3868 300820 3874
rect 300768 3810 300820 3816
rect 301964 3800 302016 3806
rect 301964 3742 302016 3748
rect 300688 3182 300808 3210
rect 300780 480 300808 3182
rect 301976 480 302004 3742
rect 303172 480 303200 4490
rect 303540 3942 303568 41806
rect 304184 38894 304212 41806
rect 304264 39976 304316 39982
rect 304264 39918 304316 39924
rect 304172 38888 304224 38894
rect 304172 38830 304224 38836
rect 304276 5370 304304 39918
rect 305104 39030 305132 41806
rect 305092 39024 305144 39030
rect 305092 38966 305144 38972
rect 306196 39024 306248 39030
rect 306196 38966 306248 38972
rect 304908 38888 304960 38894
rect 304908 38830 304960 38836
rect 304920 11762 304948 38830
rect 304908 11756 304960 11762
rect 304908 11698 304960 11704
rect 304356 9036 304408 9042
rect 304356 8978 304408 8984
rect 304264 5364 304316 5370
rect 304264 5306 304316 5312
rect 303528 3936 303580 3942
rect 303528 3878 303580 3884
rect 304368 480 304396 8978
rect 306208 6526 306236 38966
rect 306196 6520 306248 6526
rect 306196 6462 306248 6468
rect 306300 3806 306328 41806
rect 306760 39030 306788 41806
rect 307680 39574 307708 41806
rect 307668 39568 307720 39574
rect 307668 39510 307720 39516
rect 307760 39432 307812 39438
rect 307760 39374 307812 39380
rect 307024 39296 307076 39302
rect 307024 39238 307076 39244
rect 306748 39024 306800 39030
rect 306748 38966 306800 38972
rect 307036 5302 307064 39238
rect 307668 39024 307720 39030
rect 307668 38966 307720 38972
rect 307680 14482 307708 38966
rect 307668 14476 307720 14482
rect 307668 14418 307720 14424
rect 306748 5296 306800 5302
rect 306748 5238 306800 5244
rect 307024 5296 307076 5302
rect 307024 5238 307076 5244
rect 306288 3800 306340 3806
rect 306288 3742 306340 3748
rect 305552 3664 305604 3670
rect 305552 3606 305604 3612
rect 305564 480 305592 3606
rect 306760 480 306788 5238
rect 307772 3466 307800 39374
rect 308508 38962 308536 41806
rect 309336 39030 309364 41806
rect 309324 39024 309376 39030
rect 309324 38966 309376 38972
rect 308496 38956 308548 38962
rect 308496 38898 308548 38904
rect 309048 38956 309100 38962
rect 309048 38898 309100 38904
rect 309060 6914 309088 38898
rect 310348 7886 310376 41806
rect 311084 39030 311112 41806
rect 312004 39302 312032 41806
rect 311992 39296 312044 39302
rect 311992 39238 312044 39244
rect 310428 39024 310480 39030
rect 310428 38966 310480 38972
rect 311072 39024 311124 39030
rect 311072 38966 311124 38972
rect 311808 39024 311860 39030
rect 311808 38966 311860 38972
rect 310336 7880 310388 7886
rect 310336 7822 310388 7828
rect 308968 6886 309088 6914
rect 307944 4684 307996 4690
rect 307944 4626 307996 4632
rect 307760 3460 307812 3466
rect 307760 3402 307812 3408
rect 307956 480 307984 4626
rect 308968 3670 308996 6886
rect 310440 6458 310468 38966
rect 310428 6452 310480 6458
rect 310428 6394 310480 6400
rect 311440 6248 311492 6254
rect 311440 6190 311492 6196
rect 310244 5364 310296 5370
rect 310244 5306 310296 5312
rect 308956 3664 309008 3670
rect 308956 3606 309008 3612
rect 309048 3460 309100 3466
rect 309048 3402 309100 3408
rect 309060 480 309088 3402
rect 310256 480 310284 5306
rect 311452 480 311480 6190
rect 311820 3738 311848 38966
rect 313200 6390 313228 41806
rect 313660 39030 313688 41806
rect 314488 41806 314562 41834
rect 315362 41834 315390 42092
rect 316190 41834 316218 42092
rect 317110 41834 317138 42092
rect 317938 41834 317966 42092
rect 318766 41834 318794 42092
rect 319686 41834 319714 42092
rect 320514 41834 320542 42092
rect 321342 41834 321370 42092
rect 322262 41834 322290 42092
rect 323090 41834 323118 42092
rect 324010 41834 324038 42092
rect 324838 41834 324866 42092
rect 325666 41834 325694 42092
rect 326586 41834 326614 42092
rect 327414 41834 327442 42092
rect 328242 41834 328270 42092
rect 329162 41834 329190 42092
rect 329990 41834 330018 42092
rect 330818 41834 330846 42092
rect 331738 41834 331766 42092
rect 332566 41834 332594 42092
rect 333486 41834 333514 42092
rect 334314 41834 334342 42092
rect 335142 41834 335170 42092
rect 336062 41834 336090 42092
rect 336890 41834 336918 42092
rect 337718 41834 337746 42092
rect 338638 41834 338666 42092
rect 339466 41834 339494 42092
rect 340294 41834 340322 42092
rect 341214 41834 341242 42092
rect 342042 41834 342070 42092
rect 342962 41834 342990 42092
rect 343790 41834 343818 42092
rect 344618 41834 344646 42092
rect 345538 41834 345566 42092
rect 346366 41834 346394 42092
rect 347194 41834 347222 42092
rect 348114 41834 348142 42092
rect 348942 41834 348970 42092
rect 349770 41834 349798 42092
rect 350690 41834 350718 42092
rect 351518 41834 351546 42092
rect 352346 41834 352374 42092
rect 353266 41834 353294 42092
rect 354094 41834 354122 42092
rect 355014 41834 355042 42092
rect 355842 41834 355870 42092
rect 356670 41834 356698 42092
rect 357590 41834 357618 42092
rect 358418 41834 358446 42092
rect 359246 41834 359274 42092
rect 360166 41834 360194 42092
rect 360994 41834 361022 42092
rect 361822 41834 361850 42092
rect 362742 41834 362770 42092
rect 363570 41834 363598 42092
rect 364490 41834 364518 42092
rect 365318 41834 365346 42092
rect 366146 41834 366174 42092
rect 367066 41834 367094 42092
rect 367894 41834 367922 42092
rect 368722 41834 368750 42092
rect 369642 41834 369670 42092
rect 370470 41834 370498 42092
rect 371298 41834 371326 42092
rect 372218 41834 372246 42092
rect 373046 41834 373074 42092
rect 373966 41834 373994 42092
rect 374794 41834 374822 42092
rect 375622 41834 375650 42092
rect 376542 41834 376570 42092
rect 377370 41834 377398 42092
rect 378198 41834 378226 42092
rect 379118 41834 379146 42092
rect 379946 41834 379974 42092
rect 380774 41834 380802 42092
rect 381694 41834 381722 42092
rect 382522 41834 382550 42092
rect 383350 41834 383378 42092
rect 384270 41834 384298 42092
rect 385098 41834 385126 42092
rect 386018 41834 386046 42092
rect 386846 41834 386874 42092
rect 387674 41834 387702 42092
rect 388594 41834 388622 42092
rect 389422 41834 389450 42092
rect 390250 41834 390278 42092
rect 391170 41834 391198 42092
rect 391998 41834 392026 42092
rect 392826 41834 392854 42092
rect 393746 41834 393774 42092
rect 394574 41834 394602 42092
rect 395494 41834 395522 42092
rect 396322 41834 396350 42092
rect 397150 41834 397178 42092
rect 398070 41834 398098 42092
rect 398898 41834 398926 42092
rect 399726 41834 399754 42092
rect 400646 41834 400674 42092
rect 401474 41834 401502 42092
rect 315362 41806 315436 41834
rect 316190 41806 316264 41834
rect 317110 41806 317276 41834
rect 317938 41806 318012 41834
rect 318766 41806 318840 41834
rect 319686 41806 319760 41834
rect 320514 41806 320588 41834
rect 321342 41806 321508 41834
rect 322262 41806 322336 41834
rect 323090 41806 323164 41834
rect 324010 41806 324268 41834
rect 324838 41806 324912 41834
rect 325666 41806 325740 41834
rect 326586 41806 326660 41834
rect 327414 41806 327488 41834
rect 328242 41806 328408 41834
rect 329162 41806 329236 41834
rect 329990 41806 330064 41834
rect 330818 41806 330892 41834
rect 331738 41806 331812 41834
rect 332566 41806 332640 41834
rect 333486 41806 333560 41834
rect 334314 41806 334388 41834
rect 335142 41806 335216 41834
rect 336062 41806 336136 41834
rect 336890 41806 336964 41834
rect 337718 41806 337976 41834
rect 338638 41806 338712 41834
rect 339466 41806 339540 41834
rect 340294 41806 340736 41834
rect 341214 41806 341288 41834
rect 342042 41806 342208 41834
rect 342962 41806 343036 41834
rect 343790 41806 343864 41834
rect 344618 41806 344968 41834
rect 345538 41806 345612 41834
rect 346366 41806 346440 41834
rect 347194 41806 347268 41834
rect 348114 41806 348188 41834
rect 348942 41806 349016 41834
rect 349770 41806 349844 41834
rect 350690 41806 350764 41834
rect 351518 41806 351592 41834
rect 352346 41806 352420 41834
rect 353266 41806 353340 41834
rect 354094 41806 354536 41834
rect 355014 41806 355088 41834
rect 355842 41806 355916 41834
rect 356670 41806 356744 41834
rect 357590 41806 357664 41834
rect 358418 41806 358676 41834
rect 359246 41806 359320 41834
rect 360166 41806 360240 41834
rect 360994 41806 361436 41834
rect 361822 41806 361896 41834
rect 362742 41806 362908 41834
rect 363570 41806 363644 41834
rect 364490 41806 364564 41834
rect 365318 41806 365668 41834
rect 366146 41806 366220 41834
rect 367066 41806 367140 41834
rect 367894 41806 367968 41834
rect 368722 41806 368796 41834
rect 369642 41806 369716 41834
rect 370470 41806 370544 41834
rect 371298 41806 371372 41834
rect 372218 41806 372476 41834
rect 373046 41806 373120 41834
rect 373966 41806 374040 41834
rect 374794 41806 375236 41834
rect 375622 41806 375696 41834
rect 376542 41806 376616 41834
rect 377370 41806 377444 41834
rect 378198 41806 378272 41834
rect 379118 41806 379376 41834
rect 379946 41806 380020 41834
rect 380774 41806 380848 41834
rect 381694 41806 381768 41834
rect 382522 41806 382596 41834
rect 383350 41806 383608 41834
rect 384270 41806 384344 41834
rect 385098 41806 385172 41834
rect 386018 41806 386276 41834
rect 386846 41806 386920 41834
rect 387674 41806 387748 41834
rect 388594 41806 388668 41834
rect 389422 41806 389496 41834
rect 390250 41806 390416 41834
rect 391170 41806 391244 41834
rect 391998 41806 392072 41834
rect 392826 41806 393268 41834
rect 393746 41806 393820 41834
rect 394574 41806 394648 41834
rect 395494 41806 395568 41834
rect 396322 41806 396396 41834
rect 397150 41806 397224 41834
rect 398070 41806 398144 41834
rect 398898 41806 398972 41834
rect 399726 41806 400168 41834
rect 400646 41806 400720 41834
rect 313648 39024 313700 39030
rect 313648 38966 313700 38972
rect 313188 6384 313240 6390
rect 313188 6326 313240 6332
rect 314488 6322 314516 41806
rect 315408 39438 315436 41806
rect 315396 39432 315448 39438
rect 315396 39374 315448 39380
rect 316236 39030 316264 41806
rect 314568 39024 314620 39030
rect 314568 38966 314620 38972
rect 316224 39024 316276 39030
rect 316224 38966 316276 38972
rect 314476 6316 314528 6322
rect 314476 6258 314528 6264
rect 313832 5228 313884 5234
rect 313832 5170 313884 5176
rect 311808 3732 311860 3738
rect 311808 3674 311860 3680
rect 312636 3120 312688 3126
rect 312636 3062 312688 3068
rect 312648 480 312676 3062
rect 313844 480 313872 5170
rect 314580 3466 314608 38966
rect 317248 17270 317276 41806
rect 317984 39030 318012 41806
rect 318064 39908 318116 39914
rect 318064 39850 318116 39856
rect 317328 39024 317380 39030
rect 317328 38966 317380 38972
rect 317972 39024 318024 39030
rect 317972 38966 318024 38972
rect 317236 17264 317288 17270
rect 317236 17206 317288 17212
rect 317236 7676 317288 7682
rect 317236 7618 317288 7624
rect 315028 5160 315080 5166
rect 315028 5102 315080 5108
rect 314568 3460 314620 3466
rect 314568 3402 314620 3408
rect 315040 480 315068 5102
rect 316224 3528 316276 3534
rect 316224 3470 316276 3476
rect 317248 3482 317276 7618
rect 317340 3618 317368 38966
rect 318076 4214 318104 39850
rect 318812 39030 318840 41806
rect 319732 39982 319760 41806
rect 319720 39976 319772 39982
rect 319720 39918 319772 39924
rect 320560 39030 320588 41806
rect 318708 39024 318760 39030
rect 318708 38966 318760 38972
rect 318800 39024 318852 39030
rect 318800 38966 318852 38972
rect 320088 39024 320140 39030
rect 320088 38966 320140 38972
rect 320548 39024 320600 39030
rect 320548 38966 320600 38972
rect 321376 39024 321428 39030
rect 321376 38966 321428 38972
rect 318720 7818 318748 38966
rect 318708 7812 318760 7818
rect 318708 7754 318760 7760
rect 318524 6180 318576 6186
rect 318524 6122 318576 6128
rect 318064 4208 318116 4214
rect 318064 4150 318116 4156
rect 317340 3590 317460 3618
rect 317432 3534 317460 3590
rect 317420 3528 317472 3534
rect 316236 480 316264 3470
rect 317248 3454 317368 3482
rect 317420 3470 317472 3476
rect 317340 480 317368 3454
rect 318536 480 318564 6122
rect 320100 3602 320128 38966
rect 321388 7750 321416 38966
rect 321376 7744 321428 7750
rect 321376 7686 321428 7692
rect 320916 4208 320968 4214
rect 320916 4150 320968 4156
rect 319720 3596 319772 3602
rect 319720 3538 319772 3544
rect 320088 3596 320140 3602
rect 320088 3538 320140 3544
rect 319732 480 319760 3538
rect 320928 480 320956 4150
rect 321480 2854 321508 41806
rect 322204 40044 322256 40050
rect 322204 39986 322256 39992
rect 322216 7954 322244 39986
rect 322308 38962 322336 41806
rect 323136 39030 323164 41806
rect 323124 39024 323176 39030
rect 323124 38966 323176 38972
rect 324136 39024 324188 39030
rect 324136 38966 324188 38972
rect 322296 38956 322348 38962
rect 322296 38898 322348 38904
rect 322848 38956 322900 38962
rect 322848 38898 322900 38904
rect 322204 7948 322256 7954
rect 322204 7890 322256 7896
rect 322112 7608 322164 7614
rect 322112 7550 322164 7556
rect 321468 2848 321520 2854
rect 321468 2790 321520 2796
rect 322124 480 322152 7550
rect 322860 6254 322888 38898
rect 324148 7682 324176 38966
rect 324136 7676 324188 7682
rect 324136 7618 324188 7624
rect 322848 6248 322900 6254
rect 322848 6190 322900 6196
rect 324240 6186 324268 41806
rect 324884 39030 324912 41806
rect 325712 39914 325740 41806
rect 325700 39908 325752 39914
rect 325700 39850 325752 39856
rect 326632 39778 326660 41806
rect 327460 40050 327488 41806
rect 327448 40044 327500 40050
rect 327448 39986 327500 39992
rect 327724 39840 327776 39846
rect 327724 39782 327776 39788
rect 325700 39772 325752 39778
rect 325700 39714 325752 39720
rect 326620 39772 326672 39778
rect 326620 39714 326672 39720
rect 324964 39296 325016 39302
rect 324964 39238 325016 39244
rect 324872 39024 324924 39030
rect 324872 38966 324924 38972
rect 324320 21412 324372 21418
rect 324320 21354 324372 21360
rect 324228 6180 324280 6186
rect 324228 6122 324280 6128
rect 324332 3194 324360 21354
rect 324976 10334 325004 39238
rect 325608 39024 325660 39030
rect 325608 38966 325660 38972
rect 325620 21418 325648 38966
rect 325608 21412 325660 21418
rect 325608 21354 325660 21360
rect 325712 16574 325740 39714
rect 325712 16546 326384 16574
rect 324412 10328 324464 10334
rect 324412 10270 324464 10276
rect 324964 10328 325016 10334
rect 324964 10270 325016 10276
rect 323308 3188 323360 3194
rect 323308 3130 323360 3136
rect 324320 3188 324372 3194
rect 324320 3130 324372 3136
rect 323320 480 323348 3130
rect 324424 480 324452 10270
rect 325608 3188 325660 3194
rect 325608 3130 325660 3136
rect 325620 480 325648 3130
rect 326356 490 326384 16546
rect 327736 4214 327764 39782
rect 328380 22778 328408 41806
rect 329208 39030 329236 41806
rect 329932 39364 329984 39370
rect 329932 39306 329984 39312
rect 329196 39024 329248 39030
rect 329196 38966 329248 38972
rect 329748 39024 329800 39030
rect 329748 38966 329800 38972
rect 328368 22772 328420 22778
rect 328368 22714 328420 22720
rect 328000 5092 328052 5098
rect 328000 5034 328052 5040
rect 327724 4208 327776 4214
rect 327724 4150 327776 4156
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 5034
rect 329196 4208 329248 4214
rect 329196 4150 329248 4156
rect 329208 480 329236 4150
rect 329760 2922 329788 38966
rect 329944 16574 329972 39306
rect 330036 39030 330064 41806
rect 330864 39302 330892 41806
rect 331220 39704 331272 39710
rect 331220 39646 331272 39652
rect 330852 39296 330904 39302
rect 330852 39238 330904 39244
rect 330024 39024 330076 39030
rect 330024 38966 330076 38972
rect 331128 39024 331180 39030
rect 331128 38966 331180 38972
rect 329944 16546 330432 16574
rect 329748 2916 329800 2922
rect 329748 2858 329800 2864
rect 330404 480 330432 16546
rect 331140 4282 331168 38966
rect 331128 4276 331180 4282
rect 331128 4218 331180 4224
rect 331232 490 331260 39646
rect 331784 39030 331812 41806
rect 332612 39030 332640 41806
rect 333532 39710 333560 41806
rect 333520 39704 333572 39710
rect 333520 39646 333572 39652
rect 334360 39030 334388 41806
rect 331772 39024 331824 39030
rect 331772 38966 331824 38972
rect 332508 39024 332560 39030
rect 332508 38966 332560 38972
rect 332600 39024 332652 39030
rect 332600 38966 332652 38972
rect 333888 39024 333940 39030
rect 333888 38966 333940 38972
rect 334348 39024 334400 39030
rect 334348 38966 334400 38972
rect 332520 2990 332548 38966
rect 332692 4956 332744 4962
rect 332692 4898 332744 4904
rect 332508 2984 332560 2990
rect 332508 2926 332560 2932
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 4898
rect 333900 4350 333928 38966
rect 335084 5024 335136 5030
rect 335084 4966 335136 4972
rect 333888 4344 333940 4350
rect 333888 4286 333940 4292
rect 333888 3256 333940 3262
rect 333888 3198 333940 3204
rect 333900 480 333928 3198
rect 335096 480 335124 4966
rect 335188 4418 335216 41806
rect 336004 39840 336056 39846
rect 336004 39782 336056 39788
rect 335268 39024 335320 39030
rect 335268 38966 335320 38972
rect 335176 4412 335228 4418
rect 335176 4354 335228 4360
rect 335280 3058 335308 38966
rect 336016 18630 336044 39782
rect 336108 39030 336136 41806
rect 336936 39030 336964 41806
rect 336096 39024 336148 39030
rect 336096 38966 336148 38972
rect 336648 39024 336700 39030
rect 336648 38966 336700 38972
rect 336924 39024 336976 39030
rect 336924 38966 336976 38972
rect 336004 18624 336056 18630
rect 336004 18566 336056 18572
rect 335360 17332 335412 17338
rect 335360 17274 335412 17280
rect 335372 16574 335400 17274
rect 335372 16546 336320 16574
rect 335268 3052 335320 3058
rect 335268 2994 335320 3000
rect 336292 480 336320 16546
rect 336660 15910 336688 38966
rect 336648 15904 336700 15910
rect 336648 15846 336700 15852
rect 337948 4554 337976 41806
rect 338684 39030 338712 41806
rect 338764 39636 338816 39642
rect 338764 39578 338816 39584
rect 338028 39024 338080 39030
rect 338028 38966 338080 38972
rect 338672 39024 338724 39030
rect 338672 38966 338724 38972
rect 337936 4548 337988 4554
rect 337936 4490 337988 4496
rect 337476 3324 337528 3330
rect 337476 3266 337528 3272
rect 337488 480 337516 3266
rect 338040 3126 338068 38966
rect 338672 15972 338724 15978
rect 338672 15914 338724 15920
rect 338028 3120 338080 3126
rect 338028 3062 338080 3068
rect 338684 480 338712 15914
rect 338776 8294 338804 39578
rect 339512 39030 339540 41806
rect 339408 39024 339460 39030
rect 339408 38966 339460 38972
rect 339500 39024 339552 39030
rect 339500 38966 339552 38972
rect 339420 29646 339448 38966
rect 339408 29640 339460 29646
rect 339408 29582 339460 29588
rect 338764 8288 338816 8294
rect 338764 8230 338816 8236
rect 339868 8288 339920 8294
rect 339868 8230 339920 8236
rect 339880 480 339908 8230
rect 340708 4486 340736 41806
rect 341260 39030 341288 41806
rect 340788 39024 340840 39030
rect 340788 38966 340840 38972
rect 341248 39024 341300 39030
rect 341248 38966 341300 38972
rect 342076 39024 342128 39030
rect 342076 38966 342128 38972
rect 340696 4480 340748 4486
rect 340696 4422 340748 4428
rect 340800 3194 340828 38966
rect 342088 24138 342116 38966
rect 342076 24132 342128 24138
rect 342076 24074 342128 24080
rect 342180 6914 342208 41806
rect 342904 40044 342956 40050
rect 342904 39986 342956 39992
rect 342088 6886 342208 6914
rect 340972 4140 341024 4146
rect 340972 4082 341024 4088
rect 340788 3188 340840 3194
rect 340788 3130 340840 3136
rect 340984 480 341012 4082
rect 342088 3262 342116 6886
rect 342916 6050 342944 39986
rect 343008 39030 343036 41806
rect 343836 39982 343864 41806
rect 343824 39976 343876 39982
rect 343824 39918 343876 39924
rect 342996 39024 343048 39030
rect 342996 38966 343048 38972
rect 343548 39024 343600 39030
rect 343548 38966 343600 38972
rect 343364 6656 343416 6662
rect 343364 6598 343416 6604
rect 342904 6044 342956 6050
rect 342904 5986 342956 5992
rect 342168 4888 342220 4894
rect 342168 4830 342220 4836
rect 342076 3256 342128 3262
rect 342076 3198 342128 3204
rect 342180 480 342208 4830
rect 343376 480 343404 6598
rect 343560 4622 343588 38966
rect 343548 4616 343600 4622
rect 343548 4558 343600 4564
rect 344940 3398 344968 41806
rect 345020 39500 345072 39506
rect 345020 39442 345072 39448
rect 345032 16574 345060 39442
rect 345584 39030 345612 41806
rect 346412 39642 346440 41806
rect 346400 39636 346452 39642
rect 346400 39578 346452 39584
rect 347240 39030 347268 41806
rect 348160 39030 348188 41806
rect 348988 39846 349016 41806
rect 348976 39840 349028 39846
rect 348976 39782 349028 39788
rect 349712 39704 349764 39710
rect 349712 39646 349764 39652
rect 345572 39024 345624 39030
rect 345572 38966 345624 38972
rect 346308 39024 346360 39030
rect 346308 38966 346360 38972
rect 347228 39024 347280 39030
rect 347228 38966 347280 38972
rect 347688 39024 347740 39030
rect 347688 38966 347740 38972
rect 348148 39024 348200 39030
rect 348148 38966 348200 38972
rect 349068 39024 349120 39030
rect 349068 38966 349120 38972
rect 345032 16546 345336 16574
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 344928 3392 344980 3398
rect 344928 3334 344980 3340
rect 344572 480 344600 3334
rect 345308 490 345336 16546
rect 346320 4690 346348 38966
rect 346952 5296 347004 5302
rect 346952 5238 347004 5244
rect 346308 4684 346360 4690
rect 346308 4626 346360 4632
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 5238
rect 347700 4146 347728 38966
rect 349080 4758 349108 38966
rect 349724 37942 349752 39646
rect 349816 39030 349844 41806
rect 350736 39030 350764 41806
rect 351564 39710 351592 41806
rect 351552 39704 351604 39710
rect 351552 39646 351604 39652
rect 352392 39030 352420 41806
rect 352564 39976 352616 39982
rect 352564 39918 352616 39924
rect 349804 39024 349856 39030
rect 349804 38966 349856 38972
rect 350448 39024 350500 39030
rect 350448 38966 350500 38972
rect 350724 39024 350776 39030
rect 350724 38966 350776 38972
rect 351828 39024 351880 39030
rect 351828 38966 351880 38972
rect 352380 39024 352432 39030
rect 352380 38966 352432 38972
rect 349160 37936 349212 37942
rect 349160 37878 349212 37884
rect 349712 37936 349764 37942
rect 349712 37878 349764 37884
rect 349068 4752 349120 4758
rect 349068 4694 349120 4700
rect 347688 4140 347740 4146
rect 347688 4082 347740 4088
rect 348056 4004 348108 4010
rect 348056 3946 348108 3952
rect 348068 480 348096 3946
rect 349172 3330 349200 37878
rect 349252 8968 349304 8974
rect 349252 8910 349304 8916
rect 349160 3324 349212 3330
rect 349160 3266 349212 3272
rect 349264 480 349292 8910
rect 350460 4146 350488 38966
rect 351840 5438 351868 38966
rect 352576 13122 352604 39918
rect 353312 39030 353340 41806
rect 353208 39024 353260 39030
rect 353208 38966 353260 38972
rect 353300 39024 353352 39030
rect 353300 38966 353352 38972
rect 352564 13116 352616 13122
rect 352564 13058 352616 13064
rect 352840 13048 352892 13054
rect 352840 12990 352892 12996
rect 351828 5432 351880 5438
rect 351828 5374 351880 5380
rect 350448 4140 350500 4146
rect 350448 4082 350500 4088
rect 351644 4072 351696 4078
rect 351644 4014 351696 4020
rect 350448 3324 350500 3330
rect 350448 3266 350500 3272
rect 350460 480 350488 3266
rect 351656 480 351684 4014
rect 352852 480 352880 12990
rect 353220 4078 353248 38966
rect 354508 7614 354536 41806
rect 355060 39030 355088 41806
rect 354588 39024 354640 39030
rect 354588 38966 354640 38972
rect 355048 39024 355100 39030
rect 355048 38966 355100 38972
rect 354496 7608 354548 7614
rect 354496 7550 354548 7556
rect 354036 6588 354088 6594
rect 354036 6530 354088 6536
rect 353208 4072 353260 4078
rect 353208 4014 353260 4020
rect 354048 480 354076 6530
rect 354600 5506 354628 38966
rect 354588 5500 354640 5506
rect 354588 5442 354640 5448
rect 355888 5370 355916 41806
rect 356612 39568 356664 39574
rect 356612 39510 356664 39516
rect 355968 39024 356020 39030
rect 355968 38966 356020 38972
rect 355876 5364 355928 5370
rect 355876 5306 355928 5312
rect 355980 3874 356008 38966
rect 356624 35894 356652 39510
rect 356716 39030 356744 41806
rect 357636 39030 357664 41806
rect 356704 39024 356756 39030
rect 356704 38966 356756 38972
rect 357348 39024 357400 39030
rect 357348 38966 357400 38972
rect 357624 39024 357676 39030
rect 357624 38966 357676 38972
rect 356624 35866 356744 35894
rect 356336 7948 356388 7954
rect 356336 7890 356388 7896
rect 355232 3868 355284 3874
rect 355232 3810 355284 3816
rect 355968 3868 356020 3874
rect 355968 3810 356020 3816
rect 355244 480 355272 3810
rect 356348 480 356376 7890
rect 356716 6662 356744 35866
rect 357360 25566 357388 38966
rect 357348 25560 357400 25566
rect 357348 25502 357400 25508
rect 356704 6656 356756 6662
rect 356704 6598 356756 6604
rect 358648 5302 358676 41806
rect 359292 39506 359320 41806
rect 359556 39908 359608 39914
rect 359556 39850 359608 39856
rect 359464 39772 359516 39778
rect 359464 39714 359516 39720
rect 359280 39500 359332 39506
rect 359280 39442 359332 39448
rect 358728 39024 358780 39030
rect 358728 38966 358780 38972
rect 358636 5296 358688 5302
rect 358636 5238 358688 5244
rect 358740 5114 358768 38966
rect 359280 11756 359332 11762
rect 359280 11698 359332 11704
rect 358648 5086 358768 5114
rect 357532 4820 357584 4826
rect 357532 4762 357584 4768
rect 357544 480 357572 4762
rect 358648 4010 358676 5086
rect 358636 4004 358688 4010
rect 358636 3946 358688 3952
rect 358728 3936 358780 3942
rect 358728 3878 358780 3884
rect 358740 480 358768 3878
rect 359292 626 359320 11698
rect 359476 6914 359504 39714
rect 359568 8974 359596 39850
rect 360212 39030 360240 41806
rect 360200 39024 360252 39030
rect 360200 38966 360252 38972
rect 359556 8968 359608 8974
rect 359556 8910 359608 8916
rect 359384 6886 359504 6914
rect 359384 6594 359412 6886
rect 359372 6588 359424 6594
rect 359372 6530 359424 6536
rect 361120 6520 361172 6526
rect 361120 6462 361172 6468
rect 359292 598 359504 626
rect 359476 490 359504 598
rect 359752 598 359964 626
rect 359752 490 359780 598
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 462 359780 490
rect 359936 480 359964 598
rect 361132 480 361160 6462
rect 361408 5166 361436 41806
rect 361868 39778 361896 41806
rect 361856 39772 361908 39778
rect 361856 39714 361908 39720
rect 361488 39024 361540 39030
rect 361488 38966 361540 38972
rect 361396 5160 361448 5166
rect 361396 5102 361448 5108
rect 361500 3874 361528 38966
rect 361488 3868 361540 3874
rect 361488 3810 361540 3816
rect 362880 3806 362908 41806
rect 363512 39840 363564 39846
rect 363512 39782 363564 39788
rect 363524 35894 363552 39782
rect 363616 39030 363644 41806
rect 364536 39574 364564 41806
rect 364524 39568 364576 39574
rect 364524 39510 364576 39516
rect 363604 39024 363656 39030
rect 363604 38966 363656 38972
rect 364248 39024 364300 39030
rect 364248 38966 364300 38972
rect 363524 35866 363644 35894
rect 363616 14482 363644 35866
rect 363512 14476 363564 14482
rect 363512 14418 363564 14424
rect 363604 14476 363656 14482
rect 363604 14418 363656 14424
rect 362316 3800 362368 3806
rect 362316 3742 362368 3748
rect 362868 3800 362920 3806
rect 362868 3742 362920 3748
rect 362328 480 362356 3742
rect 363524 480 363552 14418
rect 364260 5234 364288 38966
rect 364616 6656 364668 6662
rect 364616 6598 364668 6604
rect 364248 5228 364300 5234
rect 364248 5170 364300 5176
rect 364628 480 364656 6598
rect 365640 3505 365668 41806
rect 366192 39030 366220 41806
rect 366180 39024 366232 39030
rect 366180 38966 366232 38972
rect 367008 39024 367060 39030
rect 367008 38966 367060 38972
rect 366916 6452 366968 6458
rect 366916 6394 366968 6400
rect 365812 3664 365864 3670
rect 365812 3606 365864 3612
rect 365626 3496 365682 3505
rect 365626 3431 365682 3440
rect 365824 480 365852 3606
rect 366928 1578 366956 6394
rect 367020 5098 367048 38966
rect 367112 38962 367140 41806
rect 367940 39030 367968 41806
rect 368768 39030 368796 41806
rect 369688 39846 369716 41806
rect 369676 39840 369728 39846
rect 369676 39782 369728 39788
rect 370412 39432 370464 39438
rect 370412 39374 370464 39380
rect 367928 39024 367980 39030
rect 367928 38966 367980 38972
rect 368388 39024 368440 39030
rect 368388 38966 368440 38972
rect 368756 39024 368808 39030
rect 368756 38966 368808 38972
rect 369768 39024 369820 39030
rect 369768 38966 369820 38972
rect 367100 38956 367152 38962
rect 367100 38898 367152 38904
rect 368296 38956 368348 38962
rect 368296 38898 368348 38904
rect 368308 11762 368336 38898
rect 368296 11756 368348 11762
rect 368296 11698 368348 11704
rect 368204 7880 368256 7886
rect 368204 7822 368256 7828
rect 367008 5092 367060 5098
rect 367008 5034 367060 5040
rect 366928 1550 367048 1578
rect 367020 480 367048 1550
rect 368216 480 368244 7822
rect 368400 3670 368428 38966
rect 369780 4962 369808 38966
rect 370424 35894 370452 39374
rect 370516 39030 370544 41806
rect 370504 39024 370556 39030
rect 370504 38966 370556 38972
rect 371148 39024 371200 39030
rect 371148 38966 371200 38972
rect 370424 35866 370544 35894
rect 370136 10328 370188 10334
rect 370136 10270 370188 10276
rect 369768 4956 369820 4962
rect 369768 4898 369820 4904
rect 369400 3732 369452 3738
rect 369400 3674 369452 3680
rect 368388 3664 368440 3670
rect 368388 3606 368440 3612
rect 369412 480 369440 3674
rect 370148 490 370176 10270
rect 370516 6934 370544 35866
rect 370504 6928 370556 6934
rect 370504 6870 370556 6876
rect 371160 3738 371188 38966
rect 371344 38962 371372 41806
rect 371332 38956 371384 38962
rect 371332 38898 371384 38904
rect 372448 26926 372476 41806
rect 373092 39030 373120 41806
rect 374012 39030 374040 41806
rect 373080 39024 373132 39030
rect 373080 38966 373132 38972
rect 373908 39024 373960 39030
rect 373908 38966 373960 38972
rect 374000 39024 374052 39030
rect 374000 38966 374052 38972
rect 372528 38956 372580 38962
rect 372528 38898 372580 38904
rect 372436 26920 372488 26926
rect 372436 26862 372488 26868
rect 371700 6384 371752 6390
rect 371700 6326 371752 6332
rect 371148 3732 371200 3738
rect 371148 3674 371200 3680
rect 370424 598 370636 626
rect 370424 490 370452 598
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 462 370452 490
rect 370608 480 370636 598
rect 371712 480 371740 6326
rect 372540 5030 372568 38898
rect 372528 5024 372580 5030
rect 372528 4966 372580 4972
rect 373920 3466 373948 38966
rect 375208 28286 375236 41806
rect 375668 39030 375696 41806
rect 375288 39024 375340 39030
rect 375288 38966 375340 38972
rect 375656 39024 375708 39030
rect 375656 38966 375708 38972
rect 375196 28280 375248 28286
rect 375196 28222 375248 28228
rect 375300 16574 375328 38966
rect 375208 16546 375328 16574
rect 374092 6316 374144 6322
rect 374092 6258 374144 6264
rect 372896 3460 372948 3466
rect 372896 3402 372948 3408
rect 373908 3460 373960 3466
rect 373908 3402 373960 3408
rect 372908 480 372936 3402
rect 374104 480 374132 6258
rect 375208 4894 375236 16546
rect 375288 6928 375340 6934
rect 375288 6870 375340 6876
rect 375196 4888 375248 4894
rect 375196 4830 375248 4836
rect 375300 480 375328 6870
rect 376588 4826 376616 41806
rect 377312 39772 377364 39778
rect 377312 39714 377364 39720
rect 376668 39024 376720 39030
rect 376668 38966 376720 38972
rect 376576 4820 376628 4826
rect 376576 4762 376628 4768
rect 376680 3534 376708 38966
rect 377324 35894 377352 39714
rect 377416 39030 377444 41806
rect 377404 39024 377456 39030
rect 377404 38966 377456 38972
rect 378048 39024 378100 39030
rect 378048 38966 378100 38972
rect 377324 35866 377444 35894
rect 377416 17270 377444 35866
rect 378060 33794 378088 38966
rect 378244 38962 378272 41806
rect 378232 38956 378284 38962
rect 378232 38898 378284 38904
rect 378048 33788 378100 33794
rect 378048 33730 378100 33736
rect 376760 17264 376812 17270
rect 376760 17206 376812 17212
rect 377404 17264 377456 17270
rect 377404 17206 377456 17212
rect 376772 16574 376800 17206
rect 376772 16546 377720 16574
rect 376484 3528 376536 3534
rect 376484 3470 376536 3476
rect 376668 3528 376720 3534
rect 376668 3470 376720 3476
rect 376496 480 376524 3470
rect 377692 480 377720 16546
rect 378876 7812 378928 7818
rect 378876 7754 378928 7760
rect 378888 480 378916 7754
rect 379348 6866 379376 41806
rect 379992 39438 380020 41806
rect 379980 39432 380032 39438
rect 379980 39374 380032 39380
rect 379428 38956 379480 38962
rect 379428 38898 379480 38904
rect 379336 6860 379388 6866
rect 379336 6802 379388 6808
rect 379440 3369 379468 38898
rect 380820 3602 380848 41806
rect 381544 39840 381596 39846
rect 381544 39782 381596 39788
rect 381556 18630 381584 39782
rect 381740 38894 381768 41806
rect 382568 39030 382596 41806
rect 382556 39024 382608 39030
rect 382556 38966 382608 38972
rect 383476 39024 383528 39030
rect 383476 38966 383528 38972
rect 381728 38888 381780 38894
rect 381728 38830 381780 38836
rect 382188 38888 382240 38894
rect 382188 38830 382240 38836
rect 380900 18624 380952 18630
rect 380900 18566 380952 18572
rect 381544 18624 381596 18630
rect 381544 18566 381596 18572
rect 380912 16574 380940 18566
rect 380912 16546 381216 16574
rect 379980 3596 380032 3602
rect 379980 3538 380032 3544
rect 380808 3596 380860 3602
rect 380808 3538 380860 3544
rect 379426 3360 379482 3369
rect 379426 3295 379482 3304
rect 379992 480 380020 3538
rect 381188 480 381216 16546
rect 382200 6118 382228 38830
rect 383488 31074 383516 38966
rect 383476 31068 383528 31074
rect 383476 31010 383528 31016
rect 382372 7744 382424 7750
rect 382372 7686 382424 7692
rect 382188 6112 382240 6118
rect 382188 6054 382240 6060
rect 382384 480 382412 7686
rect 383580 2938 383608 41806
rect 384316 39030 384344 41806
rect 384304 39024 384356 39030
rect 384304 38966 384356 38972
rect 384948 39024 385000 39030
rect 384948 38966 385000 38972
rect 384960 6798 384988 38966
rect 385144 38418 385172 41806
rect 385132 38412 385184 38418
rect 385132 38354 385184 38360
rect 385960 7676 386012 7682
rect 385960 7618 386012 7624
rect 384948 6792 385000 6798
rect 384948 6734 385000 6740
rect 384764 6248 384816 6254
rect 384764 6190 384816 6196
rect 383580 2910 383700 2938
rect 383672 2854 383700 2910
rect 383568 2848 383620 2854
rect 383568 2790 383620 2796
rect 383660 2848 383712 2854
rect 383660 2790 383712 2796
rect 383580 480 383608 2790
rect 384776 480 384804 6190
rect 385972 480 386000 7618
rect 386248 3777 386276 41806
rect 386892 38826 386920 41806
rect 387720 39302 387748 41806
rect 388444 39432 388496 39438
rect 388444 39374 388496 39380
rect 387708 39296 387760 39302
rect 387708 39238 387760 39244
rect 386880 38820 386932 38826
rect 386880 38762 386932 38768
rect 387708 38820 387760 38826
rect 387708 38762 387760 38768
rect 387720 6662 387748 38762
rect 388456 21418 388484 39374
rect 388640 39030 388668 41806
rect 389468 39030 389496 41806
rect 388628 39024 388680 39030
rect 388628 38966 388680 38972
rect 389088 39024 389140 39030
rect 389088 38966 389140 38972
rect 389456 39024 389508 39030
rect 389456 38966 389508 38972
rect 387800 21412 387852 21418
rect 387800 21354 387852 21360
rect 388444 21412 388496 21418
rect 388444 21354 388496 21360
rect 387708 6656 387760 6662
rect 387708 6598 387760 6604
rect 387156 6180 387208 6186
rect 387156 6122 387208 6128
rect 386234 3768 386290 3777
rect 386234 3703 386290 3712
rect 387168 480 387196 6122
rect 387812 490 387840 21354
rect 389100 3641 389128 38966
rect 390388 9042 390416 41806
rect 391216 39982 391244 41806
rect 391204 39976 391256 39982
rect 391204 39918 391256 39924
rect 392044 39166 392072 41806
rect 392032 39160 392084 39166
rect 392032 39102 392084 39108
rect 390468 39024 390520 39030
rect 390468 38966 390520 38972
rect 390376 9036 390428 9042
rect 390376 8978 390428 8984
rect 389456 8968 389508 8974
rect 389456 8910 389508 8916
rect 389086 3632 389142 3641
rect 389086 3567 389142 3576
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 8910
rect 390480 6730 390508 38966
rect 391940 22772 391992 22778
rect 391940 22714 391992 22720
rect 391952 16574 391980 22714
rect 391952 16546 392624 16574
rect 390468 6724 390520 6730
rect 390468 6666 390520 6672
rect 390652 6588 390704 6594
rect 390652 6530 390704 6536
rect 390664 480 390692 6530
rect 391848 6044 391900 6050
rect 391848 5986 391900 5992
rect 391860 480 391888 5986
rect 392596 490 392624 16546
rect 393240 6526 393268 41806
rect 393792 40050 393820 41806
rect 393780 40044 393832 40050
rect 393780 39986 393832 39992
rect 393964 39364 394016 39370
rect 393964 39306 394016 39312
rect 393228 6520 393280 6526
rect 393228 6462 393280 6468
rect 393976 5574 394004 39306
rect 394620 8158 394648 41806
rect 395344 39636 395396 39642
rect 395344 39578 395396 39584
rect 394608 8152 394660 8158
rect 394608 8094 394660 8100
rect 395356 7750 395384 39578
rect 395540 39030 395568 41806
rect 396368 39030 396396 41806
rect 396724 39704 396776 39710
rect 396724 39646 396776 39652
rect 395528 39024 395580 39030
rect 395528 38966 395580 38972
rect 395988 39024 396040 39030
rect 395988 38966 396040 38972
rect 396356 39024 396408 39030
rect 396356 38966 396408 38972
rect 395344 7744 395396 7750
rect 395344 7686 395396 7692
rect 396000 6594 396028 38966
rect 396736 7682 396764 39646
rect 397196 39642 397224 41806
rect 397184 39636 397236 39642
rect 397184 39578 397236 39584
rect 398116 39030 398144 41806
rect 398944 39846 398972 41806
rect 398932 39840 398984 39846
rect 398932 39782 398984 39788
rect 397368 39024 397420 39030
rect 397368 38966 397420 38972
rect 398104 39024 398156 39030
rect 398104 38966 398156 38972
rect 398748 39024 398800 39030
rect 398748 38966 398800 38972
rect 397380 35290 397408 38966
rect 397368 35284 397420 35290
rect 397368 35226 397420 35232
rect 396724 7676 396776 7682
rect 396724 7618 396776 7624
rect 395988 6588 396040 6594
rect 395988 6530 396040 6536
rect 398760 6390 398788 38966
rect 398840 37936 398892 37942
rect 398840 37878 398892 37884
rect 398748 6384 398800 6390
rect 398748 6326 398800 6332
rect 393964 5568 394016 5574
rect 393964 5510 394016 5516
rect 396540 5568 396592 5574
rect 396540 5510 396592 5516
rect 395344 4276 395396 4282
rect 395344 4218 395396 4224
rect 394240 2916 394292 2922
rect 394240 2858 394292 2864
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 2858
rect 395356 480 395384 4218
rect 396552 480 396580 5510
rect 398852 3058 398880 37878
rect 400140 8090 400168 41806
rect 400692 39030 400720 41806
rect 401428 41806 401502 41834
rect 402302 41834 402330 42092
rect 403222 41834 403250 42092
rect 404050 41834 404078 42092
rect 404970 41834 404998 42092
rect 405798 41834 405826 42092
rect 406626 41834 406654 42092
rect 407546 41834 407574 42092
rect 408374 41834 408402 42092
rect 402302 41806 402376 41834
rect 403222 41806 403296 41834
rect 404050 41806 404124 41834
rect 404970 41806 405044 41834
rect 405798 41806 405872 41834
rect 406626 41806 406700 41834
rect 407546 41806 407620 41834
rect 400680 39024 400732 39030
rect 400680 38966 400732 38972
rect 401428 22778 401456 41806
rect 402348 39778 402376 41806
rect 402336 39772 402388 39778
rect 402336 39714 402388 39720
rect 403268 39030 403296 41806
rect 404096 39710 404124 41806
rect 404084 39704 404136 39710
rect 404084 39646 404136 39652
rect 405016 39234 405044 41806
rect 405004 39228 405056 39234
rect 405004 39170 405056 39176
rect 405844 39030 405872 41806
rect 401508 39024 401560 39030
rect 401508 38966 401560 38972
rect 403256 39024 403308 39030
rect 403256 38966 403308 38972
rect 404268 39024 404320 39030
rect 404268 38966 404320 38972
rect 405832 39024 405884 39030
rect 405832 38966 405884 38972
rect 401416 22772 401468 22778
rect 401416 22714 401468 22720
rect 400128 8084 400180 8090
rect 400128 8026 400180 8032
rect 401520 6458 401548 38966
rect 403624 15904 403676 15910
rect 403624 15846 403676 15852
rect 401508 6452 401560 6458
rect 401508 6394 401560 6400
rect 402520 4412 402572 4418
rect 402520 4354 402572 4360
rect 398932 4344 398984 4350
rect 398932 4286 398984 4292
rect 398840 3052 398892 3058
rect 398840 2994 398892 3000
rect 397736 2984 397788 2990
rect 397736 2926 397788 2932
rect 397748 480 397776 2926
rect 398944 480 398972 4286
rect 400128 3052 400180 3058
rect 400128 2994 400180 3000
rect 400140 480 400168 2994
rect 401324 2984 401376 2990
rect 401324 2926 401376 2932
rect 401336 480 401364 2926
rect 402532 480 402560 4354
rect 403636 480 403664 15846
rect 404280 6322 404308 38966
rect 406672 36922 406700 41806
rect 407028 39024 407080 39030
rect 407028 38966 407080 38972
rect 406660 36916 406712 36922
rect 406660 36858 406712 36864
rect 404268 6316 404320 6322
rect 404268 6258 404320 6264
rect 407040 6254 407068 38966
rect 407592 38350 407620 41806
rect 408328 41806 408402 41834
rect 409202 41834 409230 42092
rect 410122 41834 410150 42092
rect 410950 41834 410978 42092
rect 411778 41834 411806 42092
rect 412698 41834 412726 42092
rect 413526 41834 413554 42092
rect 414354 41834 414382 42092
rect 415274 41834 415302 42092
rect 416102 41834 416130 42092
rect 417022 41834 417050 42092
rect 417850 41834 417878 42092
rect 418678 41834 418706 42092
rect 419598 41834 419626 42092
rect 420426 41834 420454 42092
rect 421254 41834 421282 42092
rect 422174 41834 422202 42092
rect 409202 41806 409276 41834
rect 410122 41806 410196 41834
rect 410950 41806 411208 41834
rect 411778 41806 411852 41834
rect 412698 41806 412772 41834
rect 413526 41806 413876 41834
rect 414354 41806 414428 41834
rect 415274 41806 415348 41834
rect 416102 41806 416176 41834
rect 417022 41806 417096 41834
rect 417850 41806 418108 41834
rect 418678 41806 418752 41834
rect 419598 41806 419672 41834
rect 420426 41806 420776 41834
rect 421254 41806 421328 41834
rect 407580 38344 407632 38350
rect 407580 38286 407632 38292
rect 407212 29640 407264 29646
rect 407212 29582 407264 29588
rect 407028 6248 407080 6254
rect 407028 6190 407080 6196
rect 406016 4548 406068 4554
rect 406016 4490 406068 4496
rect 404820 3120 404872 3126
rect 404820 3062 404872 3068
rect 404832 480 404860 3062
rect 406028 480 406056 4490
rect 407224 480 407252 29582
rect 408328 6186 408356 41806
rect 409248 39438 409276 41806
rect 409236 39432 409288 39438
rect 409236 39374 409288 39380
rect 410168 39098 410196 41806
rect 410156 39092 410208 39098
rect 410156 39034 410208 39040
rect 409880 24132 409932 24138
rect 409880 24074 409932 24080
rect 409892 16574 409920 24074
rect 409892 16546 410840 16574
rect 408316 6180 408368 6186
rect 408316 6122 408368 6128
rect 409604 4480 409656 4486
rect 409604 4422 409656 4428
rect 408408 3188 408460 3194
rect 408408 3130 408460 3136
rect 408420 480 408448 3130
rect 409616 480 409644 4422
rect 410812 480 410840 16546
rect 411180 8974 411208 41806
rect 411824 36854 411852 41806
rect 411904 39500 411956 39506
rect 411904 39442 411956 39448
rect 411812 36848 411864 36854
rect 411812 36790 411864 36796
rect 411168 8968 411220 8974
rect 411168 8910 411220 8916
rect 411916 8294 411944 39442
rect 412744 38282 412772 41806
rect 413284 39568 413336 39574
rect 413284 39510 413336 39516
rect 412732 38276 412784 38282
rect 412732 38218 412784 38224
rect 411904 8288 411956 8294
rect 411904 8230 411956 8236
rect 413296 8226 413324 39510
rect 413284 8220 413336 8226
rect 413284 8162 413336 8168
rect 413848 8022 413876 41806
rect 414400 39574 414428 41806
rect 414388 39568 414440 39574
rect 414388 39510 414440 39516
rect 414296 13116 414348 13122
rect 414296 13058 414348 13064
rect 413836 8016 413888 8022
rect 413836 7958 413888 7964
rect 413100 4616 413152 4622
rect 413100 4558 413152 4564
rect 411904 3256 411956 3262
rect 411904 3198 411956 3204
rect 411916 480 411944 3198
rect 413112 480 413140 4558
rect 414308 480 414336 13058
rect 415320 4282 415348 41806
rect 416148 39370 416176 41806
rect 416136 39364 416188 39370
rect 416136 39306 416188 39312
rect 417068 39030 417096 41806
rect 417056 39024 417108 39030
rect 417056 38966 417108 38972
rect 417976 39024 418028 39030
rect 417976 38966 418028 38972
rect 417988 35222 418016 38966
rect 417976 35216 418028 35222
rect 417976 35158 418028 35164
rect 417884 7744 417936 7750
rect 417884 7686 417936 7692
rect 416688 4684 416740 4690
rect 416688 4626 416740 4632
rect 415308 4276 415360 4282
rect 415308 4218 415360 4224
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 415504 480 415532 3334
rect 416700 480 416728 4626
rect 417896 480 417924 7686
rect 418080 4350 418108 41806
rect 418724 39030 418752 41806
rect 419644 39030 419672 41806
rect 418712 39024 418764 39030
rect 418712 38966 418764 38972
rect 419448 39024 419500 39030
rect 419448 38966 419500 38972
rect 419632 39024 419684 39030
rect 419632 38966 419684 38972
rect 419460 7954 419488 38966
rect 419448 7948 419500 7954
rect 419448 7890 419500 7896
rect 420184 4752 420236 4758
rect 420184 4694 420236 4700
rect 418068 4344 418120 4350
rect 418068 4286 418120 4292
rect 418988 3324 419040 3330
rect 418988 3266 419040 3272
rect 419000 480 419028 3266
rect 420196 480 420224 4694
rect 420748 4418 420776 41806
rect 420828 39024 420880 39030
rect 420828 38966 420880 38972
rect 420736 4412 420788 4418
rect 420736 4354 420788 4360
rect 420840 2922 420868 38966
rect 421300 38214 421328 41806
rect 422128 41806 422202 41834
rect 423002 41834 423030 42092
rect 423830 41834 423858 42092
rect 424750 41834 424778 42092
rect 425578 41834 425606 42092
rect 426498 41834 426526 42092
rect 427326 41834 427354 42092
rect 428154 41834 428182 42092
rect 429074 41834 429102 42092
rect 423002 41806 423076 41834
rect 423830 41806 423904 41834
rect 424750 41806 425008 41834
rect 425578 41806 425652 41834
rect 426498 41806 426572 41834
rect 427326 41806 427768 41834
rect 428154 41806 428228 41834
rect 421288 38208 421340 38214
rect 421288 38150 421340 38156
rect 420920 14476 420972 14482
rect 420920 14418 420972 14424
rect 420828 2916 420880 2922
rect 420828 2858 420880 2864
rect 420932 490 420960 14418
rect 422128 3058 422156 41806
rect 423048 39030 423076 41806
rect 423876 39370 423904 41806
rect 423864 39364 423916 39370
rect 423864 39306 423916 39312
rect 423036 39024 423088 39030
rect 423036 38966 423088 38972
rect 423588 39024 423640 39030
rect 423588 38966 423640 38972
rect 423600 4554 423628 38966
rect 424876 7676 424928 7682
rect 424876 7618 424928 7624
rect 423772 5432 423824 5438
rect 423772 5374 423824 5380
rect 423588 4548 423640 4554
rect 423588 4490 423640 4496
rect 422576 4140 422628 4146
rect 422576 4082 422628 4088
rect 422116 3052 422168 3058
rect 422116 2994 422168 3000
rect 421208 598 421420 626
rect 421208 490 421236 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 462 421236 490
rect 421392 480 421420 598
rect 422588 480 422616 4082
rect 423784 480 423812 5374
rect 424784 4140 424836 4146
rect 424784 4082 424836 4088
rect 424796 2990 424824 4082
rect 424888 3482 424916 7618
rect 424980 4146 425008 41806
rect 425624 39030 425652 41806
rect 425612 39024 425664 39030
rect 425612 38966 425664 38972
rect 426348 39024 426400 39030
rect 426348 38966 426400 38972
rect 426360 4486 426388 38966
rect 426544 38962 426572 41806
rect 426532 38956 426584 38962
rect 426532 38898 426584 38904
rect 427268 5500 427320 5506
rect 427268 5442 427320 5448
rect 426348 4480 426400 4486
rect 426348 4422 426400 4428
rect 424968 4140 425020 4146
rect 424968 4082 425020 4088
rect 426164 4072 426216 4078
rect 426164 4014 426216 4020
rect 424888 3454 425008 3482
rect 424784 2984 424836 2990
rect 424784 2926 424836 2932
rect 424980 480 425008 3454
rect 426176 480 426204 4014
rect 427280 480 427308 5442
rect 427740 3194 427768 41806
rect 428200 39030 428228 41806
rect 429028 41806 429102 41834
rect 429902 41834 429930 42092
rect 430730 41834 430758 42092
rect 431650 41834 431678 42092
rect 432478 41834 432506 42092
rect 433306 41834 433334 42092
rect 434226 41834 434254 42092
rect 435054 41834 435082 42092
rect 435974 41834 436002 42092
rect 429902 41806 429976 41834
rect 430730 41806 430804 41834
rect 431650 41806 431816 41834
rect 432478 41806 432552 41834
rect 433306 41806 433380 41834
rect 434226 41806 434300 41834
rect 435054 41806 435128 41834
rect 428188 39024 428240 39030
rect 428188 38966 428240 38972
rect 429028 7750 429056 41806
rect 429948 39030 429976 41806
rect 430776 39030 430804 41806
rect 429108 39024 429160 39030
rect 429108 38966 429160 38972
rect 429936 39024 429988 39030
rect 429936 38966 429988 38972
rect 430488 39024 430540 39030
rect 430488 38966 430540 38972
rect 430764 39024 430816 39030
rect 430764 38966 430816 38972
rect 429016 7744 429068 7750
rect 429016 7686 429068 7692
rect 428464 7608 428516 7614
rect 428464 7550 428516 7556
rect 427728 3188 427780 3194
rect 427728 3130 427780 3136
rect 428476 480 428504 7550
rect 429120 4622 429148 38966
rect 429844 38956 429896 38962
rect 429844 38898 429896 38904
rect 429856 7886 429884 38898
rect 429844 7880 429896 7886
rect 429844 7822 429896 7828
rect 429108 4616 429160 4622
rect 429108 4558 429160 4564
rect 429660 4004 429712 4010
rect 429660 3946 429712 3952
rect 429672 480 429700 3946
rect 430500 3126 430528 38966
rect 431788 7818 431816 41806
rect 432524 39030 432552 41806
rect 433352 39030 433380 41806
rect 434272 39370 434300 41806
rect 434260 39364 434312 39370
rect 434260 39306 434312 39312
rect 435100 39030 435128 41806
rect 435928 41806 436002 41834
rect 436802 41834 436830 42092
rect 437630 41834 437658 42092
rect 438550 41834 438578 42092
rect 439378 41834 439406 42092
rect 440206 41834 440234 42092
rect 441126 41834 441154 42092
rect 441954 41834 441982 42092
rect 442782 41834 442810 42092
rect 443702 41834 443730 42092
rect 444530 41834 444558 42092
rect 445358 41834 445386 42092
rect 446278 41834 446306 42092
rect 447106 41834 447134 42092
rect 448026 41834 448054 42092
rect 448854 41834 448882 42092
rect 449682 41834 449710 42092
rect 450602 41834 450630 42092
rect 451430 41834 451458 42092
rect 452258 41834 452286 42092
rect 453178 41834 453206 42092
rect 454006 41834 454034 42092
rect 454834 41834 454862 42092
rect 455754 41834 455782 42092
rect 456582 41834 456610 42092
rect 457502 41834 457530 42092
rect 458330 41834 458358 42092
rect 459158 41834 459186 42092
rect 460078 41834 460106 42092
rect 460906 41834 460934 42092
rect 461734 41834 461762 42092
rect 462654 41834 462682 42092
rect 463482 41834 463510 42092
rect 464310 41834 464338 42092
rect 465230 41834 465258 42092
rect 466058 41834 466086 42092
rect 436802 41806 436876 41834
rect 437630 41806 437704 41834
rect 438550 41806 438716 41834
rect 439378 41806 439452 41834
rect 440206 41806 440280 41834
rect 441126 41806 441476 41834
rect 441954 41806 442028 41834
rect 442782 41806 442948 41834
rect 443702 41806 443776 41834
rect 444530 41806 444604 41834
rect 445358 41806 445616 41834
rect 446278 41806 446352 41834
rect 447106 41806 447180 41834
rect 448026 41806 448468 41834
rect 448854 41806 448928 41834
rect 449682 41806 449756 41834
rect 450602 41806 450676 41834
rect 451430 41806 451504 41834
rect 452258 41806 452332 41834
rect 453178 41806 453252 41834
rect 454006 41806 454080 41834
rect 454834 41806 454908 41834
rect 455754 41806 455828 41834
rect 456582 41806 456656 41834
rect 457502 41806 457576 41834
rect 458330 41806 458404 41834
rect 459158 41806 459416 41834
rect 460078 41806 460152 41834
rect 460906 41806 460980 41834
rect 461734 41806 462176 41834
rect 462654 41806 462728 41834
rect 463482 41806 463648 41834
rect 464310 41806 464384 41834
rect 465230 41806 465304 41834
rect 466058 41806 466408 41834
rect 431868 39024 431920 39030
rect 431868 38966 431920 38972
rect 432512 39024 432564 39030
rect 432512 38966 432564 38972
rect 433248 39024 433300 39030
rect 433248 38966 433300 38972
rect 433340 39024 433392 39030
rect 433340 38966 433392 38972
rect 434628 39024 434680 39030
rect 434628 38966 434680 38972
rect 435088 39024 435140 39030
rect 435088 38966 435140 38972
rect 431776 7812 431828 7818
rect 431776 7754 431828 7760
rect 430856 5364 430908 5370
rect 430856 5306 430908 5312
rect 430488 3120 430540 3126
rect 430488 3062 430540 3068
rect 430868 480 430896 5306
rect 431880 4690 431908 38966
rect 432052 25560 432104 25566
rect 432052 25502 432104 25508
rect 431868 4684 431920 4690
rect 431868 4626 431920 4632
rect 432064 480 432092 25502
rect 433260 6914 433288 38966
rect 433168 6886 433288 6914
rect 433168 3262 433196 6886
rect 434444 5296 434496 5302
rect 434444 5238 434496 5244
rect 433248 3936 433300 3942
rect 433248 3878 433300 3884
rect 433156 3256 433208 3262
rect 433156 3198 433208 3204
rect 433260 480 433288 3878
rect 434456 480 434484 5238
rect 434640 4758 434668 38966
rect 435548 8288 435600 8294
rect 435548 8230 435600 8236
rect 434628 4752 434680 4758
rect 434628 4694 434680 4700
rect 435560 480 435588 8230
rect 435928 5506 435956 41806
rect 436848 39030 436876 41806
rect 437296 39364 437348 39370
rect 437296 39306 437348 39312
rect 436008 39024 436060 39030
rect 436008 38966 436060 38972
rect 436836 39024 436888 39030
rect 436836 38966 436888 38972
rect 435916 5500 435968 5506
rect 435916 5442 435968 5448
rect 436020 3330 436048 38966
rect 437308 38146 437336 39306
rect 437676 39030 437704 41806
rect 437388 39024 437440 39030
rect 437388 38966 437440 38972
rect 437664 39024 437716 39030
rect 437664 38966 437716 38972
rect 437296 38140 437348 38146
rect 437296 38082 437348 38088
rect 437400 7682 437428 38966
rect 437388 7676 437440 7682
rect 437388 7618 437440 7624
rect 438688 5438 438716 41806
rect 438768 39024 438820 39030
rect 438768 38966 438820 38972
rect 438676 5432 438728 5438
rect 438676 5374 438728 5380
rect 437940 5160 437992 5166
rect 437940 5102 437992 5108
rect 436744 3868 436796 3874
rect 436744 3810 436796 3816
rect 436008 3324 436060 3330
rect 436008 3266 436060 3272
rect 436756 480 436784 3810
rect 437952 480 437980 5102
rect 438780 3398 438808 38966
rect 439424 38758 439452 41806
rect 440252 39030 440280 41806
rect 440240 39024 440292 39030
rect 440240 38966 440292 38972
rect 439412 38752 439464 38758
rect 439412 38694 439464 38700
rect 440148 38752 440200 38758
rect 440148 38694 440200 38700
rect 438860 17264 438912 17270
rect 438860 17206 438912 17212
rect 438872 16574 438900 17206
rect 438872 16546 439176 16574
rect 438768 3392 438820 3398
rect 438768 3334 438820 3340
rect 439148 480 439176 16546
rect 440160 7614 440188 38694
rect 441344 8288 441396 8294
rect 441344 8230 441396 8236
rect 440148 7608 440200 7614
rect 440148 7550 440200 7556
rect 441356 4146 441384 8230
rect 441448 5302 441476 41806
rect 442000 39370 442028 41806
rect 441988 39364 442040 39370
rect 441988 39306 442040 39312
rect 441528 39024 441580 39030
rect 441528 38966 441580 38972
rect 441540 8294 441568 38966
rect 441528 8288 441580 8294
rect 441528 8230 441580 8236
rect 442632 8220 442684 8226
rect 442632 8162 442684 8168
rect 441436 5296 441488 5302
rect 441436 5238 441488 5244
rect 441528 5228 441580 5234
rect 441528 5170 441580 5176
rect 441344 4140 441396 4146
rect 441344 4082 441396 4088
rect 440332 3800 440384 3806
rect 440332 3742 440384 3748
rect 440344 480 440372 3742
rect 441540 480 441568 5170
rect 442644 480 442672 8162
rect 442920 4078 442948 41806
rect 443748 39030 443776 41806
rect 444196 39364 444248 39370
rect 444196 39306 444248 39312
rect 443736 39024 443788 39030
rect 443736 38966 443788 38972
rect 444208 38078 444236 39306
rect 444288 39024 444340 39030
rect 444288 38966 444340 38972
rect 444196 38072 444248 38078
rect 444196 38014 444248 38020
rect 444300 5370 444328 38966
rect 444576 38010 444604 41806
rect 444564 38004 444616 38010
rect 444564 37946 444616 37952
rect 444288 5364 444340 5370
rect 444288 5306 444340 5312
rect 445024 5092 445076 5098
rect 445024 5034 445076 5040
rect 442908 4072 442960 4078
rect 442908 4014 442960 4020
rect 443826 3496 443882 3505
rect 443826 3431 443882 3440
rect 443840 480 443868 3431
rect 445036 480 445064 5034
rect 445588 3942 445616 41806
rect 446324 39030 446352 41806
rect 446312 39024 446364 39030
rect 446312 38966 446364 38972
rect 447048 39024 447100 39030
rect 447048 38966 447100 38972
rect 445760 11756 445812 11762
rect 445760 11698 445812 11704
rect 445576 3936 445628 3942
rect 445576 3878 445628 3884
rect 445772 490 445800 11698
rect 447060 5166 447088 38966
rect 447152 36786 447180 41806
rect 447140 36780 447192 36786
rect 447140 36722 447192 36728
rect 447048 5160 447100 5166
rect 447048 5102 447100 5108
rect 448440 4010 448468 41806
rect 448900 39030 448928 41806
rect 448888 39024 448940 39030
rect 448888 38966 448940 38972
rect 449728 36718 449756 41806
rect 450648 39030 450676 41806
rect 451476 39030 451504 41806
rect 449808 39024 449860 39030
rect 449808 38966 449860 38972
rect 450636 39024 450688 39030
rect 450636 38966 450688 38972
rect 451188 39024 451240 39030
rect 451188 38966 451240 38972
rect 451464 39024 451516 39030
rect 451464 38966 451516 38972
rect 449716 36712 449768 36718
rect 449716 36654 449768 36660
rect 448520 18624 448572 18630
rect 448520 18566 448572 18572
rect 448428 4004 448480 4010
rect 448428 3946 448480 3952
rect 448532 3670 448560 18566
rect 449820 5234 449848 38966
rect 449808 5228 449860 5234
rect 449808 5170 449860 5176
rect 448612 4956 448664 4962
rect 448612 4898 448664 4904
rect 447416 3664 447468 3670
rect 447416 3606 447468 3612
rect 448520 3664 448572 3670
rect 448520 3606 448572 3612
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 3606
rect 448624 480 448652 4898
rect 451200 3874 451228 38966
rect 452304 37942 452332 41806
rect 453224 39030 453252 41806
rect 454052 39030 454080 41806
rect 452476 39024 452528 39030
rect 452476 38966 452528 38972
rect 453212 39024 453264 39030
rect 453212 38966 453264 38972
rect 453948 39024 454000 39030
rect 453948 38966 454000 38972
rect 454040 39024 454092 39030
rect 454040 38966 454092 38972
rect 452292 37936 452344 37942
rect 452292 37878 452344 37884
rect 452488 5098 452516 38966
rect 452660 26920 452712 26926
rect 452660 26862 452712 26868
rect 452672 16574 452700 26862
rect 452672 16546 453344 16574
rect 452476 5092 452528 5098
rect 452476 5034 452528 5040
rect 452108 5024 452160 5030
rect 452108 4966 452160 4972
rect 451188 3868 451240 3874
rect 451188 3810 451240 3816
rect 450912 3732 450964 3738
rect 450912 3674 450964 3680
rect 449808 3664 449860 3670
rect 449808 3606 449860 3612
rect 449820 480 449848 3606
rect 450924 480 450952 3674
rect 452120 480 452148 4966
rect 453316 480 453344 16546
rect 453960 3806 453988 38966
rect 454880 36650 454908 41806
rect 455800 39030 455828 41806
rect 455328 39024 455380 39030
rect 455328 38966 455380 38972
rect 455788 39024 455840 39030
rect 455788 38966 455840 38972
rect 454868 36644 454920 36650
rect 454868 36586 454920 36592
rect 455340 5030 455368 38966
rect 455328 5024 455380 5030
rect 455328 4966 455380 4972
rect 456628 4962 456656 41806
rect 457548 39030 457576 41806
rect 458376 39030 458404 41806
rect 456708 39024 456760 39030
rect 456708 38966 456760 38972
rect 457536 39024 457588 39030
rect 457536 38966 457588 38972
rect 458088 39024 458140 39030
rect 458088 38966 458140 38972
rect 458364 39024 458416 39030
rect 458364 38966 458416 38972
rect 456616 4956 456668 4962
rect 456616 4898 456668 4904
rect 455696 4888 455748 4894
rect 455696 4830 455748 4836
rect 453948 3800 454000 3806
rect 453948 3742 454000 3748
rect 454500 3460 454552 3466
rect 454500 3402 454552 3408
rect 454512 480 454540 3402
rect 455708 480 455736 4830
rect 456720 3738 456748 38966
rect 456892 28280 456944 28286
rect 456892 28222 456944 28228
rect 456708 3732 456760 3738
rect 456708 3674 456760 3680
rect 456904 480 456932 28222
rect 458100 10334 458128 38966
rect 458088 10328 458140 10334
rect 458088 10270 458140 10276
rect 459388 4826 459416 41806
rect 459468 39024 459520 39030
rect 459468 38966 459520 38972
rect 459192 4820 459244 4826
rect 459192 4762 459244 4768
rect 459376 4820 459428 4826
rect 459376 4762 459428 4768
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 458100 480 458128 3470
rect 459204 480 459232 4762
rect 459480 3670 459508 38966
rect 460124 36582 460152 41806
rect 460952 39030 460980 41806
rect 460940 39024 460992 39030
rect 460940 38966 460992 38972
rect 460112 36576 460164 36582
rect 460112 36518 460164 36524
rect 459560 33788 459612 33794
rect 459560 33730 459612 33736
rect 459572 16574 459600 33730
rect 459572 16546 459968 16574
rect 459468 3664 459520 3670
rect 459468 3606 459520 3612
rect 459940 490 459968 16546
rect 462148 4894 462176 41806
rect 462700 39370 462728 41806
rect 462688 39364 462740 39370
rect 462688 39306 462740 39312
rect 462228 39024 462280 39030
rect 462228 38966 462280 38972
rect 462136 4888 462188 4894
rect 462136 4830 462188 4836
rect 462240 3534 462268 38966
rect 462780 6860 462832 6866
rect 462780 6802 462832 6808
rect 462228 3528 462280 3534
rect 462228 3470 462280 3476
rect 461582 3360 461638 3369
rect 461582 3295 461638 3304
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 3295
rect 462792 480 462820 6802
rect 463620 3466 463648 41806
rect 464356 38962 464384 41806
rect 465276 39030 465304 41806
rect 465264 39024 465316 39030
rect 465264 38966 465316 38972
rect 466276 39024 466328 39030
rect 466276 38966 466328 38972
rect 464344 38956 464396 38962
rect 464344 38898 464396 38904
rect 464988 38956 465040 38962
rect 464988 38898 465040 38904
rect 463700 21412 463752 21418
rect 463700 21354 463752 21360
rect 463712 16574 463740 21354
rect 463712 16546 464016 16574
rect 463608 3460 463660 3466
rect 463608 3402 463660 3408
rect 463988 480 464016 16546
rect 465000 3505 465028 38898
rect 466288 6914 466316 38966
rect 466196 6886 466316 6914
rect 466196 3602 466224 6886
rect 466276 6112 466328 6118
rect 466276 6054 466328 6060
rect 465172 3596 465224 3602
rect 465172 3538 465224 3544
rect 466184 3596 466236 3602
rect 466184 3538 466236 3544
rect 464986 3496 465042 3505
rect 464986 3431 465042 3440
rect 465184 480 465212 3538
rect 466288 480 466316 6054
rect 466380 3369 466408 41806
rect 481640 40044 481692 40050
rect 481640 39986 481692 39992
rect 478880 39976 478932 39982
rect 478880 39918 478932 39924
rect 473360 39296 473412 39302
rect 473360 39238 473412 39244
rect 467104 39092 467156 39098
rect 467104 39034 467156 39040
rect 466460 31068 466512 31074
rect 466460 31010 466512 31016
rect 466472 6914 466500 31010
rect 467116 16574 467144 39034
rect 470600 38412 470652 38418
rect 470600 38354 470652 38360
rect 467116 16546 467236 16574
rect 466472 6886 467144 6914
rect 467116 3482 467144 6886
rect 467208 6866 467236 16546
rect 467196 6860 467248 6866
rect 467196 6802 467248 6808
rect 469864 6792 469916 6798
rect 469864 6734 469916 6740
rect 467116 3454 467512 3482
rect 466366 3360 466422 3369
rect 466366 3295 466422 3304
rect 467484 480 467512 3454
rect 468668 2848 468720 2854
rect 468668 2790 468720 2796
rect 468680 480 468708 2790
rect 469876 480 469904 6734
rect 470612 490 470640 38354
rect 473372 16574 473400 39238
rect 475384 39160 475436 39166
rect 475384 39102 475436 39108
rect 473372 16546 474136 16574
rect 473452 6656 473504 6662
rect 473452 6598 473504 6604
rect 472254 3768 472310 3777
rect 472254 3703 472310 3712
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 3703
rect 473464 480 473492 6598
rect 474108 490 474136 16546
rect 475396 5574 475424 39102
rect 478144 9036 478196 9042
rect 478144 8978 478196 8984
rect 476948 6724 477000 6730
rect 476948 6666 477000 6672
rect 475384 5568 475436 5574
rect 475384 5510 475436 5516
rect 475750 3632 475806 3641
rect 475750 3567 475806 3576
rect 474384 598 474596 626
rect 474384 490 474412 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 462 474412 490
rect 474568 480 474596 598
rect 475764 480 475792 3567
rect 476960 480 476988 6666
rect 478156 480 478184 8978
rect 478892 490 478920 39918
rect 481652 16574 481680 39986
rect 486424 39908 486476 39914
rect 486424 39850 486476 39856
rect 485780 35284 485832 35290
rect 485780 35226 485832 35232
rect 485792 16574 485820 35226
rect 481652 16546 482416 16574
rect 485792 16546 486372 16574
rect 481732 6520 481784 6526
rect 481732 6462 481784 6468
rect 480536 5568 480588 5574
rect 480536 5510 480588 5516
rect 479168 598 479380 626
rect 479168 490 479196 598
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 478892 462 479196 490
rect 479352 480 479380 598
rect 480548 480 480576 5510
rect 481744 480 481772 6462
rect 482388 490 482416 16546
rect 484032 8152 484084 8158
rect 484032 8094 484084 8100
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 8094
rect 485228 6588 485280 6594
rect 485228 6530 485280 6536
rect 485240 480 485268 6530
rect 486344 3482 486372 16546
rect 486436 5574 486464 39850
rect 489920 39840 489972 39846
rect 489920 39782 489972 39788
rect 489184 39228 489236 39234
rect 489184 39170 489236 39176
rect 489196 6390 489224 39170
rect 488816 6384 488868 6390
rect 488816 6326 488868 6332
rect 489184 6384 489236 6390
rect 489184 6326 489236 6332
rect 486424 5568 486476 5574
rect 486424 5510 486476 5516
rect 487620 5568 487672 5574
rect 487620 5510 487672 5516
rect 486344 3454 486464 3482
rect 486436 480 486464 3454
rect 487632 480 487660 5510
rect 488828 480 488856 6326
rect 489932 480 489960 39782
rect 493324 39772 493376 39778
rect 493324 39714 493376 39720
rect 492680 22772 492732 22778
rect 492680 22714 492732 22720
rect 492692 16574 492720 22714
rect 492692 16546 493088 16574
rect 491116 8084 491168 8090
rect 491116 8026 491168 8032
rect 491128 480 491156 8026
rect 492312 6452 492364 6458
rect 492312 6394 492364 6400
rect 492324 480 492352 6394
rect 493060 490 493088 16546
rect 493336 5574 493364 39714
rect 496820 39704 496872 39710
rect 496820 39646 496872 39652
rect 496832 16574 496860 39646
rect 503720 39636 503772 39642
rect 503720 39578 503772 39584
rect 500960 38344 501012 38350
rect 500960 38286 501012 38292
rect 499580 36916 499632 36922
rect 499580 36858 499632 36864
rect 499592 16574 499620 36858
rect 500972 16574 501000 38286
rect 496832 16546 497136 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 495900 6316 495952 6322
rect 495900 6258 495952 6264
rect 493324 5568 493376 5574
rect 493324 5510 493376 5516
rect 494704 5568 494756 5574
rect 494704 5510 494756 5516
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 5510
rect 495912 480 495940 6258
rect 497108 480 497136 16546
rect 498200 6384 498252 6390
rect 498200 6326 498252 6332
rect 498212 480 498240 6326
rect 499396 6248 499448 6254
rect 499396 6190 499448 6196
rect 499408 480 499436 6190
rect 500604 480 500632 16546
rect 501340 490 501368 16546
rect 502984 6180 503036 6186
rect 502984 6122 503036 6128
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 6122
rect 503732 490 503760 39578
rect 510620 39568 510672 39574
rect 510620 39510 510672 39516
rect 507860 38276 507912 38282
rect 507860 38218 507912 38224
rect 506480 36848 506532 36854
rect 506480 36790 506532 36796
rect 506492 16574 506520 36790
rect 507872 16574 507900 38218
rect 510632 16574 510660 39510
rect 512644 39500 512696 39506
rect 512644 39442 512696 39448
rect 506492 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 506480 8968 506532 8974
rect 506480 8910 506532 8916
rect 505376 6860 505428 6866
rect 505376 6802 505428 6808
rect 504008 598 504220 626
rect 504008 490 504036 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 6802
rect 506492 480 506520 8910
rect 507228 490 507256 16546
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 16546
rect 510068 8016 510120 8022
rect 510068 7958 510120 7964
rect 510080 480 510108 7958
rect 511276 480 511304 16546
rect 512656 5574 512684 39442
rect 522304 39432 522356 39438
rect 522304 39374 522356 39380
rect 520280 38208 520332 38214
rect 520280 38150 520332 38156
rect 514760 35216 514812 35222
rect 514760 35158 514812 35164
rect 512644 5568 512696 5574
rect 512644 5510 512696 5516
rect 513564 5568 513616 5574
rect 513564 5510 513616 5516
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 512472 480 512500 4218
rect 513576 480 513604 5510
rect 514772 480 514800 35158
rect 517152 7948 517204 7954
rect 517152 7890 517204 7896
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 515968 480 515996 4286
rect 517164 480 517192 7890
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 518348 2916 518400 2922
rect 518348 2858 518400 2864
rect 518360 480 518388 2858
rect 519556 480 519584 4354
rect 520292 490 520320 38150
rect 522316 4214 522344 39374
rect 574744 39364 574796 39370
rect 574744 39306 574796 39312
rect 538220 38140 538272 38146
rect 538220 38082 538272 38088
rect 538232 16574 538260 38082
rect 547880 38072 547932 38078
rect 547880 38014 547932 38020
rect 547892 16574 547920 38014
rect 551284 38004 551336 38010
rect 551284 37946 551336 37952
rect 538232 16546 538444 16574
rect 547892 16546 548656 16574
rect 527824 7880 527876 7886
rect 527824 7822 527876 7828
rect 523040 4548 523092 4554
rect 523040 4490 523092 4496
rect 522304 4208 522356 4214
rect 522304 4150 522356 4156
rect 521844 3052 521896 3058
rect 521844 2994 521896 3000
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 2994
rect 523052 480 523080 4490
rect 526628 4480 526680 4486
rect 526628 4422 526680 4428
rect 524236 4208 524288 4214
rect 524236 4150 524288 4156
rect 524248 480 524276 4150
rect 525432 2984 525484 2990
rect 525432 2926 525484 2932
rect 525444 480 525472 2926
rect 526640 480 526668 4422
rect 527836 480 527864 7822
rect 534908 7812 534960 7818
rect 534908 7754 534960 7760
rect 531320 7744 531372 7750
rect 531320 7686 531372 7692
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 529020 3188 529072 3194
rect 529020 3130 529072 3136
rect 529032 480 529060 3130
rect 530136 480 530164 4558
rect 531332 480 531360 7686
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 532516 3120 532568 3126
rect 532516 3062 532568 3068
rect 532528 480 532556 3062
rect 533724 480 533752 4626
rect 534920 480 534948 7754
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 536104 3256 536156 3262
rect 536104 3198 536156 3204
rect 536116 480 536144 3198
rect 537220 480 537248 4694
rect 538416 480 538444 16546
rect 541992 7676 542044 7682
rect 541992 7618 542044 7624
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 539600 3324 539652 3330
rect 539600 3266 539652 3272
rect 539612 480 539640 3266
rect 540808 480 540836 5442
rect 542004 480 542032 7618
rect 545488 7608 545540 7614
rect 545488 7550 545540 7556
rect 544384 5432 544436 5438
rect 544384 5374 544436 5380
rect 543188 3392 543240 3398
rect 543188 3334 543240 3340
rect 543200 480 543228 3334
rect 544396 480 544424 5374
rect 545500 480 545528 7550
rect 547880 5296 547932 5302
rect 547880 5238 547932 5244
rect 546684 4140 546736 4146
rect 546684 4082 546736 4088
rect 546696 480 546724 4082
rect 547892 480 547920 5238
rect 548628 490 548656 16546
rect 550272 4072 550324 4078
rect 550272 4014 550324 4020
rect 548904 598 549116 626
rect 548904 490 548932 598
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 462 548932 490
rect 549088 480 549116 598
rect 550284 480 550312 4014
rect 551296 3398 551324 37946
rect 560944 37936 560996 37942
rect 560944 37878 560996 37884
rect 556252 36780 556304 36786
rect 556252 36722 556304 36728
rect 556264 6914 556292 36722
rect 558184 36712 558236 36718
rect 558184 36654 558236 36660
rect 556172 6886 556292 6914
rect 551468 5364 551520 5370
rect 551468 5306 551520 5312
rect 551284 3392 551336 3398
rect 551284 3334 551336 3340
rect 551480 480 551508 5306
rect 554964 5160 555016 5166
rect 554964 5102 555016 5108
rect 553768 3936 553820 3942
rect 553768 3878 553820 3884
rect 552664 3392 552716 3398
rect 552664 3334 552716 3340
rect 552676 480 552704 3334
rect 553780 480 553808 3878
rect 554976 480 555004 5102
rect 556172 480 556200 6886
rect 557356 4004 557408 4010
rect 557356 3946 557408 3952
rect 557368 480 557396 3946
rect 558196 3398 558224 36654
rect 558552 5228 558604 5234
rect 558552 5170 558604 5176
rect 558184 3392 558236 3398
rect 558184 3334 558236 3340
rect 558564 480 558592 5170
rect 560852 3868 560904 3874
rect 560852 3810 560904 3816
rect 559748 3392 559800 3398
rect 559748 3334 559800 3340
rect 559760 480 559788 3334
rect 560864 480 560892 3810
rect 560956 3058 560984 37878
rect 565820 36644 565872 36650
rect 565820 36586 565872 36592
rect 565832 16574 565860 36586
rect 572720 36576 572772 36582
rect 572720 36518 572772 36524
rect 572732 16574 572760 36518
rect 565832 16546 566872 16574
rect 572732 16546 573496 16574
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 560944 3052 560996 3058
rect 560944 2994 560996 3000
rect 562060 480 562088 5034
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 564440 3800 564492 3806
rect 564440 3742 564492 3748
rect 563244 3052 563296 3058
rect 563244 2994 563296 3000
rect 563256 480 563284 2994
rect 564452 480 564480 3742
rect 565648 480 565676 4966
rect 566844 480 566872 16546
rect 569224 10328 569276 10334
rect 569224 10270 569276 10276
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 3732 568080 3738
rect 568028 3674 568080 3680
rect 568040 480 568068 3674
rect 569144 480 569172 4898
rect 569236 3262 569264 10270
rect 572720 4820 572772 4826
rect 572720 4762 572772 4768
rect 571524 3664 571576 3670
rect 571524 3606 571576 3612
rect 569224 3256 569276 3262
rect 569224 3198 569276 3204
rect 570328 3256 570380 3262
rect 570328 3198 570380 3204
rect 570340 480 570368 3198
rect 571536 480 571564 3606
rect 572732 480 572760 4762
rect 573468 490 573496 16546
rect 574756 4146 574784 39306
rect 576308 4888 576360 4894
rect 576308 4830 576360 4836
rect 574744 4140 574796 4146
rect 574744 4082 574796 4088
rect 575112 3528 575164 3534
rect 575112 3470 575164 3476
rect 573744 598 573956 626
rect 573744 490 573772 598
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 462 573772 490
rect 573928 480 573956 598
rect 575124 480 575152 3470
rect 576320 480 576348 4830
rect 577412 4140 577464 4146
rect 577412 4082 577464 4088
rect 577424 480 577452 4082
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 580998 3496 581054 3505
rect 578608 3460 578660 3466
rect 580998 3431 581054 3440
rect 578608 3402 578660 3408
rect 578620 480 578648 3402
rect 581012 480 581040 3431
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3422 462576 3478 462632
rect 3330 449520 3386 449576
rect 2962 410488 3018 410544
rect 3238 397432 3294 397488
rect 2778 371356 2780 371376
rect 2780 371356 2832 371376
rect 2832 371356 2834 371376
rect 2778 371320 2834 371356
rect 3330 358400 3386 358456
rect 3146 345344 3202 345400
rect 3054 293120 3110 293176
rect 3146 254088 3202 254144
rect 3514 423544 3570 423600
rect 3514 319232 3570 319288
rect 3514 306176 3570 306232
rect 3514 267144 3570 267200
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 2778 136720 2834 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 2870 32408 2926 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 13818 467744 13874 467800
rect 35254 467608 35310 467664
rect 43994 468016 44050 468072
rect 47858 468016 47914 468072
rect 51538 468016 51594 468072
rect 62762 468016 62818 468072
rect 73802 468016 73858 468072
rect 126058 468016 126114 468072
rect 137282 468016 137338 468072
rect 363878 468016 363934 468072
rect 374918 468016 374974 468072
rect 397458 468016 397514 468072
rect 40774 466928 40830 466984
rect 504362 467472 504418 467528
rect 502982 467336 503038 467392
rect 508502 467200 508558 467256
rect 507122 467064 507178 467120
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 579618 404912 579674 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 579618 298696 579674 298752
rect 579894 272176 579950 272232
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 579894 219000 579950 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 579986 179152 580042 179208
rect 580170 165824 580226 165880
rect 580446 431568 580502 431624
rect 580354 418240 580410 418296
rect 580262 152632 580318 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 365626 3440 365682 3496
rect 379426 3304 379482 3360
rect 386234 3712 386290 3768
rect 389086 3576 389142 3632
rect 443826 3440 443882 3496
rect 461582 3304 461638 3360
rect 464986 3440 465042 3496
rect 466366 3304 466422 3360
rect 472254 3712 472310 3768
rect 475750 3576 475806 3632
rect 580998 3440 581054 3496
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect 43989 468076 44055 468077
rect 43989 468072 44036 468076
rect 44100 468074 44106 468076
rect 47853 468074 47919 468077
rect 48078 468074 48084 468076
rect 43989 468016 43994 468072
rect 43989 468012 44036 468016
rect 44100 468014 44146 468074
rect 47853 468072 48084 468074
rect 47853 468016 47858 468072
rect 47914 468016 48084 468072
rect 47853 468014 48084 468016
rect 44100 468012 44106 468014
rect 43989 468011 44055 468012
rect 47853 468011 47919 468014
rect 48078 468012 48084 468014
rect 48148 468012 48154 468076
rect 51533 468074 51599 468077
rect 62757 468076 62823 468077
rect 73797 468076 73863 468077
rect 126053 468076 126119 468077
rect 137277 468076 137343 468077
rect 52310 468074 52316 468076
rect 51533 468072 52316 468074
rect 51533 468016 51538 468072
rect 51594 468016 52316 468072
rect 51533 468014 52316 468016
rect 51533 468011 51599 468014
rect 52310 468012 52316 468014
rect 52380 468012 52386 468076
rect 62757 468072 62804 468076
rect 62868 468074 62874 468076
rect 62757 468016 62762 468072
rect 62757 468012 62804 468016
rect 62868 468014 62914 468074
rect 73797 468072 73844 468076
rect 73908 468074 73914 468076
rect 73797 468016 73802 468072
rect 62868 468012 62874 468014
rect 73797 468012 73844 468016
rect 73908 468014 73954 468074
rect 126053 468072 126100 468076
rect 126164 468074 126170 468076
rect 126053 468016 126058 468072
rect 73908 468012 73914 468014
rect 126053 468012 126100 468016
rect 126164 468014 126210 468074
rect 137277 468072 137324 468076
rect 137388 468074 137394 468076
rect 363873 468074 363939 468077
rect 374913 468076 374979 468077
rect 374862 468074 374868 468076
rect 137277 468016 137282 468072
rect 126164 468012 126170 468014
rect 137277 468012 137324 468016
rect 137388 468014 137434 468074
rect 363830 468072 363939 468074
rect 363830 468016 363878 468072
rect 363934 468016 363939 468072
rect 137388 468012 137394 468014
rect 62757 468011 62823 468012
rect 73797 468011 73863 468012
rect 126053 468011 126119 468012
rect 137277 468011 137343 468012
rect 363830 468011 363939 468016
rect 374822 468014 374868 468074
rect 374932 468072 374979 468076
rect 397453 468074 397519 468077
rect 374974 468016 374979 468072
rect 374862 468012 374868 468014
rect 374932 468012 374979 468016
rect 374913 468011 374979 468012
rect 397318 468072 397519 468074
rect 397318 468016 397458 468072
rect 397514 468016 397519 468072
rect 397318 468014 397519 468016
rect 13813 467802 13879 467805
rect 363830 467802 363890 468011
rect 13813 467800 363890 467802
rect 13813 467744 13818 467800
rect 13874 467744 363890 467800
rect 13813 467742 363890 467744
rect 13813 467739 13879 467742
rect 35249 467666 35315 467669
rect 397318 467666 397378 468014
rect 397453 468011 397519 468014
rect 35249 467664 397378 467666
rect 35249 467608 35254 467664
rect 35310 467608 397378 467664
rect 35249 467606 397378 467608
rect 35249 467603 35315 467606
rect 137318 467468 137324 467532
rect 137388 467530 137394 467532
rect 504357 467530 504423 467533
rect 137388 467528 504423 467530
rect 137388 467472 504362 467528
rect 504418 467472 504423 467528
rect 137388 467470 504423 467472
rect 137388 467468 137394 467470
rect 504357 467467 504423 467470
rect 126094 467332 126100 467396
rect 126164 467394 126170 467396
rect 502977 467394 503043 467397
rect 126164 467392 503043 467394
rect 126164 467336 502982 467392
rect 503038 467336 503043 467392
rect 126164 467334 503043 467336
rect 126164 467332 126170 467334
rect 502977 467331 503043 467334
rect 73838 467196 73844 467260
rect 73908 467258 73914 467260
rect 508497 467258 508563 467261
rect 73908 467256 508563 467258
rect 73908 467200 508502 467256
rect 508558 467200 508563 467256
rect 73908 467198 508563 467200
rect 73908 467196 73914 467198
rect 508497 467195 508563 467198
rect 62798 467060 62804 467124
rect 62868 467122 62874 467124
rect 507117 467122 507183 467125
rect 62868 467120 507183 467122
rect 62868 467064 507122 467120
rect 507178 467064 507183 467120
rect 62868 467062 507183 467064
rect 62868 467060 62874 467062
rect 507117 467059 507183 467062
rect 40769 466986 40835 466989
rect 374862 466986 374868 466988
rect 40769 466984 374868 466986
rect 40769 466928 40774 466984
rect 40830 466928 374868 466984
rect 40769 466926 374868 466928
rect 40769 466923 40835 466926
rect 374862 466924 374868 466926
rect 374932 466924 374938 466988
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580441 431626 580507 431629
rect 583520 431626 584960 431716
rect 580441 431624 584960 431626
rect 580441 431568 580446 431624
rect 580502 431568 584960 431624
rect 580441 431566 584960 431568
rect 580441 431563 580507 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580349 418298 580415 418301
rect 583520 418298 584960 418388
rect 580349 418296 584960 418298
rect 580349 418240 580354 418296
rect 580410 418240 584960 418296
rect 580349 418238 584960 418240
rect 580349 418235 580415 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 579613 404970 579679 404973
rect 583520 404970 584960 405060
rect 579613 404968 584960 404970
rect 579613 404912 579618 404968
rect 579674 404912 584960 404968
rect 579613 404910 584960 404912
rect 579613 404907 579679 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3233 397490 3299 397493
rect -960 397488 3299 397490
rect -960 397432 3238 397488
rect 3294 397432 3299 397488
rect -960 397430 3299 397432
rect -960 397340 480 397430
rect 3233 397427 3299 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2773 371378 2839 371381
rect -960 371376 2839 371378
rect -960 371320 2778 371376
rect 2834 371320 2839 371376
rect -960 371318 2839 371320
rect -960 371228 480 371318
rect 2773 371315 2839 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579889 219058 579955 219061
rect 583520 219058 584960 219148
rect 579889 219056 584960 219058
rect 579889 219000 579894 219056
rect 579950 219000 584960 219056
rect 579889 218998 584960 219000
rect 579889 218995 579955 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 2773 136778 2839 136781
rect -960 136776 2839 136778
rect -960 136720 2778 136776
rect 2834 136720 2839 136776
rect -960 136718 2839 136720
rect -960 136628 480 136718
rect 2773 136715 2839 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 48078 31724 48084 31788
rect 48148 31786 48154 31788
rect 583526 31786 583586 32950
rect 48148 31726 583586 31786
rect 48148 31724 48154 31726
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 52310 19348 52316 19412
rect 52380 19410 52386 19412
rect 583526 19410 583586 19622
rect 52380 19350 583586 19410
rect 52380 19348 52386 19350
rect 583520 6626 584960 6716
rect -960 6490 480 6580
rect 583342 6566 584960 6626
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect 583342 6490 583402 6566
rect 583520 6490 584960 6566
rect 583342 6476 584960 6490
rect 583342 6430 583586 6476
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 44030 5612 44036 5676
rect 44100 5674 44106 5676
rect 583526 5674 583586 6430
rect 44100 5614 583586 5674
rect 44100 5612 44106 5614
rect 386229 3770 386295 3773
rect 472249 3770 472315 3773
rect 386229 3768 472315 3770
rect 386229 3712 386234 3768
rect 386290 3712 472254 3768
rect 472310 3712 472315 3768
rect 386229 3710 472315 3712
rect 386229 3707 386295 3710
rect 472249 3707 472315 3710
rect 389081 3634 389147 3637
rect 475745 3634 475811 3637
rect 389081 3632 475811 3634
rect 389081 3576 389086 3632
rect 389142 3576 475750 3632
rect 475806 3576 475811 3632
rect 389081 3574 475811 3576
rect 389081 3571 389147 3574
rect 475745 3571 475811 3574
rect 365621 3498 365687 3501
rect 443821 3498 443887 3501
rect 365621 3496 443887 3498
rect 365621 3440 365626 3496
rect 365682 3440 443826 3496
rect 443882 3440 443887 3496
rect 365621 3438 443887 3440
rect 365621 3435 365687 3438
rect 443821 3435 443887 3438
rect 464981 3498 465047 3501
rect 580993 3498 581059 3501
rect 464981 3496 581059 3498
rect 464981 3440 464986 3496
rect 465042 3440 580998 3496
rect 581054 3440 581059 3496
rect 464981 3438 581059 3440
rect 464981 3435 465047 3438
rect 580993 3435 581059 3438
rect 379421 3362 379487 3365
rect 461577 3362 461643 3365
rect 379421 3360 461643 3362
rect 379421 3304 379426 3360
rect 379482 3304 461582 3360
rect 461638 3304 461643 3360
rect 379421 3302 461643 3304
rect 379421 3299 379487 3302
rect 461577 3299 461643 3302
rect 466361 3362 466427 3365
rect 583385 3362 583451 3365
rect 466361 3360 583451 3362
rect 466361 3304 466366 3360
rect 466422 3304 583390 3360
rect 583446 3304 583451 3360
rect 466361 3302 583451 3304
rect 466361 3299 466427 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 44036 468072 44100 468076
rect 44036 468016 44050 468072
rect 44050 468016 44100 468072
rect 44036 468012 44100 468016
rect 48084 468012 48148 468076
rect 52316 468012 52380 468076
rect 62804 468072 62868 468076
rect 62804 468016 62818 468072
rect 62818 468016 62868 468072
rect 62804 468012 62868 468016
rect 73844 468072 73908 468076
rect 73844 468016 73858 468072
rect 73858 468016 73908 468072
rect 73844 468012 73908 468016
rect 126100 468072 126164 468076
rect 126100 468016 126114 468072
rect 126114 468016 126164 468072
rect 126100 468012 126164 468016
rect 137324 468072 137388 468076
rect 137324 468016 137338 468072
rect 137338 468016 137388 468072
rect 137324 468012 137388 468016
rect 374868 468072 374932 468076
rect 374868 468016 374918 468072
rect 374918 468016 374932 468072
rect 374868 468012 374932 468016
rect 137324 467468 137388 467532
rect 126100 467332 126164 467396
rect 73844 467196 73908 467260
rect 62804 467060 62868 467124
rect 374868 466924 374932 466988
rect 48084 31724 48148 31788
rect 52316 19348 52380 19412
rect 44036 5612 44100 5676
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 470704 42134 474618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 470704 45854 478338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 470704 49574 482058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 470704 56414 488898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 470704 60134 492618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 470704 63854 496338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 470704 67574 500058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 470704 74414 470898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 470704 78134 474618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 470704 81854 478338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 470704 85574 482058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 470704 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 470704 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 470704 99854 496338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 470704 103574 500058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 470704 110414 470898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 470704 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 470704 117854 478338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 470704 121574 482058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 470704 128414 488898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 470704 132134 492618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 470704 135854 496338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 470704 139574 500058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 470704 146414 470898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 470704 150134 474618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 470704 153854 478338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 470704 157574 482058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 470704 164414 488898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 470704 168134 492618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 470704 171854 496338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 470704 175574 500058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 470704 182414 470898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 470704 186134 474618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 470704 189854 478338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 470704 193574 482058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 470704 200414 488898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 470704 204134 492618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 470704 207854 496338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 470704 211574 500058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 470704 218414 470898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 470704 222134 474618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 470704 225854 478338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 470704 229574 482058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 470704 236414 488898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 470704 240134 492618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 470704 243854 496338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 470704 247574 500058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 470704 254414 470898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 470704 258134 474618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 470704 261854 478338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 470704 265574 482058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 470704 272414 488898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 470704 276134 492618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 470704 279854 496338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 470704 283574 500058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 470704 290414 470898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 470704 294134 474618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 470704 297854 478338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 470704 301574 482058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 470704 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 470704 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 470704 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 470704 319574 500058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 470704 326414 470898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 470704 330134 474618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 470704 333854 478338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 470704 337574 482058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 470704 344414 488898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 470704 348134 492618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 470704 351854 496338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 470704 355574 500058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 470704 362414 470898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 470704 366134 474618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 470704 369854 478338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 470704 373574 482058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 470704 380414 488898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 470704 384134 492618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 470704 387854 496338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 470704 391574 500058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 470704 398414 470898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 470704 402134 474618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 470704 405854 478338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 470704 409574 482058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 470704 416414 488898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 470704 420134 492618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 470704 423854 496338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 470704 427574 500058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 470704 434414 470898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 470704 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 470704 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 470704 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 470704 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 470704 456134 492618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 470704 459854 496338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 470704 463574 500058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 44035 468076 44101 468077
rect 44035 468012 44036 468076
rect 44100 468012 44101 468076
rect 44035 468011 44101 468012
rect 48083 468076 48149 468077
rect 48083 468012 48084 468076
rect 48148 468012 48149 468076
rect 48083 468011 48149 468012
rect 52315 468076 52381 468077
rect 52315 468012 52316 468076
rect 52380 468012 52381 468076
rect 52315 468011 52381 468012
rect 62803 468076 62869 468077
rect 62803 468012 62804 468076
rect 62868 468012 62869 468076
rect 62803 468011 62869 468012
rect 73843 468076 73909 468077
rect 73843 468012 73844 468076
rect 73908 468012 73909 468076
rect 73843 468011 73909 468012
rect 126099 468076 126165 468077
rect 126099 468012 126100 468076
rect 126164 468012 126165 468076
rect 126099 468011 126165 468012
rect 137323 468076 137389 468077
rect 137323 468012 137324 468076
rect 137388 468012 137389 468076
rect 137323 468011 137389 468012
rect 374867 468076 374933 468077
rect 374867 468012 374868 468076
rect 374932 468012 374933 468076
rect 374867 468011 374933 468012
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 7174 42134 40000
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 44038 5677 44098 468011
rect 46208 435454 46528 435486
rect 46208 435218 46250 435454
rect 46486 435218 46528 435454
rect 46208 435134 46528 435218
rect 46208 434898 46250 435134
rect 46486 434898 46528 435134
rect 46208 434866 46528 434898
rect 46208 399454 46528 399486
rect 46208 399218 46250 399454
rect 46486 399218 46528 399454
rect 46208 399134 46528 399218
rect 46208 398898 46250 399134
rect 46486 398898 46528 399134
rect 46208 398866 46528 398898
rect 46208 363454 46528 363486
rect 46208 363218 46250 363454
rect 46486 363218 46528 363454
rect 46208 363134 46528 363218
rect 46208 362898 46250 363134
rect 46486 362898 46528 363134
rect 46208 362866 46528 362898
rect 46208 327454 46528 327486
rect 46208 327218 46250 327454
rect 46486 327218 46528 327454
rect 46208 327134 46528 327218
rect 46208 326898 46250 327134
rect 46486 326898 46528 327134
rect 46208 326866 46528 326898
rect 46208 291454 46528 291486
rect 46208 291218 46250 291454
rect 46486 291218 46528 291454
rect 46208 291134 46528 291218
rect 46208 290898 46250 291134
rect 46486 290898 46528 291134
rect 46208 290866 46528 290898
rect 46208 255454 46528 255486
rect 46208 255218 46250 255454
rect 46486 255218 46528 255454
rect 46208 255134 46528 255218
rect 46208 254898 46250 255134
rect 46486 254898 46528 255134
rect 46208 254866 46528 254898
rect 46208 219454 46528 219486
rect 46208 219218 46250 219454
rect 46486 219218 46528 219454
rect 46208 219134 46528 219218
rect 46208 218898 46250 219134
rect 46486 218898 46528 219134
rect 46208 218866 46528 218898
rect 46208 183454 46528 183486
rect 46208 183218 46250 183454
rect 46486 183218 46528 183454
rect 46208 183134 46528 183218
rect 46208 182898 46250 183134
rect 46486 182898 46528 183134
rect 46208 182866 46528 182898
rect 46208 147454 46528 147486
rect 46208 147218 46250 147454
rect 46486 147218 46528 147454
rect 46208 147134 46528 147218
rect 46208 146898 46250 147134
rect 46486 146898 46528 147134
rect 46208 146866 46528 146898
rect 46208 111454 46528 111486
rect 46208 111218 46250 111454
rect 46486 111218 46528 111454
rect 46208 111134 46528 111218
rect 46208 110898 46250 111134
rect 46486 110898 46528 111134
rect 46208 110866 46528 110898
rect 46208 75454 46528 75486
rect 46208 75218 46250 75454
rect 46486 75218 46528 75454
rect 46208 75134 46528 75218
rect 46208 74898 46250 75134
rect 46486 74898 46528 75134
rect 46208 74866 46528 74898
rect 45234 10894 45854 40000
rect 48086 31789 48146 468011
rect 48083 31788 48149 31789
rect 48083 31724 48084 31788
rect 48148 31724 48149 31788
rect 48083 31723 48149 31724
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 44035 5676 44101 5677
rect 44035 5612 44036 5676
rect 44100 5612 44101 5676
rect 44035 5611 44101 5612
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 40000
rect 52318 19413 52378 468011
rect 62806 467125 62866 468011
rect 73846 467261 73906 468011
rect 126102 467397 126162 468011
rect 137326 467533 137386 468011
rect 137323 467532 137389 467533
rect 137323 467468 137324 467532
rect 137388 467468 137389 467532
rect 137323 467467 137389 467468
rect 126099 467396 126165 467397
rect 126099 467332 126100 467396
rect 126164 467332 126165 467396
rect 126099 467331 126165 467332
rect 73843 467260 73909 467261
rect 73843 467196 73844 467260
rect 73908 467196 73909 467260
rect 73843 467195 73909 467196
rect 62803 467124 62869 467125
rect 62803 467060 62804 467124
rect 62868 467060 62869 467124
rect 62803 467059 62869 467060
rect 374870 466989 374930 468011
rect 374867 466988 374933 466989
rect 374867 466924 374868 466988
rect 374932 466924 374933 466988
rect 374867 466923 374933 466924
rect 61568 453454 61888 453486
rect 61568 453218 61610 453454
rect 61846 453218 61888 453454
rect 61568 453134 61888 453218
rect 61568 452898 61610 453134
rect 61846 452898 61888 453134
rect 61568 452866 61888 452898
rect 92288 453454 92608 453486
rect 92288 453218 92330 453454
rect 92566 453218 92608 453454
rect 92288 453134 92608 453218
rect 92288 452898 92330 453134
rect 92566 452898 92608 453134
rect 92288 452866 92608 452898
rect 123008 453454 123328 453486
rect 123008 453218 123050 453454
rect 123286 453218 123328 453454
rect 123008 453134 123328 453218
rect 123008 452898 123050 453134
rect 123286 452898 123328 453134
rect 123008 452866 123328 452898
rect 153728 453454 154048 453486
rect 153728 453218 153770 453454
rect 154006 453218 154048 453454
rect 153728 453134 154048 453218
rect 153728 452898 153770 453134
rect 154006 452898 154048 453134
rect 153728 452866 154048 452898
rect 184448 453454 184768 453486
rect 184448 453218 184490 453454
rect 184726 453218 184768 453454
rect 184448 453134 184768 453218
rect 184448 452898 184490 453134
rect 184726 452898 184768 453134
rect 184448 452866 184768 452898
rect 215168 453454 215488 453486
rect 215168 453218 215210 453454
rect 215446 453218 215488 453454
rect 215168 453134 215488 453218
rect 215168 452898 215210 453134
rect 215446 452898 215488 453134
rect 215168 452866 215488 452898
rect 245888 453454 246208 453486
rect 245888 453218 245930 453454
rect 246166 453218 246208 453454
rect 245888 453134 246208 453218
rect 245888 452898 245930 453134
rect 246166 452898 246208 453134
rect 245888 452866 246208 452898
rect 276608 453454 276928 453486
rect 276608 453218 276650 453454
rect 276886 453218 276928 453454
rect 276608 453134 276928 453218
rect 276608 452898 276650 453134
rect 276886 452898 276928 453134
rect 276608 452866 276928 452898
rect 307328 453454 307648 453486
rect 307328 453218 307370 453454
rect 307606 453218 307648 453454
rect 307328 453134 307648 453218
rect 307328 452898 307370 453134
rect 307606 452898 307648 453134
rect 307328 452866 307648 452898
rect 338048 453454 338368 453486
rect 338048 453218 338090 453454
rect 338326 453218 338368 453454
rect 338048 453134 338368 453218
rect 338048 452898 338090 453134
rect 338326 452898 338368 453134
rect 338048 452866 338368 452898
rect 368768 453454 369088 453486
rect 368768 453218 368810 453454
rect 369046 453218 369088 453454
rect 368768 453134 369088 453218
rect 368768 452898 368810 453134
rect 369046 452898 369088 453134
rect 368768 452866 369088 452898
rect 399488 453454 399808 453486
rect 399488 453218 399530 453454
rect 399766 453218 399808 453454
rect 399488 453134 399808 453218
rect 399488 452898 399530 453134
rect 399766 452898 399808 453134
rect 399488 452866 399808 452898
rect 430208 453454 430528 453486
rect 430208 453218 430250 453454
rect 430486 453218 430528 453454
rect 430208 453134 430528 453218
rect 430208 452898 430250 453134
rect 430486 452898 430528 453134
rect 430208 452866 430528 452898
rect 460928 453454 461248 453486
rect 460928 453218 460970 453454
rect 461206 453218 461248 453454
rect 460928 453134 461248 453218
rect 460928 452898 460970 453134
rect 461206 452898 461248 453134
rect 460928 452866 461248 452898
rect 76928 435454 77248 435486
rect 76928 435218 76970 435454
rect 77206 435218 77248 435454
rect 76928 435134 77248 435218
rect 76928 434898 76970 435134
rect 77206 434898 77248 435134
rect 76928 434866 77248 434898
rect 107648 435454 107968 435486
rect 107648 435218 107690 435454
rect 107926 435218 107968 435454
rect 107648 435134 107968 435218
rect 107648 434898 107690 435134
rect 107926 434898 107968 435134
rect 107648 434866 107968 434898
rect 138368 435454 138688 435486
rect 138368 435218 138410 435454
rect 138646 435218 138688 435454
rect 138368 435134 138688 435218
rect 138368 434898 138410 435134
rect 138646 434898 138688 435134
rect 138368 434866 138688 434898
rect 169088 435454 169408 435486
rect 169088 435218 169130 435454
rect 169366 435218 169408 435454
rect 169088 435134 169408 435218
rect 169088 434898 169130 435134
rect 169366 434898 169408 435134
rect 169088 434866 169408 434898
rect 199808 435454 200128 435486
rect 199808 435218 199850 435454
rect 200086 435218 200128 435454
rect 199808 435134 200128 435218
rect 199808 434898 199850 435134
rect 200086 434898 200128 435134
rect 199808 434866 200128 434898
rect 230528 435454 230848 435486
rect 230528 435218 230570 435454
rect 230806 435218 230848 435454
rect 230528 435134 230848 435218
rect 230528 434898 230570 435134
rect 230806 434898 230848 435134
rect 230528 434866 230848 434898
rect 261248 435454 261568 435486
rect 261248 435218 261290 435454
rect 261526 435218 261568 435454
rect 261248 435134 261568 435218
rect 261248 434898 261290 435134
rect 261526 434898 261568 435134
rect 261248 434866 261568 434898
rect 291968 435454 292288 435486
rect 291968 435218 292010 435454
rect 292246 435218 292288 435454
rect 291968 435134 292288 435218
rect 291968 434898 292010 435134
rect 292246 434898 292288 435134
rect 291968 434866 292288 434898
rect 322688 435454 323008 435486
rect 322688 435218 322730 435454
rect 322966 435218 323008 435454
rect 322688 435134 323008 435218
rect 322688 434898 322730 435134
rect 322966 434898 323008 435134
rect 322688 434866 323008 434898
rect 353408 435454 353728 435486
rect 353408 435218 353450 435454
rect 353686 435218 353728 435454
rect 353408 435134 353728 435218
rect 353408 434898 353450 435134
rect 353686 434898 353728 435134
rect 353408 434866 353728 434898
rect 384128 435454 384448 435486
rect 384128 435218 384170 435454
rect 384406 435218 384448 435454
rect 384128 435134 384448 435218
rect 384128 434898 384170 435134
rect 384406 434898 384448 435134
rect 384128 434866 384448 434898
rect 414848 435454 415168 435486
rect 414848 435218 414890 435454
rect 415126 435218 415168 435454
rect 414848 435134 415168 435218
rect 414848 434898 414890 435134
rect 415126 434898 415168 435134
rect 414848 434866 415168 434898
rect 445568 435454 445888 435486
rect 445568 435218 445610 435454
rect 445846 435218 445888 435454
rect 445568 435134 445888 435218
rect 445568 434898 445610 435134
rect 445846 434898 445888 435134
rect 445568 434866 445888 434898
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 61568 417454 61888 417486
rect 61568 417218 61610 417454
rect 61846 417218 61888 417454
rect 61568 417134 61888 417218
rect 61568 416898 61610 417134
rect 61846 416898 61888 417134
rect 61568 416866 61888 416898
rect 92288 417454 92608 417486
rect 92288 417218 92330 417454
rect 92566 417218 92608 417454
rect 92288 417134 92608 417218
rect 92288 416898 92330 417134
rect 92566 416898 92608 417134
rect 92288 416866 92608 416898
rect 123008 417454 123328 417486
rect 123008 417218 123050 417454
rect 123286 417218 123328 417454
rect 123008 417134 123328 417218
rect 123008 416898 123050 417134
rect 123286 416898 123328 417134
rect 123008 416866 123328 416898
rect 153728 417454 154048 417486
rect 153728 417218 153770 417454
rect 154006 417218 154048 417454
rect 153728 417134 154048 417218
rect 153728 416898 153770 417134
rect 154006 416898 154048 417134
rect 153728 416866 154048 416898
rect 184448 417454 184768 417486
rect 184448 417218 184490 417454
rect 184726 417218 184768 417454
rect 184448 417134 184768 417218
rect 184448 416898 184490 417134
rect 184726 416898 184768 417134
rect 184448 416866 184768 416898
rect 215168 417454 215488 417486
rect 215168 417218 215210 417454
rect 215446 417218 215488 417454
rect 215168 417134 215488 417218
rect 215168 416898 215210 417134
rect 215446 416898 215488 417134
rect 215168 416866 215488 416898
rect 245888 417454 246208 417486
rect 245888 417218 245930 417454
rect 246166 417218 246208 417454
rect 245888 417134 246208 417218
rect 245888 416898 245930 417134
rect 246166 416898 246208 417134
rect 245888 416866 246208 416898
rect 276608 417454 276928 417486
rect 276608 417218 276650 417454
rect 276886 417218 276928 417454
rect 276608 417134 276928 417218
rect 276608 416898 276650 417134
rect 276886 416898 276928 417134
rect 276608 416866 276928 416898
rect 307328 417454 307648 417486
rect 307328 417218 307370 417454
rect 307606 417218 307648 417454
rect 307328 417134 307648 417218
rect 307328 416898 307370 417134
rect 307606 416898 307648 417134
rect 307328 416866 307648 416898
rect 338048 417454 338368 417486
rect 338048 417218 338090 417454
rect 338326 417218 338368 417454
rect 338048 417134 338368 417218
rect 338048 416898 338090 417134
rect 338326 416898 338368 417134
rect 338048 416866 338368 416898
rect 368768 417454 369088 417486
rect 368768 417218 368810 417454
rect 369046 417218 369088 417454
rect 368768 417134 369088 417218
rect 368768 416898 368810 417134
rect 369046 416898 369088 417134
rect 368768 416866 369088 416898
rect 399488 417454 399808 417486
rect 399488 417218 399530 417454
rect 399766 417218 399808 417454
rect 399488 417134 399808 417218
rect 399488 416898 399530 417134
rect 399766 416898 399808 417134
rect 399488 416866 399808 416898
rect 430208 417454 430528 417486
rect 430208 417218 430250 417454
rect 430486 417218 430528 417454
rect 430208 417134 430528 417218
rect 430208 416898 430250 417134
rect 430486 416898 430528 417134
rect 430208 416866 430528 416898
rect 460928 417454 461248 417486
rect 460928 417218 460970 417454
rect 461206 417218 461248 417454
rect 460928 417134 461248 417218
rect 460928 416898 460970 417134
rect 461206 416898 461248 417134
rect 460928 416866 461248 416898
rect 76928 399454 77248 399486
rect 76928 399218 76970 399454
rect 77206 399218 77248 399454
rect 76928 399134 77248 399218
rect 76928 398898 76970 399134
rect 77206 398898 77248 399134
rect 76928 398866 77248 398898
rect 107648 399454 107968 399486
rect 107648 399218 107690 399454
rect 107926 399218 107968 399454
rect 107648 399134 107968 399218
rect 107648 398898 107690 399134
rect 107926 398898 107968 399134
rect 107648 398866 107968 398898
rect 138368 399454 138688 399486
rect 138368 399218 138410 399454
rect 138646 399218 138688 399454
rect 138368 399134 138688 399218
rect 138368 398898 138410 399134
rect 138646 398898 138688 399134
rect 138368 398866 138688 398898
rect 169088 399454 169408 399486
rect 169088 399218 169130 399454
rect 169366 399218 169408 399454
rect 169088 399134 169408 399218
rect 169088 398898 169130 399134
rect 169366 398898 169408 399134
rect 169088 398866 169408 398898
rect 199808 399454 200128 399486
rect 199808 399218 199850 399454
rect 200086 399218 200128 399454
rect 199808 399134 200128 399218
rect 199808 398898 199850 399134
rect 200086 398898 200128 399134
rect 199808 398866 200128 398898
rect 230528 399454 230848 399486
rect 230528 399218 230570 399454
rect 230806 399218 230848 399454
rect 230528 399134 230848 399218
rect 230528 398898 230570 399134
rect 230806 398898 230848 399134
rect 230528 398866 230848 398898
rect 261248 399454 261568 399486
rect 261248 399218 261290 399454
rect 261526 399218 261568 399454
rect 261248 399134 261568 399218
rect 261248 398898 261290 399134
rect 261526 398898 261568 399134
rect 261248 398866 261568 398898
rect 291968 399454 292288 399486
rect 291968 399218 292010 399454
rect 292246 399218 292288 399454
rect 291968 399134 292288 399218
rect 291968 398898 292010 399134
rect 292246 398898 292288 399134
rect 291968 398866 292288 398898
rect 322688 399454 323008 399486
rect 322688 399218 322730 399454
rect 322966 399218 323008 399454
rect 322688 399134 323008 399218
rect 322688 398898 322730 399134
rect 322966 398898 323008 399134
rect 322688 398866 323008 398898
rect 353408 399454 353728 399486
rect 353408 399218 353450 399454
rect 353686 399218 353728 399454
rect 353408 399134 353728 399218
rect 353408 398898 353450 399134
rect 353686 398898 353728 399134
rect 353408 398866 353728 398898
rect 384128 399454 384448 399486
rect 384128 399218 384170 399454
rect 384406 399218 384448 399454
rect 384128 399134 384448 399218
rect 384128 398898 384170 399134
rect 384406 398898 384448 399134
rect 384128 398866 384448 398898
rect 414848 399454 415168 399486
rect 414848 399218 414890 399454
rect 415126 399218 415168 399454
rect 414848 399134 415168 399218
rect 414848 398898 414890 399134
rect 415126 398898 415168 399134
rect 414848 398866 415168 398898
rect 445568 399454 445888 399486
rect 445568 399218 445610 399454
rect 445846 399218 445888 399454
rect 445568 399134 445888 399218
rect 445568 398898 445610 399134
rect 445846 398898 445888 399134
rect 445568 398866 445888 398898
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 61568 381454 61888 381486
rect 61568 381218 61610 381454
rect 61846 381218 61888 381454
rect 61568 381134 61888 381218
rect 61568 380898 61610 381134
rect 61846 380898 61888 381134
rect 61568 380866 61888 380898
rect 92288 381454 92608 381486
rect 92288 381218 92330 381454
rect 92566 381218 92608 381454
rect 92288 381134 92608 381218
rect 92288 380898 92330 381134
rect 92566 380898 92608 381134
rect 92288 380866 92608 380898
rect 123008 381454 123328 381486
rect 123008 381218 123050 381454
rect 123286 381218 123328 381454
rect 123008 381134 123328 381218
rect 123008 380898 123050 381134
rect 123286 380898 123328 381134
rect 123008 380866 123328 380898
rect 153728 381454 154048 381486
rect 153728 381218 153770 381454
rect 154006 381218 154048 381454
rect 153728 381134 154048 381218
rect 153728 380898 153770 381134
rect 154006 380898 154048 381134
rect 153728 380866 154048 380898
rect 184448 381454 184768 381486
rect 184448 381218 184490 381454
rect 184726 381218 184768 381454
rect 184448 381134 184768 381218
rect 184448 380898 184490 381134
rect 184726 380898 184768 381134
rect 184448 380866 184768 380898
rect 215168 381454 215488 381486
rect 215168 381218 215210 381454
rect 215446 381218 215488 381454
rect 215168 381134 215488 381218
rect 215168 380898 215210 381134
rect 215446 380898 215488 381134
rect 215168 380866 215488 380898
rect 245888 381454 246208 381486
rect 245888 381218 245930 381454
rect 246166 381218 246208 381454
rect 245888 381134 246208 381218
rect 245888 380898 245930 381134
rect 246166 380898 246208 381134
rect 245888 380866 246208 380898
rect 276608 381454 276928 381486
rect 276608 381218 276650 381454
rect 276886 381218 276928 381454
rect 276608 381134 276928 381218
rect 276608 380898 276650 381134
rect 276886 380898 276928 381134
rect 276608 380866 276928 380898
rect 307328 381454 307648 381486
rect 307328 381218 307370 381454
rect 307606 381218 307648 381454
rect 307328 381134 307648 381218
rect 307328 380898 307370 381134
rect 307606 380898 307648 381134
rect 307328 380866 307648 380898
rect 338048 381454 338368 381486
rect 338048 381218 338090 381454
rect 338326 381218 338368 381454
rect 338048 381134 338368 381218
rect 338048 380898 338090 381134
rect 338326 380898 338368 381134
rect 338048 380866 338368 380898
rect 368768 381454 369088 381486
rect 368768 381218 368810 381454
rect 369046 381218 369088 381454
rect 368768 381134 369088 381218
rect 368768 380898 368810 381134
rect 369046 380898 369088 381134
rect 368768 380866 369088 380898
rect 399488 381454 399808 381486
rect 399488 381218 399530 381454
rect 399766 381218 399808 381454
rect 399488 381134 399808 381218
rect 399488 380898 399530 381134
rect 399766 380898 399808 381134
rect 399488 380866 399808 380898
rect 430208 381454 430528 381486
rect 430208 381218 430250 381454
rect 430486 381218 430528 381454
rect 430208 381134 430528 381218
rect 430208 380898 430250 381134
rect 430486 380898 430528 381134
rect 430208 380866 430528 380898
rect 460928 381454 461248 381486
rect 460928 381218 460970 381454
rect 461206 381218 461248 381454
rect 460928 381134 461248 381218
rect 460928 380898 460970 381134
rect 461206 380898 461248 381134
rect 460928 380866 461248 380898
rect 76928 363454 77248 363486
rect 76928 363218 76970 363454
rect 77206 363218 77248 363454
rect 76928 363134 77248 363218
rect 76928 362898 76970 363134
rect 77206 362898 77248 363134
rect 76928 362866 77248 362898
rect 107648 363454 107968 363486
rect 107648 363218 107690 363454
rect 107926 363218 107968 363454
rect 107648 363134 107968 363218
rect 107648 362898 107690 363134
rect 107926 362898 107968 363134
rect 107648 362866 107968 362898
rect 138368 363454 138688 363486
rect 138368 363218 138410 363454
rect 138646 363218 138688 363454
rect 138368 363134 138688 363218
rect 138368 362898 138410 363134
rect 138646 362898 138688 363134
rect 138368 362866 138688 362898
rect 169088 363454 169408 363486
rect 169088 363218 169130 363454
rect 169366 363218 169408 363454
rect 169088 363134 169408 363218
rect 169088 362898 169130 363134
rect 169366 362898 169408 363134
rect 169088 362866 169408 362898
rect 199808 363454 200128 363486
rect 199808 363218 199850 363454
rect 200086 363218 200128 363454
rect 199808 363134 200128 363218
rect 199808 362898 199850 363134
rect 200086 362898 200128 363134
rect 199808 362866 200128 362898
rect 230528 363454 230848 363486
rect 230528 363218 230570 363454
rect 230806 363218 230848 363454
rect 230528 363134 230848 363218
rect 230528 362898 230570 363134
rect 230806 362898 230848 363134
rect 230528 362866 230848 362898
rect 261248 363454 261568 363486
rect 261248 363218 261290 363454
rect 261526 363218 261568 363454
rect 261248 363134 261568 363218
rect 261248 362898 261290 363134
rect 261526 362898 261568 363134
rect 261248 362866 261568 362898
rect 291968 363454 292288 363486
rect 291968 363218 292010 363454
rect 292246 363218 292288 363454
rect 291968 363134 292288 363218
rect 291968 362898 292010 363134
rect 292246 362898 292288 363134
rect 291968 362866 292288 362898
rect 322688 363454 323008 363486
rect 322688 363218 322730 363454
rect 322966 363218 323008 363454
rect 322688 363134 323008 363218
rect 322688 362898 322730 363134
rect 322966 362898 323008 363134
rect 322688 362866 323008 362898
rect 353408 363454 353728 363486
rect 353408 363218 353450 363454
rect 353686 363218 353728 363454
rect 353408 363134 353728 363218
rect 353408 362898 353450 363134
rect 353686 362898 353728 363134
rect 353408 362866 353728 362898
rect 384128 363454 384448 363486
rect 384128 363218 384170 363454
rect 384406 363218 384448 363454
rect 384128 363134 384448 363218
rect 384128 362898 384170 363134
rect 384406 362898 384448 363134
rect 384128 362866 384448 362898
rect 414848 363454 415168 363486
rect 414848 363218 414890 363454
rect 415126 363218 415168 363454
rect 414848 363134 415168 363218
rect 414848 362898 414890 363134
rect 415126 362898 415168 363134
rect 414848 362866 415168 362898
rect 445568 363454 445888 363486
rect 445568 363218 445610 363454
rect 445846 363218 445888 363454
rect 445568 363134 445888 363218
rect 445568 362898 445610 363134
rect 445846 362898 445888 363134
rect 445568 362866 445888 362898
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 61568 345454 61888 345486
rect 61568 345218 61610 345454
rect 61846 345218 61888 345454
rect 61568 345134 61888 345218
rect 61568 344898 61610 345134
rect 61846 344898 61888 345134
rect 61568 344866 61888 344898
rect 92288 345454 92608 345486
rect 92288 345218 92330 345454
rect 92566 345218 92608 345454
rect 92288 345134 92608 345218
rect 92288 344898 92330 345134
rect 92566 344898 92608 345134
rect 92288 344866 92608 344898
rect 123008 345454 123328 345486
rect 123008 345218 123050 345454
rect 123286 345218 123328 345454
rect 123008 345134 123328 345218
rect 123008 344898 123050 345134
rect 123286 344898 123328 345134
rect 123008 344866 123328 344898
rect 153728 345454 154048 345486
rect 153728 345218 153770 345454
rect 154006 345218 154048 345454
rect 153728 345134 154048 345218
rect 153728 344898 153770 345134
rect 154006 344898 154048 345134
rect 153728 344866 154048 344898
rect 184448 345454 184768 345486
rect 184448 345218 184490 345454
rect 184726 345218 184768 345454
rect 184448 345134 184768 345218
rect 184448 344898 184490 345134
rect 184726 344898 184768 345134
rect 184448 344866 184768 344898
rect 215168 345454 215488 345486
rect 215168 345218 215210 345454
rect 215446 345218 215488 345454
rect 215168 345134 215488 345218
rect 215168 344898 215210 345134
rect 215446 344898 215488 345134
rect 215168 344866 215488 344898
rect 245888 345454 246208 345486
rect 245888 345218 245930 345454
rect 246166 345218 246208 345454
rect 245888 345134 246208 345218
rect 245888 344898 245930 345134
rect 246166 344898 246208 345134
rect 245888 344866 246208 344898
rect 276608 345454 276928 345486
rect 276608 345218 276650 345454
rect 276886 345218 276928 345454
rect 276608 345134 276928 345218
rect 276608 344898 276650 345134
rect 276886 344898 276928 345134
rect 276608 344866 276928 344898
rect 307328 345454 307648 345486
rect 307328 345218 307370 345454
rect 307606 345218 307648 345454
rect 307328 345134 307648 345218
rect 307328 344898 307370 345134
rect 307606 344898 307648 345134
rect 307328 344866 307648 344898
rect 338048 345454 338368 345486
rect 338048 345218 338090 345454
rect 338326 345218 338368 345454
rect 338048 345134 338368 345218
rect 338048 344898 338090 345134
rect 338326 344898 338368 345134
rect 338048 344866 338368 344898
rect 368768 345454 369088 345486
rect 368768 345218 368810 345454
rect 369046 345218 369088 345454
rect 368768 345134 369088 345218
rect 368768 344898 368810 345134
rect 369046 344898 369088 345134
rect 368768 344866 369088 344898
rect 399488 345454 399808 345486
rect 399488 345218 399530 345454
rect 399766 345218 399808 345454
rect 399488 345134 399808 345218
rect 399488 344898 399530 345134
rect 399766 344898 399808 345134
rect 399488 344866 399808 344898
rect 430208 345454 430528 345486
rect 430208 345218 430250 345454
rect 430486 345218 430528 345454
rect 430208 345134 430528 345218
rect 430208 344898 430250 345134
rect 430486 344898 430528 345134
rect 430208 344866 430528 344898
rect 460928 345454 461248 345486
rect 460928 345218 460970 345454
rect 461206 345218 461248 345454
rect 460928 345134 461248 345218
rect 460928 344898 460970 345134
rect 461206 344898 461248 345134
rect 460928 344866 461248 344898
rect 76928 327454 77248 327486
rect 76928 327218 76970 327454
rect 77206 327218 77248 327454
rect 76928 327134 77248 327218
rect 76928 326898 76970 327134
rect 77206 326898 77248 327134
rect 76928 326866 77248 326898
rect 107648 327454 107968 327486
rect 107648 327218 107690 327454
rect 107926 327218 107968 327454
rect 107648 327134 107968 327218
rect 107648 326898 107690 327134
rect 107926 326898 107968 327134
rect 107648 326866 107968 326898
rect 138368 327454 138688 327486
rect 138368 327218 138410 327454
rect 138646 327218 138688 327454
rect 138368 327134 138688 327218
rect 138368 326898 138410 327134
rect 138646 326898 138688 327134
rect 138368 326866 138688 326898
rect 169088 327454 169408 327486
rect 169088 327218 169130 327454
rect 169366 327218 169408 327454
rect 169088 327134 169408 327218
rect 169088 326898 169130 327134
rect 169366 326898 169408 327134
rect 169088 326866 169408 326898
rect 199808 327454 200128 327486
rect 199808 327218 199850 327454
rect 200086 327218 200128 327454
rect 199808 327134 200128 327218
rect 199808 326898 199850 327134
rect 200086 326898 200128 327134
rect 199808 326866 200128 326898
rect 230528 327454 230848 327486
rect 230528 327218 230570 327454
rect 230806 327218 230848 327454
rect 230528 327134 230848 327218
rect 230528 326898 230570 327134
rect 230806 326898 230848 327134
rect 230528 326866 230848 326898
rect 261248 327454 261568 327486
rect 261248 327218 261290 327454
rect 261526 327218 261568 327454
rect 261248 327134 261568 327218
rect 261248 326898 261290 327134
rect 261526 326898 261568 327134
rect 261248 326866 261568 326898
rect 291968 327454 292288 327486
rect 291968 327218 292010 327454
rect 292246 327218 292288 327454
rect 291968 327134 292288 327218
rect 291968 326898 292010 327134
rect 292246 326898 292288 327134
rect 291968 326866 292288 326898
rect 322688 327454 323008 327486
rect 322688 327218 322730 327454
rect 322966 327218 323008 327454
rect 322688 327134 323008 327218
rect 322688 326898 322730 327134
rect 322966 326898 323008 327134
rect 322688 326866 323008 326898
rect 353408 327454 353728 327486
rect 353408 327218 353450 327454
rect 353686 327218 353728 327454
rect 353408 327134 353728 327218
rect 353408 326898 353450 327134
rect 353686 326898 353728 327134
rect 353408 326866 353728 326898
rect 384128 327454 384448 327486
rect 384128 327218 384170 327454
rect 384406 327218 384448 327454
rect 384128 327134 384448 327218
rect 384128 326898 384170 327134
rect 384406 326898 384448 327134
rect 384128 326866 384448 326898
rect 414848 327454 415168 327486
rect 414848 327218 414890 327454
rect 415126 327218 415168 327454
rect 414848 327134 415168 327218
rect 414848 326898 414890 327134
rect 415126 326898 415168 327134
rect 414848 326866 415168 326898
rect 445568 327454 445888 327486
rect 445568 327218 445610 327454
rect 445846 327218 445888 327454
rect 445568 327134 445888 327218
rect 445568 326898 445610 327134
rect 445846 326898 445888 327134
rect 445568 326866 445888 326898
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 61568 309454 61888 309486
rect 61568 309218 61610 309454
rect 61846 309218 61888 309454
rect 61568 309134 61888 309218
rect 61568 308898 61610 309134
rect 61846 308898 61888 309134
rect 61568 308866 61888 308898
rect 92288 309454 92608 309486
rect 92288 309218 92330 309454
rect 92566 309218 92608 309454
rect 92288 309134 92608 309218
rect 92288 308898 92330 309134
rect 92566 308898 92608 309134
rect 92288 308866 92608 308898
rect 123008 309454 123328 309486
rect 123008 309218 123050 309454
rect 123286 309218 123328 309454
rect 123008 309134 123328 309218
rect 123008 308898 123050 309134
rect 123286 308898 123328 309134
rect 123008 308866 123328 308898
rect 153728 309454 154048 309486
rect 153728 309218 153770 309454
rect 154006 309218 154048 309454
rect 153728 309134 154048 309218
rect 153728 308898 153770 309134
rect 154006 308898 154048 309134
rect 153728 308866 154048 308898
rect 184448 309454 184768 309486
rect 184448 309218 184490 309454
rect 184726 309218 184768 309454
rect 184448 309134 184768 309218
rect 184448 308898 184490 309134
rect 184726 308898 184768 309134
rect 184448 308866 184768 308898
rect 215168 309454 215488 309486
rect 215168 309218 215210 309454
rect 215446 309218 215488 309454
rect 215168 309134 215488 309218
rect 215168 308898 215210 309134
rect 215446 308898 215488 309134
rect 215168 308866 215488 308898
rect 245888 309454 246208 309486
rect 245888 309218 245930 309454
rect 246166 309218 246208 309454
rect 245888 309134 246208 309218
rect 245888 308898 245930 309134
rect 246166 308898 246208 309134
rect 245888 308866 246208 308898
rect 276608 309454 276928 309486
rect 276608 309218 276650 309454
rect 276886 309218 276928 309454
rect 276608 309134 276928 309218
rect 276608 308898 276650 309134
rect 276886 308898 276928 309134
rect 276608 308866 276928 308898
rect 307328 309454 307648 309486
rect 307328 309218 307370 309454
rect 307606 309218 307648 309454
rect 307328 309134 307648 309218
rect 307328 308898 307370 309134
rect 307606 308898 307648 309134
rect 307328 308866 307648 308898
rect 338048 309454 338368 309486
rect 338048 309218 338090 309454
rect 338326 309218 338368 309454
rect 338048 309134 338368 309218
rect 338048 308898 338090 309134
rect 338326 308898 338368 309134
rect 338048 308866 338368 308898
rect 368768 309454 369088 309486
rect 368768 309218 368810 309454
rect 369046 309218 369088 309454
rect 368768 309134 369088 309218
rect 368768 308898 368810 309134
rect 369046 308898 369088 309134
rect 368768 308866 369088 308898
rect 399488 309454 399808 309486
rect 399488 309218 399530 309454
rect 399766 309218 399808 309454
rect 399488 309134 399808 309218
rect 399488 308898 399530 309134
rect 399766 308898 399808 309134
rect 399488 308866 399808 308898
rect 430208 309454 430528 309486
rect 430208 309218 430250 309454
rect 430486 309218 430528 309454
rect 430208 309134 430528 309218
rect 430208 308898 430250 309134
rect 430486 308898 430528 309134
rect 430208 308866 430528 308898
rect 460928 309454 461248 309486
rect 460928 309218 460970 309454
rect 461206 309218 461248 309454
rect 460928 309134 461248 309218
rect 460928 308898 460970 309134
rect 461206 308898 461248 309134
rect 460928 308866 461248 308898
rect 76928 291454 77248 291486
rect 76928 291218 76970 291454
rect 77206 291218 77248 291454
rect 76928 291134 77248 291218
rect 76928 290898 76970 291134
rect 77206 290898 77248 291134
rect 76928 290866 77248 290898
rect 107648 291454 107968 291486
rect 107648 291218 107690 291454
rect 107926 291218 107968 291454
rect 107648 291134 107968 291218
rect 107648 290898 107690 291134
rect 107926 290898 107968 291134
rect 107648 290866 107968 290898
rect 138368 291454 138688 291486
rect 138368 291218 138410 291454
rect 138646 291218 138688 291454
rect 138368 291134 138688 291218
rect 138368 290898 138410 291134
rect 138646 290898 138688 291134
rect 138368 290866 138688 290898
rect 169088 291454 169408 291486
rect 169088 291218 169130 291454
rect 169366 291218 169408 291454
rect 169088 291134 169408 291218
rect 169088 290898 169130 291134
rect 169366 290898 169408 291134
rect 169088 290866 169408 290898
rect 199808 291454 200128 291486
rect 199808 291218 199850 291454
rect 200086 291218 200128 291454
rect 199808 291134 200128 291218
rect 199808 290898 199850 291134
rect 200086 290898 200128 291134
rect 199808 290866 200128 290898
rect 230528 291454 230848 291486
rect 230528 291218 230570 291454
rect 230806 291218 230848 291454
rect 230528 291134 230848 291218
rect 230528 290898 230570 291134
rect 230806 290898 230848 291134
rect 230528 290866 230848 290898
rect 261248 291454 261568 291486
rect 261248 291218 261290 291454
rect 261526 291218 261568 291454
rect 261248 291134 261568 291218
rect 261248 290898 261290 291134
rect 261526 290898 261568 291134
rect 261248 290866 261568 290898
rect 291968 291454 292288 291486
rect 291968 291218 292010 291454
rect 292246 291218 292288 291454
rect 291968 291134 292288 291218
rect 291968 290898 292010 291134
rect 292246 290898 292288 291134
rect 291968 290866 292288 290898
rect 322688 291454 323008 291486
rect 322688 291218 322730 291454
rect 322966 291218 323008 291454
rect 322688 291134 323008 291218
rect 322688 290898 322730 291134
rect 322966 290898 323008 291134
rect 322688 290866 323008 290898
rect 353408 291454 353728 291486
rect 353408 291218 353450 291454
rect 353686 291218 353728 291454
rect 353408 291134 353728 291218
rect 353408 290898 353450 291134
rect 353686 290898 353728 291134
rect 353408 290866 353728 290898
rect 384128 291454 384448 291486
rect 384128 291218 384170 291454
rect 384406 291218 384448 291454
rect 384128 291134 384448 291218
rect 384128 290898 384170 291134
rect 384406 290898 384448 291134
rect 384128 290866 384448 290898
rect 414848 291454 415168 291486
rect 414848 291218 414890 291454
rect 415126 291218 415168 291454
rect 414848 291134 415168 291218
rect 414848 290898 414890 291134
rect 415126 290898 415168 291134
rect 414848 290866 415168 290898
rect 445568 291454 445888 291486
rect 445568 291218 445610 291454
rect 445846 291218 445888 291454
rect 445568 291134 445888 291218
rect 445568 290898 445610 291134
rect 445846 290898 445888 291134
rect 445568 290866 445888 290898
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 61568 273454 61888 273486
rect 61568 273218 61610 273454
rect 61846 273218 61888 273454
rect 61568 273134 61888 273218
rect 61568 272898 61610 273134
rect 61846 272898 61888 273134
rect 61568 272866 61888 272898
rect 92288 273454 92608 273486
rect 92288 273218 92330 273454
rect 92566 273218 92608 273454
rect 92288 273134 92608 273218
rect 92288 272898 92330 273134
rect 92566 272898 92608 273134
rect 92288 272866 92608 272898
rect 123008 273454 123328 273486
rect 123008 273218 123050 273454
rect 123286 273218 123328 273454
rect 123008 273134 123328 273218
rect 123008 272898 123050 273134
rect 123286 272898 123328 273134
rect 123008 272866 123328 272898
rect 153728 273454 154048 273486
rect 153728 273218 153770 273454
rect 154006 273218 154048 273454
rect 153728 273134 154048 273218
rect 153728 272898 153770 273134
rect 154006 272898 154048 273134
rect 153728 272866 154048 272898
rect 184448 273454 184768 273486
rect 184448 273218 184490 273454
rect 184726 273218 184768 273454
rect 184448 273134 184768 273218
rect 184448 272898 184490 273134
rect 184726 272898 184768 273134
rect 184448 272866 184768 272898
rect 215168 273454 215488 273486
rect 215168 273218 215210 273454
rect 215446 273218 215488 273454
rect 215168 273134 215488 273218
rect 215168 272898 215210 273134
rect 215446 272898 215488 273134
rect 215168 272866 215488 272898
rect 245888 273454 246208 273486
rect 245888 273218 245930 273454
rect 246166 273218 246208 273454
rect 245888 273134 246208 273218
rect 245888 272898 245930 273134
rect 246166 272898 246208 273134
rect 245888 272866 246208 272898
rect 276608 273454 276928 273486
rect 276608 273218 276650 273454
rect 276886 273218 276928 273454
rect 276608 273134 276928 273218
rect 276608 272898 276650 273134
rect 276886 272898 276928 273134
rect 276608 272866 276928 272898
rect 307328 273454 307648 273486
rect 307328 273218 307370 273454
rect 307606 273218 307648 273454
rect 307328 273134 307648 273218
rect 307328 272898 307370 273134
rect 307606 272898 307648 273134
rect 307328 272866 307648 272898
rect 338048 273454 338368 273486
rect 338048 273218 338090 273454
rect 338326 273218 338368 273454
rect 338048 273134 338368 273218
rect 338048 272898 338090 273134
rect 338326 272898 338368 273134
rect 338048 272866 338368 272898
rect 368768 273454 369088 273486
rect 368768 273218 368810 273454
rect 369046 273218 369088 273454
rect 368768 273134 369088 273218
rect 368768 272898 368810 273134
rect 369046 272898 369088 273134
rect 368768 272866 369088 272898
rect 399488 273454 399808 273486
rect 399488 273218 399530 273454
rect 399766 273218 399808 273454
rect 399488 273134 399808 273218
rect 399488 272898 399530 273134
rect 399766 272898 399808 273134
rect 399488 272866 399808 272898
rect 430208 273454 430528 273486
rect 430208 273218 430250 273454
rect 430486 273218 430528 273454
rect 430208 273134 430528 273218
rect 430208 272898 430250 273134
rect 430486 272898 430528 273134
rect 430208 272866 430528 272898
rect 460928 273454 461248 273486
rect 460928 273218 460970 273454
rect 461206 273218 461248 273454
rect 460928 273134 461248 273218
rect 460928 272898 460970 273134
rect 461206 272898 461248 273134
rect 460928 272866 461248 272898
rect 76928 255454 77248 255486
rect 76928 255218 76970 255454
rect 77206 255218 77248 255454
rect 76928 255134 77248 255218
rect 76928 254898 76970 255134
rect 77206 254898 77248 255134
rect 76928 254866 77248 254898
rect 107648 255454 107968 255486
rect 107648 255218 107690 255454
rect 107926 255218 107968 255454
rect 107648 255134 107968 255218
rect 107648 254898 107690 255134
rect 107926 254898 107968 255134
rect 107648 254866 107968 254898
rect 138368 255454 138688 255486
rect 138368 255218 138410 255454
rect 138646 255218 138688 255454
rect 138368 255134 138688 255218
rect 138368 254898 138410 255134
rect 138646 254898 138688 255134
rect 138368 254866 138688 254898
rect 169088 255454 169408 255486
rect 169088 255218 169130 255454
rect 169366 255218 169408 255454
rect 169088 255134 169408 255218
rect 169088 254898 169130 255134
rect 169366 254898 169408 255134
rect 169088 254866 169408 254898
rect 199808 255454 200128 255486
rect 199808 255218 199850 255454
rect 200086 255218 200128 255454
rect 199808 255134 200128 255218
rect 199808 254898 199850 255134
rect 200086 254898 200128 255134
rect 199808 254866 200128 254898
rect 230528 255454 230848 255486
rect 230528 255218 230570 255454
rect 230806 255218 230848 255454
rect 230528 255134 230848 255218
rect 230528 254898 230570 255134
rect 230806 254898 230848 255134
rect 230528 254866 230848 254898
rect 261248 255454 261568 255486
rect 261248 255218 261290 255454
rect 261526 255218 261568 255454
rect 261248 255134 261568 255218
rect 261248 254898 261290 255134
rect 261526 254898 261568 255134
rect 261248 254866 261568 254898
rect 291968 255454 292288 255486
rect 291968 255218 292010 255454
rect 292246 255218 292288 255454
rect 291968 255134 292288 255218
rect 291968 254898 292010 255134
rect 292246 254898 292288 255134
rect 291968 254866 292288 254898
rect 322688 255454 323008 255486
rect 322688 255218 322730 255454
rect 322966 255218 323008 255454
rect 322688 255134 323008 255218
rect 322688 254898 322730 255134
rect 322966 254898 323008 255134
rect 322688 254866 323008 254898
rect 353408 255454 353728 255486
rect 353408 255218 353450 255454
rect 353686 255218 353728 255454
rect 353408 255134 353728 255218
rect 353408 254898 353450 255134
rect 353686 254898 353728 255134
rect 353408 254866 353728 254898
rect 384128 255454 384448 255486
rect 384128 255218 384170 255454
rect 384406 255218 384448 255454
rect 384128 255134 384448 255218
rect 384128 254898 384170 255134
rect 384406 254898 384448 255134
rect 384128 254866 384448 254898
rect 414848 255454 415168 255486
rect 414848 255218 414890 255454
rect 415126 255218 415168 255454
rect 414848 255134 415168 255218
rect 414848 254898 414890 255134
rect 415126 254898 415168 255134
rect 414848 254866 415168 254898
rect 445568 255454 445888 255486
rect 445568 255218 445610 255454
rect 445846 255218 445888 255454
rect 445568 255134 445888 255218
rect 445568 254898 445610 255134
rect 445846 254898 445888 255134
rect 445568 254866 445888 254898
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 61568 237454 61888 237486
rect 61568 237218 61610 237454
rect 61846 237218 61888 237454
rect 61568 237134 61888 237218
rect 61568 236898 61610 237134
rect 61846 236898 61888 237134
rect 61568 236866 61888 236898
rect 92288 237454 92608 237486
rect 92288 237218 92330 237454
rect 92566 237218 92608 237454
rect 92288 237134 92608 237218
rect 92288 236898 92330 237134
rect 92566 236898 92608 237134
rect 92288 236866 92608 236898
rect 123008 237454 123328 237486
rect 123008 237218 123050 237454
rect 123286 237218 123328 237454
rect 123008 237134 123328 237218
rect 123008 236898 123050 237134
rect 123286 236898 123328 237134
rect 123008 236866 123328 236898
rect 153728 237454 154048 237486
rect 153728 237218 153770 237454
rect 154006 237218 154048 237454
rect 153728 237134 154048 237218
rect 153728 236898 153770 237134
rect 154006 236898 154048 237134
rect 153728 236866 154048 236898
rect 184448 237454 184768 237486
rect 184448 237218 184490 237454
rect 184726 237218 184768 237454
rect 184448 237134 184768 237218
rect 184448 236898 184490 237134
rect 184726 236898 184768 237134
rect 184448 236866 184768 236898
rect 215168 237454 215488 237486
rect 215168 237218 215210 237454
rect 215446 237218 215488 237454
rect 215168 237134 215488 237218
rect 215168 236898 215210 237134
rect 215446 236898 215488 237134
rect 215168 236866 215488 236898
rect 245888 237454 246208 237486
rect 245888 237218 245930 237454
rect 246166 237218 246208 237454
rect 245888 237134 246208 237218
rect 245888 236898 245930 237134
rect 246166 236898 246208 237134
rect 245888 236866 246208 236898
rect 276608 237454 276928 237486
rect 276608 237218 276650 237454
rect 276886 237218 276928 237454
rect 276608 237134 276928 237218
rect 276608 236898 276650 237134
rect 276886 236898 276928 237134
rect 276608 236866 276928 236898
rect 307328 237454 307648 237486
rect 307328 237218 307370 237454
rect 307606 237218 307648 237454
rect 307328 237134 307648 237218
rect 307328 236898 307370 237134
rect 307606 236898 307648 237134
rect 307328 236866 307648 236898
rect 338048 237454 338368 237486
rect 338048 237218 338090 237454
rect 338326 237218 338368 237454
rect 338048 237134 338368 237218
rect 338048 236898 338090 237134
rect 338326 236898 338368 237134
rect 338048 236866 338368 236898
rect 368768 237454 369088 237486
rect 368768 237218 368810 237454
rect 369046 237218 369088 237454
rect 368768 237134 369088 237218
rect 368768 236898 368810 237134
rect 369046 236898 369088 237134
rect 368768 236866 369088 236898
rect 399488 237454 399808 237486
rect 399488 237218 399530 237454
rect 399766 237218 399808 237454
rect 399488 237134 399808 237218
rect 399488 236898 399530 237134
rect 399766 236898 399808 237134
rect 399488 236866 399808 236898
rect 430208 237454 430528 237486
rect 430208 237218 430250 237454
rect 430486 237218 430528 237454
rect 430208 237134 430528 237218
rect 430208 236898 430250 237134
rect 430486 236898 430528 237134
rect 430208 236866 430528 236898
rect 460928 237454 461248 237486
rect 460928 237218 460970 237454
rect 461206 237218 461248 237454
rect 460928 237134 461248 237218
rect 460928 236898 460970 237134
rect 461206 236898 461248 237134
rect 460928 236866 461248 236898
rect 76928 219454 77248 219486
rect 76928 219218 76970 219454
rect 77206 219218 77248 219454
rect 76928 219134 77248 219218
rect 76928 218898 76970 219134
rect 77206 218898 77248 219134
rect 76928 218866 77248 218898
rect 107648 219454 107968 219486
rect 107648 219218 107690 219454
rect 107926 219218 107968 219454
rect 107648 219134 107968 219218
rect 107648 218898 107690 219134
rect 107926 218898 107968 219134
rect 107648 218866 107968 218898
rect 138368 219454 138688 219486
rect 138368 219218 138410 219454
rect 138646 219218 138688 219454
rect 138368 219134 138688 219218
rect 138368 218898 138410 219134
rect 138646 218898 138688 219134
rect 138368 218866 138688 218898
rect 169088 219454 169408 219486
rect 169088 219218 169130 219454
rect 169366 219218 169408 219454
rect 169088 219134 169408 219218
rect 169088 218898 169130 219134
rect 169366 218898 169408 219134
rect 169088 218866 169408 218898
rect 199808 219454 200128 219486
rect 199808 219218 199850 219454
rect 200086 219218 200128 219454
rect 199808 219134 200128 219218
rect 199808 218898 199850 219134
rect 200086 218898 200128 219134
rect 199808 218866 200128 218898
rect 230528 219454 230848 219486
rect 230528 219218 230570 219454
rect 230806 219218 230848 219454
rect 230528 219134 230848 219218
rect 230528 218898 230570 219134
rect 230806 218898 230848 219134
rect 230528 218866 230848 218898
rect 261248 219454 261568 219486
rect 261248 219218 261290 219454
rect 261526 219218 261568 219454
rect 261248 219134 261568 219218
rect 261248 218898 261290 219134
rect 261526 218898 261568 219134
rect 261248 218866 261568 218898
rect 291968 219454 292288 219486
rect 291968 219218 292010 219454
rect 292246 219218 292288 219454
rect 291968 219134 292288 219218
rect 291968 218898 292010 219134
rect 292246 218898 292288 219134
rect 291968 218866 292288 218898
rect 322688 219454 323008 219486
rect 322688 219218 322730 219454
rect 322966 219218 323008 219454
rect 322688 219134 323008 219218
rect 322688 218898 322730 219134
rect 322966 218898 323008 219134
rect 322688 218866 323008 218898
rect 353408 219454 353728 219486
rect 353408 219218 353450 219454
rect 353686 219218 353728 219454
rect 353408 219134 353728 219218
rect 353408 218898 353450 219134
rect 353686 218898 353728 219134
rect 353408 218866 353728 218898
rect 384128 219454 384448 219486
rect 384128 219218 384170 219454
rect 384406 219218 384448 219454
rect 384128 219134 384448 219218
rect 384128 218898 384170 219134
rect 384406 218898 384448 219134
rect 384128 218866 384448 218898
rect 414848 219454 415168 219486
rect 414848 219218 414890 219454
rect 415126 219218 415168 219454
rect 414848 219134 415168 219218
rect 414848 218898 414890 219134
rect 415126 218898 415168 219134
rect 414848 218866 415168 218898
rect 445568 219454 445888 219486
rect 445568 219218 445610 219454
rect 445846 219218 445888 219454
rect 445568 219134 445888 219218
rect 445568 218898 445610 219134
rect 445846 218898 445888 219134
rect 445568 218866 445888 218898
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 61568 201454 61888 201486
rect 61568 201218 61610 201454
rect 61846 201218 61888 201454
rect 61568 201134 61888 201218
rect 61568 200898 61610 201134
rect 61846 200898 61888 201134
rect 61568 200866 61888 200898
rect 92288 201454 92608 201486
rect 92288 201218 92330 201454
rect 92566 201218 92608 201454
rect 92288 201134 92608 201218
rect 92288 200898 92330 201134
rect 92566 200898 92608 201134
rect 92288 200866 92608 200898
rect 123008 201454 123328 201486
rect 123008 201218 123050 201454
rect 123286 201218 123328 201454
rect 123008 201134 123328 201218
rect 123008 200898 123050 201134
rect 123286 200898 123328 201134
rect 123008 200866 123328 200898
rect 153728 201454 154048 201486
rect 153728 201218 153770 201454
rect 154006 201218 154048 201454
rect 153728 201134 154048 201218
rect 153728 200898 153770 201134
rect 154006 200898 154048 201134
rect 153728 200866 154048 200898
rect 184448 201454 184768 201486
rect 184448 201218 184490 201454
rect 184726 201218 184768 201454
rect 184448 201134 184768 201218
rect 184448 200898 184490 201134
rect 184726 200898 184768 201134
rect 184448 200866 184768 200898
rect 215168 201454 215488 201486
rect 215168 201218 215210 201454
rect 215446 201218 215488 201454
rect 215168 201134 215488 201218
rect 215168 200898 215210 201134
rect 215446 200898 215488 201134
rect 215168 200866 215488 200898
rect 245888 201454 246208 201486
rect 245888 201218 245930 201454
rect 246166 201218 246208 201454
rect 245888 201134 246208 201218
rect 245888 200898 245930 201134
rect 246166 200898 246208 201134
rect 245888 200866 246208 200898
rect 276608 201454 276928 201486
rect 276608 201218 276650 201454
rect 276886 201218 276928 201454
rect 276608 201134 276928 201218
rect 276608 200898 276650 201134
rect 276886 200898 276928 201134
rect 276608 200866 276928 200898
rect 307328 201454 307648 201486
rect 307328 201218 307370 201454
rect 307606 201218 307648 201454
rect 307328 201134 307648 201218
rect 307328 200898 307370 201134
rect 307606 200898 307648 201134
rect 307328 200866 307648 200898
rect 338048 201454 338368 201486
rect 338048 201218 338090 201454
rect 338326 201218 338368 201454
rect 338048 201134 338368 201218
rect 338048 200898 338090 201134
rect 338326 200898 338368 201134
rect 338048 200866 338368 200898
rect 368768 201454 369088 201486
rect 368768 201218 368810 201454
rect 369046 201218 369088 201454
rect 368768 201134 369088 201218
rect 368768 200898 368810 201134
rect 369046 200898 369088 201134
rect 368768 200866 369088 200898
rect 399488 201454 399808 201486
rect 399488 201218 399530 201454
rect 399766 201218 399808 201454
rect 399488 201134 399808 201218
rect 399488 200898 399530 201134
rect 399766 200898 399808 201134
rect 399488 200866 399808 200898
rect 430208 201454 430528 201486
rect 430208 201218 430250 201454
rect 430486 201218 430528 201454
rect 430208 201134 430528 201218
rect 430208 200898 430250 201134
rect 430486 200898 430528 201134
rect 430208 200866 430528 200898
rect 460928 201454 461248 201486
rect 460928 201218 460970 201454
rect 461206 201218 461248 201454
rect 460928 201134 461248 201218
rect 460928 200898 460970 201134
rect 461206 200898 461248 201134
rect 460928 200866 461248 200898
rect 76928 183454 77248 183486
rect 76928 183218 76970 183454
rect 77206 183218 77248 183454
rect 76928 183134 77248 183218
rect 76928 182898 76970 183134
rect 77206 182898 77248 183134
rect 76928 182866 77248 182898
rect 107648 183454 107968 183486
rect 107648 183218 107690 183454
rect 107926 183218 107968 183454
rect 107648 183134 107968 183218
rect 107648 182898 107690 183134
rect 107926 182898 107968 183134
rect 107648 182866 107968 182898
rect 138368 183454 138688 183486
rect 138368 183218 138410 183454
rect 138646 183218 138688 183454
rect 138368 183134 138688 183218
rect 138368 182898 138410 183134
rect 138646 182898 138688 183134
rect 138368 182866 138688 182898
rect 169088 183454 169408 183486
rect 169088 183218 169130 183454
rect 169366 183218 169408 183454
rect 169088 183134 169408 183218
rect 169088 182898 169130 183134
rect 169366 182898 169408 183134
rect 169088 182866 169408 182898
rect 199808 183454 200128 183486
rect 199808 183218 199850 183454
rect 200086 183218 200128 183454
rect 199808 183134 200128 183218
rect 199808 182898 199850 183134
rect 200086 182898 200128 183134
rect 199808 182866 200128 182898
rect 230528 183454 230848 183486
rect 230528 183218 230570 183454
rect 230806 183218 230848 183454
rect 230528 183134 230848 183218
rect 230528 182898 230570 183134
rect 230806 182898 230848 183134
rect 230528 182866 230848 182898
rect 261248 183454 261568 183486
rect 261248 183218 261290 183454
rect 261526 183218 261568 183454
rect 261248 183134 261568 183218
rect 261248 182898 261290 183134
rect 261526 182898 261568 183134
rect 261248 182866 261568 182898
rect 291968 183454 292288 183486
rect 291968 183218 292010 183454
rect 292246 183218 292288 183454
rect 291968 183134 292288 183218
rect 291968 182898 292010 183134
rect 292246 182898 292288 183134
rect 291968 182866 292288 182898
rect 322688 183454 323008 183486
rect 322688 183218 322730 183454
rect 322966 183218 323008 183454
rect 322688 183134 323008 183218
rect 322688 182898 322730 183134
rect 322966 182898 323008 183134
rect 322688 182866 323008 182898
rect 353408 183454 353728 183486
rect 353408 183218 353450 183454
rect 353686 183218 353728 183454
rect 353408 183134 353728 183218
rect 353408 182898 353450 183134
rect 353686 182898 353728 183134
rect 353408 182866 353728 182898
rect 384128 183454 384448 183486
rect 384128 183218 384170 183454
rect 384406 183218 384448 183454
rect 384128 183134 384448 183218
rect 384128 182898 384170 183134
rect 384406 182898 384448 183134
rect 384128 182866 384448 182898
rect 414848 183454 415168 183486
rect 414848 183218 414890 183454
rect 415126 183218 415168 183454
rect 414848 183134 415168 183218
rect 414848 182898 414890 183134
rect 415126 182898 415168 183134
rect 414848 182866 415168 182898
rect 445568 183454 445888 183486
rect 445568 183218 445610 183454
rect 445846 183218 445888 183454
rect 445568 183134 445888 183218
rect 445568 182898 445610 183134
rect 445846 182898 445888 183134
rect 445568 182866 445888 182898
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 61568 165454 61888 165486
rect 61568 165218 61610 165454
rect 61846 165218 61888 165454
rect 61568 165134 61888 165218
rect 61568 164898 61610 165134
rect 61846 164898 61888 165134
rect 61568 164866 61888 164898
rect 92288 165454 92608 165486
rect 92288 165218 92330 165454
rect 92566 165218 92608 165454
rect 92288 165134 92608 165218
rect 92288 164898 92330 165134
rect 92566 164898 92608 165134
rect 92288 164866 92608 164898
rect 123008 165454 123328 165486
rect 123008 165218 123050 165454
rect 123286 165218 123328 165454
rect 123008 165134 123328 165218
rect 123008 164898 123050 165134
rect 123286 164898 123328 165134
rect 123008 164866 123328 164898
rect 153728 165454 154048 165486
rect 153728 165218 153770 165454
rect 154006 165218 154048 165454
rect 153728 165134 154048 165218
rect 153728 164898 153770 165134
rect 154006 164898 154048 165134
rect 153728 164866 154048 164898
rect 184448 165454 184768 165486
rect 184448 165218 184490 165454
rect 184726 165218 184768 165454
rect 184448 165134 184768 165218
rect 184448 164898 184490 165134
rect 184726 164898 184768 165134
rect 184448 164866 184768 164898
rect 215168 165454 215488 165486
rect 215168 165218 215210 165454
rect 215446 165218 215488 165454
rect 215168 165134 215488 165218
rect 215168 164898 215210 165134
rect 215446 164898 215488 165134
rect 215168 164866 215488 164898
rect 245888 165454 246208 165486
rect 245888 165218 245930 165454
rect 246166 165218 246208 165454
rect 245888 165134 246208 165218
rect 245888 164898 245930 165134
rect 246166 164898 246208 165134
rect 245888 164866 246208 164898
rect 276608 165454 276928 165486
rect 276608 165218 276650 165454
rect 276886 165218 276928 165454
rect 276608 165134 276928 165218
rect 276608 164898 276650 165134
rect 276886 164898 276928 165134
rect 276608 164866 276928 164898
rect 307328 165454 307648 165486
rect 307328 165218 307370 165454
rect 307606 165218 307648 165454
rect 307328 165134 307648 165218
rect 307328 164898 307370 165134
rect 307606 164898 307648 165134
rect 307328 164866 307648 164898
rect 338048 165454 338368 165486
rect 338048 165218 338090 165454
rect 338326 165218 338368 165454
rect 338048 165134 338368 165218
rect 338048 164898 338090 165134
rect 338326 164898 338368 165134
rect 338048 164866 338368 164898
rect 368768 165454 369088 165486
rect 368768 165218 368810 165454
rect 369046 165218 369088 165454
rect 368768 165134 369088 165218
rect 368768 164898 368810 165134
rect 369046 164898 369088 165134
rect 368768 164866 369088 164898
rect 399488 165454 399808 165486
rect 399488 165218 399530 165454
rect 399766 165218 399808 165454
rect 399488 165134 399808 165218
rect 399488 164898 399530 165134
rect 399766 164898 399808 165134
rect 399488 164866 399808 164898
rect 430208 165454 430528 165486
rect 430208 165218 430250 165454
rect 430486 165218 430528 165454
rect 430208 165134 430528 165218
rect 430208 164898 430250 165134
rect 430486 164898 430528 165134
rect 430208 164866 430528 164898
rect 460928 165454 461248 165486
rect 460928 165218 460970 165454
rect 461206 165218 461248 165454
rect 460928 165134 461248 165218
rect 460928 164898 460970 165134
rect 461206 164898 461248 165134
rect 460928 164866 461248 164898
rect 76928 147454 77248 147486
rect 76928 147218 76970 147454
rect 77206 147218 77248 147454
rect 76928 147134 77248 147218
rect 76928 146898 76970 147134
rect 77206 146898 77248 147134
rect 76928 146866 77248 146898
rect 107648 147454 107968 147486
rect 107648 147218 107690 147454
rect 107926 147218 107968 147454
rect 107648 147134 107968 147218
rect 107648 146898 107690 147134
rect 107926 146898 107968 147134
rect 107648 146866 107968 146898
rect 138368 147454 138688 147486
rect 138368 147218 138410 147454
rect 138646 147218 138688 147454
rect 138368 147134 138688 147218
rect 138368 146898 138410 147134
rect 138646 146898 138688 147134
rect 138368 146866 138688 146898
rect 169088 147454 169408 147486
rect 169088 147218 169130 147454
rect 169366 147218 169408 147454
rect 169088 147134 169408 147218
rect 169088 146898 169130 147134
rect 169366 146898 169408 147134
rect 169088 146866 169408 146898
rect 199808 147454 200128 147486
rect 199808 147218 199850 147454
rect 200086 147218 200128 147454
rect 199808 147134 200128 147218
rect 199808 146898 199850 147134
rect 200086 146898 200128 147134
rect 199808 146866 200128 146898
rect 230528 147454 230848 147486
rect 230528 147218 230570 147454
rect 230806 147218 230848 147454
rect 230528 147134 230848 147218
rect 230528 146898 230570 147134
rect 230806 146898 230848 147134
rect 230528 146866 230848 146898
rect 261248 147454 261568 147486
rect 261248 147218 261290 147454
rect 261526 147218 261568 147454
rect 261248 147134 261568 147218
rect 261248 146898 261290 147134
rect 261526 146898 261568 147134
rect 261248 146866 261568 146898
rect 291968 147454 292288 147486
rect 291968 147218 292010 147454
rect 292246 147218 292288 147454
rect 291968 147134 292288 147218
rect 291968 146898 292010 147134
rect 292246 146898 292288 147134
rect 291968 146866 292288 146898
rect 322688 147454 323008 147486
rect 322688 147218 322730 147454
rect 322966 147218 323008 147454
rect 322688 147134 323008 147218
rect 322688 146898 322730 147134
rect 322966 146898 323008 147134
rect 322688 146866 323008 146898
rect 353408 147454 353728 147486
rect 353408 147218 353450 147454
rect 353686 147218 353728 147454
rect 353408 147134 353728 147218
rect 353408 146898 353450 147134
rect 353686 146898 353728 147134
rect 353408 146866 353728 146898
rect 384128 147454 384448 147486
rect 384128 147218 384170 147454
rect 384406 147218 384448 147454
rect 384128 147134 384448 147218
rect 384128 146898 384170 147134
rect 384406 146898 384448 147134
rect 384128 146866 384448 146898
rect 414848 147454 415168 147486
rect 414848 147218 414890 147454
rect 415126 147218 415168 147454
rect 414848 147134 415168 147218
rect 414848 146898 414890 147134
rect 415126 146898 415168 147134
rect 414848 146866 415168 146898
rect 445568 147454 445888 147486
rect 445568 147218 445610 147454
rect 445846 147218 445888 147454
rect 445568 147134 445888 147218
rect 445568 146898 445610 147134
rect 445846 146898 445888 147134
rect 445568 146866 445888 146898
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 61568 129454 61888 129486
rect 61568 129218 61610 129454
rect 61846 129218 61888 129454
rect 61568 129134 61888 129218
rect 61568 128898 61610 129134
rect 61846 128898 61888 129134
rect 61568 128866 61888 128898
rect 92288 129454 92608 129486
rect 92288 129218 92330 129454
rect 92566 129218 92608 129454
rect 92288 129134 92608 129218
rect 92288 128898 92330 129134
rect 92566 128898 92608 129134
rect 92288 128866 92608 128898
rect 123008 129454 123328 129486
rect 123008 129218 123050 129454
rect 123286 129218 123328 129454
rect 123008 129134 123328 129218
rect 123008 128898 123050 129134
rect 123286 128898 123328 129134
rect 123008 128866 123328 128898
rect 153728 129454 154048 129486
rect 153728 129218 153770 129454
rect 154006 129218 154048 129454
rect 153728 129134 154048 129218
rect 153728 128898 153770 129134
rect 154006 128898 154048 129134
rect 153728 128866 154048 128898
rect 184448 129454 184768 129486
rect 184448 129218 184490 129454
rect 184726 129218 184768 129454
rect 184448 129134 184768 129218
rect 184448 128898 184490 129134
rect 184726 128898 184768 129134
rect 184448 128866 184768 128898
rect 215168 129454 215488 129486
rect 215168 129218 215210 129454
rect 215446 129218 215488 129454
rect 215168 129134 215488 129218
rect 215168 128898 215210 129134
rect 215446 128898 215488 129134
rect 215168 128866 215488 128898
rect 245888 129454 246208 129486
rect 245888 129218 245930 129454
rect 246166 129218 246208 129454
rect 245888 129134 246208 129218
rect 245888 128898 245930 129134
rect 246166 128898 246208 129134
rect 245888 128866 246208 128898
rect 276608 129454 276928 129486
rect 276608 129218 276650 129454
rect 276886 129218 276928 129454
rect 276608 129134 276928 129218
rect 276608 128898 276650 129134
rect 276886 128898 276928 129134
rect 276608 128866 276928 128898
rect 307328 129454 307648 129486
rect 307328 129218 307370 129454
rect 307606 129218 307648 129454
rect 307328 129134 307648 129218
rect 307328 128898 307370 129134
rect 307606 128898 307648 129134
rect 307328 128866 307648 128898
rect 338048 129454 338368 129486
rect 338048 129218 338090 129454
rect 338326 129218 338368 129454
rect 338048 129134 338368 129218
rect 338048 128898 338090 129134
rect 338326 128898 338368 129134
rect 338048 128866 338368 128898
rect 368768 129454 369088 129486
rect 368768 129218 368810 129454
rect 369046 129218 369088 129454
rect 368768 129134 369088 129218
rect 368768 128898 368810 129134
rect 369046 128898 369088 129134
rect 368768 128866 369088 128898
rect 399488 129454 399808 129486
rect 399488 129218 399530 129454
rect 399766 129218 399808 129454
rect 399488 129134 399808 129218
rect 399488 128898 399530 129134
rect 399766 128898 399808 129134
rect 399488 128866 399808 128898
rect 430208 129454 430528 129486
rect 430208 129218 430250 129454
rect 430486 129218 430528 129454
rect 430208 129134 430528 129218
rect 430208 128898 430250 129134
rect 430486 128898 430528 129134
rect 430208 128866 430528 128898
rect 460928 129454 461248 129486
rect 460928 129218 460970 129454
rect 461206 129218 461248 129454
rect 460928 129134 461248 129218
rect 460928 128898 460970 129134
rect 461206 128898 461248 129134
rect 460928 128866 461248 128898
rect 76928 111454 77248 111486
rect 76928 111218 76970 111454
rect 77206 111218 77248 111454
rect 76928 111134 77248 111218
rect 76928 110898 76970 111134
rect 77206 110898 77248 111134
rect 76928 110866 77248 110898
rect 107648 111454 107968 111486
rect 107648 111218 107690 111454
rect 107926 111218 107968 111454
rect 107648 111134 107968 111218
rect 107648 110898 107690 111134
rect 107926 110898 107968 111134
rect 107648 110866 107968 110898
rect 138368 111454 138688 111486
rect 138368 111218 138410 111454
rect 138646 111218 138688 111454
rect 138368 111134 138688 111218
rect 138368 110898 138410 111134
rect 138646 110898 138688 111134
rect 138368 110866 138688 110898
rect 169088 111454 169408 111486
rect 169088 111218 169130 111454
rect 169366 111218 169408 111454
rect 169088 111134 169408 111218
rect 169088 110898 169130 111134
rect 169366 110898 169408 111134
rect 169088 110866 169408 110898
rect 199808 111454 200128 111486
rect 199808 111218 199850 111454
rect 200086 111218 200128 111454
rect 199808 111134 200128 111218
rect 199808 110898 199850 111134
rect 200086 110898 200128 111134
rect 199808 110866 200128 110898
rect 230528 111454 230848 111486
rect 230528 111218 230570 111454
rect 230806 111218 230848 111454
rect 230528 111134 230848 111218
rect 230528 110898 230570 111134
rect 230806 110898 230848 111134
rect 230528 110866 230848 110898
rect 261248 111454 261568 111486
rect 261248 111218 261290 111454
rect 261526 111218 261568 111454
rect 261248 111134 261568 111218
rect 261248 110898 261290 111134
rect 261526 110898 261568 111134
rect 261248 110866 261568 110898
rect 291968 111454 292288 111486
rect 291968 111218 292010 111454
rect 292246 111218 292288 111454
rect 291968 111134 292288 111218
rect 291968 110898 292010 111134
rect 292246 110898 292288 111134
rect 291968 110866 292288 110898
rect 322688 111454 323008 111486
rect 322688 111218 322730 111454
rect 322966 111218 323008 111454
rect 322688 111134 323008 111218
rect 322688 110898 322730 111134
rect 322966 110898 323008 111134
rect 322688 110866 323008 110898
rect 353408 111454 353728 111486
rect 353408 111218 353450 111454
rect 353686 111218 353728 111454
rect 353408 111134 353728 111218
rect 353408 110898 353450 111134
rect 353686 110898 353728 111134
rect 353408 110866 353728 110898
rect 384128 111454 384448 111486
rect 384128 111218 384170 111454
rect 384406 111218 384448 111454
rect 384128 111134 384448 111218
rect 384128 110898 384170 111134
rect 384406 110898 384448 111134
rect 384128 110866 384448 110898
rect 414848 111454 415168 111486
rect 414848 111218 414890 111454
rect 415126 111218 415168 111454
rect 414848 111134 415168 111218
rect 414848 110898 414890 111134
rect 415126 110898 415168 111134
rect 414848 110866 415168 110898
rect 445568 111454 445888 111486
rect 445568 111218 445610 111454
rect 445846 111218 445888 111454
rect 445568 111134 445888 111218
rect 445568 110898 445610 111134
rect 445846 110898 445888 111134
rect 445568 110866 445888 110898
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 61568 93454 61888 93486
rect 61568 93218 61610 93454
rect 61846 93218 61888 93454
rect 61568 93134 61888 93218
rect 61568 92898 61610 93134
rect 61846 92898 61888 93134
rect 61568 92866 61888 92898
rect 92288 93454 92608 93486
rect 92288 93218 92330 93454
rect 92566 93218 92608 93454
rect 92288 93134 92608 93218
rect 92288 92898 92330 93134
rect 92566 92898 92608 93134
rect 92288 92866 92608 92898
rect 123008 93454 123328 93486
rect 123008 93218 123050 93454
rect 123286 93218 123328 93454
rect 123008 93134 123328 93218
rect 123008 92898 123050 93134
rect 123286 92898 123328 93134
rect 123008 92866 123328 92898
rect 153728 93454 154048 93486
rect 153728 93218 153770 93454
rect 154006 93218 154048 93454
rect 153728 93134 154048 93218
rect 153728 92898 153770 93134
rect 154006 92898 154048 93134
rect 153728 92866 154048 92898
rect 184448 93454 184768 93486
rect 184448 93218 184490 93454
rect 184726 93218 184768 93454
rect 184448 93134 184768 93218
rect 184448 92898 184490 93134
rect 184726 92898 184768 93134
rect 184448 92866 184768 92898
rect 215168 93454 215488 93486
rect 215168 93218 215210 93454
rect 215446 93218 215488 93454
rect 215168 93134 215488 93218
rect 215168 92898 215210 93134
rect 215446 92898 215488 93134
rect 215168 92866 215488 92898
rect 245888 93454 246208 93486
rect 245888 93218 245930 93454
rect 246166 93218 246208 93454
rect 245888 93134 246208 93218
rect 245888 92898 245930 93134
rect 246166 92898 246208 93134
rect 245888 92866 246208 92898
rect 276608 93454 276928 93486
rect 276608 93218 276650 93454
rect 276886 93218 276928 93454
rect 276608 93134 276928 93218
rect 276608 92898 276650 93134
rect 276886 92898 276928 93134
rect 276608 92866 276928 92898
rect 307328 93454 307648 93486
rect 307328 93218 307370 93454
rect 307606 93218 307648 93454
rect 307328 93134 307648 93218
rect 307328 92898 307370 93134
rect 307606 92898 307648 93134
rect 307328 92866 307648 92898
rect 338048 93454 338368 93486
rect 338048 93218 338090 93454
rect 338326 93218 338368 93454
rect 338048 93134 338368 93218
rect 338048 92898 338090 93134
rect 338326 92898 338368 93134
rect 338048 92866 338368 92898
rect 368768 93454 369088 93486
rect 368768 93218 368810 93454
rect 369046 93218 369088 93454
rect 368768 93134 369088 93218
rect 368768 92898 368810 93134
rect 369046 92898 369088 93134
rect 368768 92866 369088 92898
rect 399488 93454 399808 93486
rect 399488 93218 399530 93454
rect 399766 93218 399808 93454
rect 399488 93134 399808 93218
rect 399488 92898 399530 93134
rect 399766 92898 399808 93134
rect 399488 92866 399808 92898
rect 430208 93454 430528 93486
rect 430208 93218 430250 93454
rect 430486 93218 430528 93454
rect 430208 93134 430528 93218
rect 430208 92898 430250 93134
rect 430486 92898 430528 93134
rect 430208 92866 430528 92898
rect 460928 93454 461248 93486
rect 460928 93218 460970 93454
rect 461206 93218 461248 93454
rect 460928 93134 461248 93218
rect 460928 92898 460970 93134
rect 461206 92898 461248 93134
rect 460928 92866 461248 92898
rect 76928 75454 77248 75486
rect 76928 75218 76970 75454
rect 77206 75218 77248 75454
rect 76928 75134 77248 75218
rect 76928 74898 76970 75134
rect 77206 74898 77248 75134
rect 76928 74866 77248 74898
rect 107648 75454 107968 75486
rect 107648 75218 107690 75454
rect 107926 75218 107968 75454
rect 107648 75134 107968 75218
rect 107648 74898 107690 75134
rect 107926 74898 107968 75134
rect 107648 74866 107968 74898
rect 138368 75454 138688 75486
rect 138368 75218 138410 75454
rect 138646 75218 138688 75454
rect 138368 75134 138688 75218
rect 138368 74898 138410 75134
rect 138646 74898 138688 75134
rect 138368 74866 138688 74898
rect 169088 75454 169408 75486
rect 169088 75218 169130 75454
rect 169366 75218 169408 75454
rect 169088 75134 169408 75218
rect 169088 74898 169130 75134
rect 169366 74898 169408 75134
rect 169088 74866 169408 74898
rect 199808 75454 200128 75486
rect 199808 75218 199850 75454
rect 200086 75218 200128 75454
rect 199808 75134 200128 75218
rect 199808 74898 199850 75134
rect 200086 74898 200128 75134
rect 199808 74866 200128 74898
rect 230528 75454 230848 75486
rect 230528 75218 230570 75454
rect 230806 75218 230848 75454
rect 230528 75134 230848 75218
rect 230528 74898 230570 75134
rect 230806 74898 230848 75134
rect 230528 74866 230848 74898
rect 261248 75454 261568 75486
rect 261248 75218 261290 75454
rect 261526 75218 261568 75454
rect 261248 75134 261568 75218
rect 261248 74898 261290 75134
rect 261526 74898 261568 75134
rect 261248 74866 261568 74898
rect 291968 75454 292288 75486
rect 291968 75218 292010 75454
rect 292246 75218 292288 75454
rect 291968 75134 292288 75218
rect 291968 74898 292010 75134
rect 292246 74898 292288 75134
rect 291968 74866 292288 74898
rect 322688 75454 323008 75486
rect 322688 75218 322730 75454
rect 322966 75218 323008 75454
rect 322688 75134 323008 75218
rect 322688 74898 322730 75134
rect 322966 74898 323008 75134
rect 322688 74866 323008 74898
rect 353408 75454 353728 75486
rect 353408 75218 353450 75454
rect 353686 75218 353728 75454
rect 353408 75134 353728 75218
rect 353408 74898 353450 75134
rect 353686 74898 353728 75134
rect 353408 74866 353728 74898
rect 384128 75454 384448 75486
rect 384128 75218 384170 75454
rect 384406 75218 384448 75454
rect 384128 75134 384448 75218
rect 384128 74898 384170 75134
rect 384406 74898 384448 75134
rect 384128 74866 384448 74898
rect 414848 75454 415168 75486
rect 414848 75218 414890 75454
rect 415126 75218 415168 75454
rect 414848 75134 415168 75218
rect 414848 74898 414890 75134
rect 415126 74898 415168 75134
rect 414848 74866 415168 74898
rect 445568 75454 445888 75486
rect 445568 75218 445610 75454
rect 445846 75218 445888 75454
rect 445568 75134 445888 75218
rect 445568 74898 445610 75134
rect 445846 74898 445888 75134
rect 445568 74866 445888 74898
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 61568 57454 61888 57486
rect 61568 57218 61610 57454
rect 61846 57218 61888 57454
rect 61568 57134 61888 57218
rect 61568 56898 61610 57134
rect 61846 56898 61888 57134
rect 61568 56866 61888 56898
rect 92288 57454 92608 57486
rect 92288 57218 92330 57454
rect 92566 57218 92608 57454
rect 92288 57134 92608 57218
rect 92288 56898 92330 57134
rect 92566 56898 92608 57134
rect 92288 56866 92608 56898
rect 123008 57454 123328 57486
rect 123008 57218 123050 57454
rect 123286 57218 123328 57454
rect 123008 57134 123328 57218
rect 123008 56898 123050 57134
rect 123286 56898 123328 57134
rect 123008 56866 123328 56898
rect 153728 57454 154048 57486
rect 153728 57218 153770 57454
rect 154006 57218 154048 57454
rect 153728 57134 154048 57218
rect 153728 56898 153770 57134
rect 154006 56898 154048 57134
rect 153728 56866 154048 56898
rect 184448 57454 184768 57486
rect 184448 57218 184490 57454
rect 184726 57218 184768 57454
rect 184448 57134 184768 57218
rect 184448 56898 184490 57134
rect 184726 56898 184768 57134
rect 184448 56866 184768 56898
rect 215168 57454 215488 57486
rect 215168 57218 215210 57454
rect 215446 57218 215488 57454
rect 215168 57134 215488 57218
rect 215168 56898 215210 57134
rect 215446 56898 215488 57134
rect 215168 56866 215488 56898
rect 245888 57454 246208 57486
rect 245888 57218 245930 57454
rect 246166 57218 246208 57454
rect 245888 57134 246208 57218
rect 245888 56898 245930 57134
rect 246166 56898 246208 57134
rect 245888 56866 246208 56898
rect 276608 57454 276928 57486
rect 276608 57218 276650 57454
rect 276886 57218 276928 57454
rect 276608 57134 276928 57218
rect 276608 56898 276650 57134
rect 276886 56898 276928 57134
rect 276608 56866 276928 56898
rect 307328 57454 307648 57486
rect 307328 57218 307370 57454
rect 307606 57218 307648 57454
rect 307328 57134 307648 57218
rect 307328 56898 307370 57134
rect 307606 56898 307648 57134
rect 307328 56866 307648 56898
rect 338048 57454 338368 57486
rect 338048 57218 338090 57454
rect 338326 57218 338368 57454
rect 338048 57134 338368 57218
rect 338048 56898 338090 57134
rect 338326 56898 338368 57134
rect 338048 56866 338368 56898
rect 368768 57454 369088 57486
rect 368768 57218 368810 57454
rect 369046 57218 369088 57454
rect 368768 57134 369088 57218
rect 368768 56898 368810 57134
rect 369046 56898 369088 57134
rect 368768 56866 369088 56898
rect 399488 57454 399808 57486
rect 399488 57218 399530 57454
rect 399766 57218 399808 57454
rect 399488 57134 399808 57218
rect 399488 56898 399530 57134
rect 399766 56898 399808 57134
rect 399488 56866 399808 56898
rect 430208 57454 430528 57486
rect 430208 57218 430250 57454
rect 430486 57218 430528 57454
rect 430208 57134 430528 57218
rect 430208 56898 430250 57134
rect 430486 56898 430528 57134
rect 430208 56866 430528 56898
rect 460928 57454 461248 57486
rect 460928 57218 460970 57454
rect 461206 57218 461248 57454
rect 460928 57134 461248 57218
rect 460928 56898 460970 57134
rect 461206 56898 461248 57134
rect 460928 56866 461248 56898
rect 55794 21454 56414 40000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 52315 19412 52381 19413
rect 52315 19348 52316 19412
rect 52380 19348 52381 19412
rect 52315 19347 52381 19348
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 40000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 40000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 40000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 40000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 40000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 40000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 40000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 40000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 40000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 40000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 40000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 40000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 40000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 40000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 40000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 40000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 40000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 40000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 40000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 40000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 7174 150134 40000
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 40000
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 40000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 40000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 40000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 40000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 40000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 40000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 40000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 40000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 40000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 40000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 40000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 40000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 40000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 40000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 40000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 40000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 40000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 40000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 40000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 40000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 40000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 40000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 40000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 40000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 40000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 40000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 40000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 40000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 40000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 40000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 40000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 40000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 40000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 40000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 40000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 40000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 40000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 40000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 40000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 40000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 40000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 40000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 40000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 40000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 40000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 40000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 40000
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 40000
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 40000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 40000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 40000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 40000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 40000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 40000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 40000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 40000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 40000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 40000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 40000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 40000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 40000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 40000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 40000
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 40000
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 40000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 40000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 40000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 40000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 40000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 46250 435218 46486 435454
rect 46250 434898 46486 435134
rect 46250 399218 46486 399454
rect 46250 398898 46486 399134
rect 46250 363218 46486 363454
rect 46250 362898 46486 363134
rect 46250 327218 46486 327454
rect 46250 326898 46486 327134
rect 46250 291218 46486 291454
rect 46250 290898 46486 291134
rect 46250 255218 46486 255454
rect 46250 254898 46486 255134
rect 46250 219218 46486 219454
rect 46250 218898 46486 219134
rect 46250 183218 46486 183454
rect 46250 182898 46486 183134
rect 46250 147218 46486 147454
rect 46250 146898 46486 147134
rect 46250 111218 46486 111454
rect 46250 110898 46486 111134
rect 46250 75218 46486 75454
rect 46250 74898 46486 75134
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 61610 453218 61846 453454
rect 61610 452898 61846 453134
rect 92330 453218 92566 453454
rect 92330 452898 92566 453134
rect 123050 453218 123286 453454
rect 123050 452898 123286 453134
rect 153770 453218 154006 453454
rect 153770 452898 154006 453134
rect 184490 453218 184726 453454
rect 184490 452898 184726 453134
rect 215210 453218 215446 453454
rect 215210 452898 215446 453134
rect 245930 453218 246166 453454
rect 245930 452898 246166 453134
rect 276650 453218 276886 453454
rect 276650 452898 276886 453134
rect 307370 453218 307606 453454
rect 307370 452898 307606 453134
rect 338090 453218 338326 453454
rect 338090 452898 338326 453134
rect 368810 453218 369046 453454
rect 368810 452898 369046 453134
rect 399530 453218 399766 453454
rect 399530 452898 399766 453134
rect 430250 453218 430486 453454
rect 430250 452898 430486 453134
rect 460970 453218 461206 453454
rect 460970 452898 461206 453134
rect 76970 435218 77206 435454
rect 76970 434898 77206 435134
rect 107690 435218 107926 435454
rect 107690 434898 107926 435134
rect 138410 435218 138646 435454
rect 138410 434898 138646 435134
rect 169130 435218 169366 435454
rect 169130 434898 169366 435134
rect 199850 435218 200086 435454
rect 199850 434898 200086 435134
rect 230570 435218 230806 435454
rect 230570 434898 230806 435134
rect 261290 435218 261526 435454
rect 261290 434898 261526 435134
rect 292010 435218 292246 435454
rect 292010 434898 292246 435134
rect 322730 435218 322966 435454
rect 322730 434898 322966 435134
rect 353450 435218 353686 435454
rect 353450 434898 353686 435134
rect 384170 435218 384406 435454
rect 384170 434898 384406 435134
rect 414890 435218 415126 435454
rect 414890 434898 415126 435134
rect 445610 435218 445846 435454
rect 445610 434898 445846 435134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 61610 417218 61846 417454
rect 61610 416898 61846 417134
rect 92330 417218 92566 417454
rect 92330 416898 92566 417134
rect 123050 417218 123286 417454
rect 123050 416898 123286 417134
rect 153770 417218 154006 417454
rect 153770 416898 154006 417134
rect 184490 417218 184726 417454
rect 184490 416898 184726 417134
rect 215210 417218 215446 417454
rect 215210 416898 215446 417134
rect 245930 417218 246166 417454
rect 245930 416898 246166 417134
rect 276650 417218 276886 417454
rect 276650 416898 276886 417134
rect 307370 417218 307606 417454
rect 307370 416898 307606 417134
rect 338090 417218 338326 417454
rect 338090 416898 338326 417134
rect 368810 417218 369046 417454
rect 368810 416898 369046 417134
rect 399530 417218 399766 417454
rect 399530 416898 399766 417134
rect 430250 417218 430486 417454
rect 430250 416898 430486 417134
rect 460970 417218 461206 417454
rect 460970 416898 461206 417134
rect 76970 399218 77206 399454
rect 76970 398898 77206 399134
rect 107690 399218 107926 399454
rect 107690 398898 107926 399134
rect 138410 399218 138646 399454
rect 138410 398898 138646 399134
rect 169130 399218 169366 399454
rect 169130 398898 169366 399134
rect 199850 399218 200086 399454
rect 199850 398898 200086 399134
rect 230570 399218 230806 399454
rect 230570 398898 230806 399134
rect 261290 399218 261526 399454
rect 261290 398898 261526 399134
rect 292010 399218 292246 399454
rect 292010 398898 292246 399134
rect 322730 399218 322966 399454
rect 322730 398898 322966 399134
rect 353450 399218 353686 399454
rect 353450 398898 353686 399134
rect 384170 399218 384406 399454
rect 384170 398898 384406 399134
rect 414890 399218 415126 399454
rect 414890 398898 415126 399134
rect 445610 399218 445846 399454
rect 445610 398898 445846 399134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 61610 381218 61846 381454
rect 61610 380898 61846 381134
rect 92330 381218 92566 381454
rect 92330 380898 92566 381134
rect 123050 381218 123286 381454
rect 123050 380898 123286 381134
rect 153770 381218 154006 381454
rect 153770 380898 154006 381134
rect 184490 381218 184726 381454
rect 184490 380898 184726 381134
rect 215210 381218 215446 381454
rect 215210 380898 215446 381134
rect 245930 381218 246166 381454
rect 245930 380898 246166 381134
rect 276650 381218 276886 381454
rect 276650 380898 276886 381134
rect 307370 381218 307606 381454
rect 307370 380898 307606 381134
rect 338090 381218 338326 381454
rect 338090 380898 338326 381134
rect 368810 381218 369046 381454
rect 368810 380898 369046 381134
rect 399530 381218 399766 381454
rect 399530 380898 399766 381134
rect 430250 381218 430486 381454
rect 430250 380898 430486 381134
rect 460970 381218 461206 381454
rect 460970 380898 461206 381134
rect 76970 363218 77206 363454
rect 76970 362898 77206 363134
rect 107690 363218 107926 363454
rect 107690 362898 107926 363134
rect 138410 363218 138646 363454
rect 138410 362898 138646 363134
rect 169130 363218 169366 363454
rect 169130 362898 169366 363134
rect 199850 363218 200086 363454
rect 199850 362898 200086 363134
rect 230570 363218 230806 363454
rect 230570 362898 230806 363134
rect 261290 363218 261526 363454
rect 261290 362898 261526 363134
rect 292010 363218 292246 363454
rect 292010 362898 292246 363134
rect 322730 363218 322966 363454
rect 322730 362898 322966 363134
rect 353450 363218 353686 363454
rect 353450 362898 353686 363134
rect 384170 363218 384406 363454
rect 384170 362898 384406 363134
rect 414890 363218 415126 363454
rect 414890 362898 415126 363134
rect 445610 363218 445846 363454
rect 445610 362898 445846 363134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 61610 345218 61846 345454
rect 61610 344898 61846 345134
rect 92330 345218 92566 345454
rect 92330 344898 92566 345134
rect 123050 345218 123286 345454
rect 123050 344898 123286 345134
rect 153770 345218 154006 345454
rect 153770 344898 154006 345134
rect 184490 345218 184726 345454
rect 184490 344898 184726 345134
rect 215210 345218 215446 345454
rect 215210 344898 215446 345134
rect 245930 345218 246166 345454
rect 245930 344898 246166 345134
rect 276650 345218 276886 345454
rect 276650 344898 276886 345134
rect 307370 345218 307606 345454
rect 307370 344898 307606 345134
rect 338090 345218 338326 345454
rect 338090 344898 338326 345134
rect 368810 345218 369046 345454
rect 368810 344898 369046 345134
rect 399530 345218 399766 345454
rect 399530 344898 399766 345134
rect 430250 345218 430486 345454
rect 430250 344898 430486 345134
rect 460970 345218 461206 345454
rect 460970 344898 461206 345134
rect 76970 327218 77206 327454
rect 76970 326898 77206 327134
rect 107690 327218 107926 327454
rect 107690 326898 107926 327134
rect 138410 327218 138646 327454
rect 138410 326898 138646 327134
rect 169130 327218 169366 327454
rect 169130 326898 169366 327134
rect 199850 327218 200086 327454
rect 199850 326898 200086 327134
rect 230570 327218 230806 327454
rect 230570 326898 230806 327134
rect 261290 327218 261526 327454
rect 261290 326898 261526 327134
rect 292010 327218 292246 327454
rect 292010 326898 292246 327134
rect 322730 327218 322966 327454
rect 322730 326898 322966 327134
rect 353450 327218 353686 327454
rect 353450 326898 353686 327134
rect 384170 327218 384406 327454
rect 384170 326898 384406 327134
rect 414890 327218 415126 327454
rect 414890 326898 415126 327134
rect 445610 327218 445846 327454
rect 445610 326898 445846 327134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 61610 309218 61846 309454
rect 61610 308898 61846 309134
rect 92330 309218 92566 309454
rect 92330 308898 92566 309134
rect 123050 309218 123286 309454
rect 123050 308898 123286 309134
rect 153770 309218 154006 309454
rect 153770 308898 154006 309134
rect 184490 309218 184726 309454
rect 184490 308898 184726 309134
rect 215210 309218 215446 309454
rect 215210 308898 215446 309134
rect 245930 309218 246166 309454
rect 245930 308898 246166 309134
rect 276650 309218 276886 309454
rect 276650 308898 276886 309134
rect 307370 309218 307606 309454
rect 307370 308898 307606 309134
rect 338090 309218 338326 309454
rect 338090 308898 338326 309134
rect 368810 309218 369046 309454
rect 368810 308898 369046 309134
rect 399530 309218 399766 309454
rect 399530 308898 399766 309134
rect 430250 309218 430486 309454
rect 430250 308898 430486 309134
rect 460970 309218 461206 309454
rect 460970 308898 461206 309134
rect 76970 291218 77206 291454
rect 76970 290898 77206 291134
rect 107690 291218 107926 291454
rect 107690 290898 107926 291134
rect 138410 291218 138646 291454
rect 138410 290898 138646 291134
rect 169130 291218 169366 291454
rect 169130 290898 169366 291134
rect 199850 291218 200086 291454
rect 199850 290898 200086 291134
rect 230570 291218 230806 291454
rect 230570 290898 230806 291134
rect 261290 291218 261526 291454
rect 261290 290898 261526 291134
rect 292010 291218 292246 291454
rect 292010 290898 292246 291134
rect 322730 291218 322966 291454
rect 322730 290898 322966 291134
rect 353450 291218 353686 291454
rect 353450 290898 353686 291134
rect 384170 291218 384406 291454
rect 384170 290898 384406 291134
rect 414890 291218 415126 291454
rect 414890 290898 415126 291134
rect 445610 291218 445846 291454
rect 445610 290898 445846 291134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 61610 273218 61846 273454
rect 61610 272898 61846 273134
rect 92330 273218 92566 273454
rect 92330 272898 92566 273134
rect 123050 273218 123286 273454
rect 123050 272898 123286 273134
rect 153770 273218 154006 273454
rect 153770 272898 154006 273134
rect 184490 273218 184726 273454
rect 184490 272898 184726 273134
rect 215210 273218 215446 273454
rect 215210 272898 215446 273134
rect 245930 273218 246166 273454
rect 245930 272898 246166 273134
rect 276650 273218 276886 273454
rect 276650 272898 276886 273134
rect 307370 273218 307606 273454
rect 307370 272898 307606 273134
rect 338090 273218 338326 273454
rect 338090 272898 338326 273134
rect 368810 273218 369046 273454
rect 368810 272898 369046 273134
rect 399530 273218 399766 273454
rect 399530 272898 399766 273134
rect 430250 273218 430486 273454
rect 430250 272898 430486 273134
rect 460970 273218 461206 273454
rect 460970 272898 461206 273134
rect 76970 255218 77206 255454
rect 76970 254898 77206 255134
rect 107690 255218 107926 255454
rect 107690 254898 107926 255134
rect 138410 255218 138646 255454
rect 138410 254898 138646 255134
rect 169130 255218 169366 255454
rect 169130 254898 169366 255134
rect 199850 255218 200086 255454
rect 199850 254898 200086 255134
rect 230570 255218 230806 255454
rect 230570 254898 230806 255134
rect 261290 255218 261526 255454
rect 261290 254898 261526 255134
rect 292010 255218 292246 255454
rect 292010 254898 292246 255134
rect 322730 255218 322966 255454
rect 322730 254898 322966 255134
rect 353450 255218 353686 255454
rect 353450 254898 353686 255134
rect 384170 255218 384406 255454
rect 384170 254898 384406 255134
rect 414890 255218 415126 255454
rect 414890 254898 415126 255134
rect 445610 255218 445846 255454
rect 445610 254898 445846 255134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 61610 237218 61846 237454
rect 61610 236898 61846 237134
rect 92330 237218 92566 237454
rect 92330 236898 92566 237134
rect 123050 237218 123286 237454
rect 123050 236898 123286 237134
rect 153770 237218 154006 237454
rect 153770 236898 154006 237134
rect 184490 237218 184726 237454
rect 184490 236898 184726 237134
rect 215210 237218 215446 237454
rect 215210 236898 215446 237134
rect 245930 237218 246166 237454
rect 245930 236898 246166 237134
rect 276650 237218 276886 237454
rect 276650 236898 276886 237134
rect 307370 237218 307606 237454
rect 307370 236898 307606 237134
rect 338090 237218 338326 237454
rect 338090 236898 338326 237134
rect 368810 237218 369046 237454
rect 368810 236898 369046 237134
rect 399530 237218 399766 237454
rect 399530 236898 399766 237134
rect 430250 237218 430486 237454
rect 430250 236898 430486 237134
rect 460970 237218 461206 237454
rect 460970 236898 461206 237134
rect 76970 219218 77206 219454
rect 76970 218898 77206 219134
rect 107690 219218 107926 219454
rect 107690 218898 107926 219134
rect 138410 219218 138646 219454
rect 138410 218898 138646 219134
rect 169130 219218 169366 219454
rect 169130 218898 169366 219134
rect 199850 219218 200086 219454
rect 199850 218898 200086 219134
rect 230570 219218 230806 219454
rect 230570 218898 230806 219134
rect 261290 219218 261526 219454
rect 261290 218898 261526 219134
rect 292010 219218 292246 219454
rect 292010 218898 292246 219134
rect 322730 219218 322966 219454
rect 322730 218898 322966 219134
rect 353450 219218 353686 219454
rect 353450 218898 353686 219134
rect 384170 219218 384406 219454
rect 384170 218898 384406 219134
rect 414890 219218 415126 219454
rect 414890 218898 415126 219134
rect 445610 219218 445846 219454
rect 445610 218898 445846 219134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 61610 201218 61846 201454
rect 61610 200898 61846 201134
rect 92330 201218 92566 201454
rect 92330 200898 92566 201134
rect 123050 201218 123286 201454
rect 123050 200898 123286 201134
rect 153770 201218 154006 201454
rect 153770 200898 154006 201134
rect 184490 201218 184726 201454
rect 184490 200898 184726 201134
rect 215210 201218 215446 201454
rect 215210 200898 215446 201134
rect 245930 201218 246166 201454
rect 245930 200898 246166 201134
rect 276650 201218 276886 201454
rect 276650 200898 276886 201134
rect 307370 201218 307606 201454
rect 307370 200898 307606 201134
rect 338090 201218 338326 201454
rect 338090 200898 338326 201134
rect 368810 201218 369046 201454
rect 368810 200898 369046 201134
rect 399530 201218 399766 201454
rect 399530 200898 399766 201134
rect 430250 201218 430486 201454
rect 430250 200898 430486 201134
rect 460970 201218 461206 201454
rect 460970 200898 461206 201134
rect 76970 183218 77206 183454
rect 76970 182898 77206 183134
rect 107690 183218 107926 183454
rect 107690 182898 107926 183134
rect 138410 183218 138646 183454
rect 138410 182898 138646 183134
rect 169130 183218 169366 183454
rect 169130 182898 169366 183134
rect 199850 183218 200086 183454
rect 199850 182898 200086 183134
rect 230570 183218 230806 183454
rect 230570 182898 230806 183134
rect 261290 183218 261526 183454
rect 261290 182898 261526 183134
rect 292010 183218 292246 183454
rect 292010 182898 292246 183134
rect 322730 183218 322966 183454
rect 322730 182898 322966 183134
rect 353450 183218 353686 183454
rect 353450 182898 353686 183134
rect 384170 183218 384406 183454
rect 384170 182898 384406 183134
rect 414890 183218 415126 183454
rect 414890 182898 415126 183134
rect 445610 183218 445846 183454
rect 445610 182898 445846 183134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 61610 165218 61846 165454
rect 61610 164898 61846 165134
rect 92330 165218 92566 165454
rect 92330 164898 92566 165134
rect 123050 165218 123286 165454
rect 123050 164898 123286 165134
rect 153770 165218 154006 165454
rect 153770 164898 154006 165134
rect 184490 165218 184726 165454
rect 184490 164898 184726 165134
rect 215210 165218 215446 165454
rect 215210 164898 215446 165134
rect 245930 165218 246166 165454
rect 245930 164898 246166 165134
rect 276650 165218 276886 165454
rect 276650 164898 276886 165134
rect 307370 165218 307606 165454
rect 307370 164898 307606 165134
rect 338090 165218 338326 165454
rect 338090 164898 338326 165134
rect 368810 165218 369046 165454
rect 368810 164898 369046 165134
rect 399530 165218 399766 165454
rect 399530 164898 399766 165134
rect 430250 165218 430486 165454
rect 430250 164898 430486 165134
rect 460970 165218 461206 165454
rect 460970 164898 461206 165134
rect 76970 147218 77206 147454
rect 76970 146898 77206 147134
rect 107690 147218 107926 147454
rect 107690 146898 107926 147134
rect 138410 147218 138646 147454
rect 138410 146898 138646 147134
rect 169130 147218 169366 147454
rect 169130 146898 169366 147134
rect 199850 147218 200086 147454
rect 199850 146898 200086 147134
rect 230570 147218 230806 147454
rect 230570 146898 230806 147134
rect 261290 147218 261526 147454
rect 261290 146898 261526 147134
rect 292010 147218 292246 147454
rect 292010 146898 292246 147134
rect 322730 147218 322966 147454
rect 322730 146898 322966 147134
rect 353450 147218 353686 147454
rect 353450 146898 353686 147134
rect 384170 147218 384406 147454
rect 384170 146898 384406 147134
rect 414890 147218 415126 147454
rect 414890 146898 415126 147134
rect 445610 147218 445846 147454
rect 445610 146898 445846 147134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 61610 129218 61846 129454
rect 61610 128898 61846 129134
rect 92330 129218 92566 129454
rect 92330 128898 92566 129134
rect 123050 129218 123286 129454
rect 123050 128898 123286 129134
rect 153770 129218 154006 129454
rect 153770 128898 154006 129134
rect 184490 129218 184726 129454
rect 184490 128898 184726 129134
rect 215210 129218 215446 129454
rect 215210 128898 215446 129134
rect 245930 129218 246166 129454
rect 245930 128898 246166 129134
rect 276650 129218 276886 129454
rect 276650 128898 276886 129134
rect 307370 129218 307606 129454
rect 307370 128898 307606 129134
rect 338090 129218 338326 129454
rect 338090 128898 338326 129134
rect 368810 129218 369046 129454
rect 368810 128898 369046 129134
rect 399530 129218 399766 129454
rect 399530 128898 399766 129134
rect 430250 129218 430486 129454
rect 430250 128898 430486 129134
rect 460970 129218 461206 129454
rect 460970 128898 461206 129134
rect 76970 111218 77206 111454
rect 76970 110898 77206 111134
rect 107690 111218 107926 111454
rect 107690 110898 107926 111134
rect 138410 111218 138646 111454
rect 138410 110898 138646 111134
rect 169130 111218 169366 111454
rect 169130 110898 169366 111134
rect 199850 111218 200086 111454
rect 199850 110898 200086 111134
rect 230570 111218 230806 111454
rect 230570 110898 230806 111134
rect 261290 111218 261526 111454
rect 261290 110898 261526 111134
rect 292010 111218 292246 111454
rect 292010 110898 292246 111134
rect 322730 111218 322966 111454
rect 322730 110898 322966 111134
rect 353450 111218 353686 111454
rect 353450 110898 353686 111134
rect 384170 111218 384406 111454
rect 384170 110898 384406 111134
rect 414890 111218 415126 111454
rect 414890 110898 415126 111134
rect 445610 111218 445846 111454
rect 445610 110898 445846 111134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 61610 93218 61846 93454
rect 61610 92898 61846 93134
rect 92330 93218 92566 93454
rect 92330 92898 92566 93134
rect 123050 93218 123286 93454
rect 123050 92898 123286 93134
rect 153770 93218 154006 93454
rect 153770 92898 154006 93134
rect 184490 93218 184726 93454
rect 184490 92898 184726 93134
rect 215210 93218 215446 93454
rect 215210 92898 215446 93134
rect 245930 93218 246166 93454
rect 245930 92898 246166 93134
rect 276650 93218 276886 93454
rect 276650 92898 276886 93134
rect 307370 93218 307606 93454
rect 307370 92898 307606 93134
rect 338090 93218 338326 93454
rect 338090 92898 338326 93134
rect 368810 93218 369046 93454
rect 368810 92898 369046 93134
rect 399530 93218 399766 93454
rect 399530 92898 399766 93134
rect 430250 93218 430486 93454
rect 430250 92898 430486 93134
rect 460970 93218 461206 93454
rect 460970 92898 461206 93134
rect 76970 75218 77206 75454
rect 76970 74898 77206 75134
rect 107690 75218 107926 75454
rect 107690 74898 107926 75134
rect 138410 75218 138646 75454
rect 138410 74898 138646 75134
rect 169130 75218 169366 75454
rect 169130 74898 169366 75134
rect 199850 75218 200086 75454
rect 199850 74898 200086 75134
rect 230570 75218 230806 75454
rect 230570 74898 230806 75134
rect 261290 75218 261526 75454
rect 261290 74898 261526 75134
rect 292010 75218 292246 75454
rect 292010 74898 292246 75134
rect 322730 75218 322966 75454
rect 322730 74898 322966 75134
rect 353450 75218 353686 75454
rect 353450 74898 353686 75134
rect 384170 75218 384406 75454
rect 384170 74898 384406 75134
rect 414890 75218 415126 75454
rect 414890 74898 415126 75134
rect 445610 75218 445846 75454
rect 445610 74898 445846 75134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 61610 57218 61846 57454
rect 61610 56898 61846 57134
rect 92330 57218 92566 57454
rect 92330 56898 92566 57134
rect 123050 57218 123286 57454
rect 123050 56898 123286 57134
rect 153770 57218 154006 57454
rect 153770 56898 154006 57134
rect 184490 57218 184726 57454
rect 184490 56898 184726 57134
rect 215210 57218 215446 57454
rect 215210 56898 215446 57134
rect 245930 57218 246166 57454
rect 245930 56898 246166 57134
rect 276650 57218 276886 57454
rect 276650 56898 276886 57134
rect 307370 57218 307606 57454
rect 307370 56898 307606 57134
rect 338090 57218 338326 57454
rect 338090 56898 338326 57134
rect 368810 57218 369046 57454
rect 368810 56898 369046 57134
rect 399530 57218 399766 57454
rect 399530 56898 399766 57134
rect 430250 57218 430486 57454
rect 430250 56898 430486 57134
rect 460970 57218 461206 57454
rect 460970 56898 461206 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 61610 453454
rect 61846 453218 92330 453454
rect 92566 453218 123050 453454
rect 123286 453218 153770 453454
rect 154006 453218 184490 453454
rect 184726 453218 215210 453454
rect 215446 453218 245930 453454
rect 246166 453218 276650 453454
rect 276886 453218 307370 453454
rect 307606 453218 338090 453454
rect 338326 453218 368810 453454
rect 369046 453218 399530 453454
rect 399766 453218 430250 453454
rect 430486 453218 460970 453454
rect 461206 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 61610 453134
rect 61846 452898 92330 453134
rect 92566 452898 123050 453134
rect 123286 452898 153770 453134
rect 154006 452898 184490 453134
rect 184726 452898 215210 453134
rect 215446 452898 245930 453134
rect 246166 452898 276650 453134
rect 276886 452898 307370 453134
rect 307606 452898 338090 453134
rect 338326 452898 368810 453134
rect 369046 452898 399530 453134
rect 399766 452898 430250 453134
rect 430486 452898 460970 453134
rect 461206 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 46250 435454
rect 46486 435218 76970 435454
rect 77206 435218 107690 435454
rect 107926 435218 138410 435454
rect 138646 435218 169130 435454
rect 169366 435218 199850 435454
rect 200086 435218 230570 435454
rect 230806 435218 261290 435454
rect 261526 435218 292010 435454
rect 292246 435218 322730 435454
rect 322966 435218 353450 435454
rect 353686 435218 384170 435454
rect 384406 435218 414890 435454
rect 415126 435218 445610 435454
rect 445846 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 46250 435134
rect 46486 434898 76970 435134
rect 77206 434898 107690 435134
rect 107926 434898 138410 435134
rect 138646 434898 169130 435134
rect 169366 434898 199850 435134
rect 200086 434898 230570 435134
rect 230806 434898 261290 435134
rect 261526 434898 292010 435134
rect 292246 434898 322730 435134
rect 322966 434898 353450 435134
rect 353686 434898 384170 435134
rect 384406 434898 414890 435134
rect 415126 434898 445610 435134
rect 445846 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 61610 417454
rect 61846 417218 92330 417454
rect 92566 417218 123050 417454
rect 123286 417218 153770 417454
rect 154006 417218 184490 417454
rect 184726 417218 215210 417454
rect 215446 417218 245930 417454
rect 246166 417218 276650 417454
rect 276886 417218 307370 417454
rect 307606 417218 338090 417454
rect 338326 417218 368810 417454
rect 369046 417218 399530 417454
rect 399766 417218 430250 417454
rect 430486 417218 460970 417454
rect 461206 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 61610 417134
rect 61846 416898 92330 417134
rect 92566 416898 123050 417134
rect 123286 416898 153770 417134
rect 154006 416898 184490 417134
rect 184726 416898 215210 417134
rect 215446 416898 245930 417134
rect 246166 416898 276650 417134
rect 276886 416898 307370 417134
rect 307606 416898 338090 417134
rect 338326 416898 368810 417134
rect 369046 416898 399530 417134
rect 399766 416898 430250 417134
rect 430486 416898 460970 417134
rect 461206 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 46250 399454
rect 46486 399218 76970 399454
rect 77206 399218 107690 399454
rect 107926 399218 138410 399454
rect 138646 399218 169130 399454
rect 169366 399218 199850 399454
rect 200086 399218 230570 399454
rect 230806 399218 261290 399454
rect 261526 399218 292010 399454
rect 292246 399218 322730 399454
rect 322966 399218 353450 399454
rect 353686 399218 384170 399454
rect 384406 399218 414890 399454
rect 415126 399218 445610 399454
rect 445846 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 46250 399134
rect 46486 398898 76970 399134
rect 77206 398898 107690 399134
rect 107926 398898 138410 399134
rect 138646 398898 169130 399134
rect 169366 398898 199850 399134
rect 200086 398898 230570 399134
rect 230806 398898 261290 399134
rect 261526 398898 292010 399134
rect 292246 398898 322730 399134
rect 322966 398898 353450 399134
rect 353686 398898 384170 399134
rect 384406 398898 414890 399134
rect 415126 398898 445610 399134
rect 445846 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 61610 381454
rect 61846 381218 92330 381454
rect 92566 381218 123050 381454
rect 123286 381218 153770 381454
rect 154006 381218 184490 381454
rect 184726 381218 215210 381454
rect 215446 381218 245930 381454
rect 246166 381218 276650 381454
rect 276886 381218 307370 381454
rect 307606 381218 338090 381454
rect 338326 381218 368810 381454
rect 369046 381218 399530 381454
rect 399766 381218 430250 381454
rect 430486 381218 460970 381454
rect 461206 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 61610 381134
rect 61846 380898 92330 381134
rect 92566 380898 123050 381134
rect 123286 380898 153770 381134
rect 154006 380898 184490 381134
rect 184726 380898 215210 381134
rect 215446 380898 245930 381134
rect 246166 380898 276650 381134
rect 276886 380898 307370 381134
rect 307606 380898 338090 381134
rect 338326 380898 368810 381134
rect 369046 380898 399530 381134
rect 399766 380898 430250 381134
rect 430486 380898 460970 381134
rect 461206 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 46250 363454
rect 46486 363218 76970 363454
rect 77206 363218 107690 363454
rect 107926 363218 138410 363454
rect 138646 363218 169130 363454
rect 169366 363218 199850 363454
rect 200086 363218 230570 363454
rect 230806 363218 261290 363454
rect 261526 363218 292010 363454
rect 292246 363218 322730 363454
rect 322966 363218 353450 363454
rect 353686 363218 384170 363454
rect 384406 363218 414890 363454
rect 415126 363218 445610 363454
rect 445846 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 46250 363134
rect 46486 362898 76970 363134
rect 77206 362898 107690 363134
rect 107926 362898 138410 363134
rect 138646 362898 169130 363134
rect 169366 362898 199850 363134
rect 200086 362898 230570 363134
rect 230806 362898 261290 363134
rect 261526 362898 292010 363134
rect 292246 362898 322730 363134
rect 322966 362898 353450 363134
rect 353686 362898 384170 363134
rect 384406 362898 414890 363134
rect 415126 362898 445610 363134
rect 445846 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 61610 345454
rect 61846 345218 92330 345454
rect 92566 345218 123050 345454
rect 123286 345218 153770 345454
rect 154006 345218 184490 345454
rect 184726 345218 215210 345454
rect 215446 345218 245930 345454
rect 246166 345218 276650 345454
rect 276886 345218 307370 345454
rect 307606 345218 338090 345454
rect 338326 345218 368810 345454
rect 369046 345218 399530 345454
rect 399766 345218 430250 345454
rect 430486 345218 460970 345454
rect 461206 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 61610 345134
rect 61846 344898 92330 345134
rect 92566 344898 123050 345134
rect 123286 344898 153770 345134
rect 154006 344898 184490 345134
rect 184726 344898 215210 345134
rect 215446 344898 245930 345134
rect 246166 344898 276650 345134
rect 276886 344898 307370 345134
rect 307606 344898 338090 345134
rect 338326 344898 368810 345134
rect 369046 344898 399530 345134
rect 399766 344898 430250 345134
rect 430486 344898 460970 345134
rect 461206 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 46250 327454
rect 46486 327218 76970 327454
rect 77206 327218 107690 327454
rect 107926 327218 138410 327454
rect 138646 327218 169130 327454
rect 169366 327218 199850 327454
rect 200086 327218 230570 327454
rect 230806 327218 261290 327454
rect 261526 327218 292010 327454
rect 292246 327218 322730 327454
rect 322966 327218 353450 327454
rect 353686 327218 384170 327454
rect 384406 327218 414890 327454
rect 415126 327218 445610 327454
rect 445846 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 46250 327134
rect 46486 326898 76970 327134
rect 77206 326898 107690 327134
rect 107926 326898 138410 327134
rect 138646 326898 169130 327134
rect 169366 326898 199850 327134
rect 200086 326898 230570 327134
rect 230806 326898 261290 327134
rect 261526 326898 292010 327134
rect 292246 326898 322730 327134
rect 322966 326898 353450 327134
rect 353686 326898 384170 327134
rect 384406 326898 414890 327134
rect 415126 326898 445610 327134
rect 445846 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 61610 309454
rect 61846 309218 92330 309454
rect 92566 309218 123050 309454
rect 123286 309218 153770 309454
rect 154006 309218 184490 309454
rect 184726 309218 215210 309454
rect 215446 309218 245930 309454
rect 246166 309218 276650 309454
rect 276886 309218 307370 309454
rect 307606 309218 338090 309454
rect 338326 309218 368810 309454
rect 369046 309218 399530 309454
rect 399766 309218 430250 309454
rect 430486 309218 460970 309454
rect 461206 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 61610 309134
rect 61846 308898 92330 309134
rect 92566 308898 123050 309134
rect 123286 308898 153770 309134
rect 154006 308898 184490 309134
rect 184726 308898 215210 309134
rect 215446 308898 245930 309134
rect 246166 308898 276650 309134
rect 276886 308898 307370 309134
rect 307606 308898 338090 309134
rect 338326 308898 368810 309134
rect 369046 308898 399530 309134
rect 399766 308898 430250 309134
rect 430486 308898 460970 309134
rect 461206 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 46250 291454
rect 46486 291218 76970 291454
rect 77206 291218 107690 291454
rect 107926 291218 138410 291454
rect 138646 291218 169130 291454
rect 169366 291218 199850 291454
rect 200086 291218 230570 291454
rect 230806 291218 261290 291454
rect 261526 291218 292010 291454
rect 292246 291218 322730 291454
rect 322966 291218 353450 291454
rect 353686 291218 384170 291454
rect 384406 291218 414890 291454
rect 415126 291218 445610 291454
rect 445846 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 46250 291134
rect 46486 290898 76970 291134
rect 77206 290898 107690 291134
rect 107926 290898 138410 291134
rect 138646 290898 169130 291134
rect 169366 290898 199850 291134
rect 200086 290898 230570 291134
rect 230806 290898 261290 291134
rect 261526 290898 292010 291134
rect 292246 290898 322730 291134
rect 322966 290898 353450 291134
rect 353686 290898 384170 291134
rect 384406 290898 414890 291134
rect 415126 290898 445610 291134
rect 445846 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 61610 273454
rect 61846 273218 92330 273454
rect 92566 273218 123050 273454
rect 123286 273218 153770 273454
rect 154006 273218 184490 273454
rect 184726 273218 215210 273454
rect 215446 273218 245930 273454
rect 246166 273218 276650 273454
rect 276886 273218 307370 273454
rect 307606 273218 338090 273454
rect 338326 273218 368810 273454
rect 369046 273218 399530 273454
rect 399766 273218 430250 273454
rect 430486 273218 460970 273454
rect 461206 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 61610 273134
rect 61846 272898 92330 273134
rect 92566 272898 123050 273134
rect 123286 272898 153770 273134
rect 154006 272898 184490 273134
rect 184726 272898 215210 273134
rect 215446 272898 245930 273134
rect 246166 272898 276650 273134
rect 276886 272898 307370 273134
rect 307606 272898 338090 273134
rect 338326 272898 368810 273134
rect 369046 272898 399530 273134
rect 399766 272898 430250 273134
rect 430486 272898 460970 273134
rect 461206 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 46250 255454
rect 46486 255218 76970 255454
rect 77206 255218 107690 255454
rect 107926 255218 138410 255454
rect 138646 255218 169130 255454
rect 169366 255218 199850 255454
rect 200086 255218 230570 255454
rect 230806 255218 261290 255454
rect 261526 255218 292010 255454
rect 292246 255218 322730 255454
rect 322966 255218 353450 255454
rect 353686 255218 384170 255454
rect 384406 255218 414890 255454
rect 415126 255218 445610 255454
rect 445846 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 46250 255134
rect 46486 254898 76970 255134
rect 77206 254898 107690 255134
rect 107926 254898 138410 255134
rect 138646 254898 169130 255134
rect 169366 254898 199850 255134
rect 200086 254898 230570 255134
rect 230806 254898 261290 255134
rect 261526 254898 292010 255134
rect 292246 254898 322730 255134
rect 322966 254898 353450 255134
rect 353686 254898 384170 255134
rect 384406 254898 414890 255134
rect 415126 254898 445610 255134
rect 445846 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 61610 237454
rect 61846 237218 92330 237454
rect 92566 237218 123050 237454
rect 123286 237218 153770 237454
rect 154006 237218 184490 237454
rect 184726 237218 215210 237454
rect 215446 237218 245930 237454
rect 246166 237218 276650 237454
rect 276886 237218 307370 237454
rect 307606 237218 338090 237454
rect 338326 237218 368810 237454
rect 369046 237218 399530 237454
rect 399766 237218 430250 237454
rect 430486 237218 460970 237454
rect 461206 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 61610 237134
rect 61846 236898 92330 237134
rect 92566 236898 123050 237134
rect 123286 236898 153770 237134
rect 154006 236898 184490 237134
rect 184726 236898 215210 237134
rect 215446 236898 245930 237134
rect 246166 236898 276650 237134
rect 276886 236898 307370 237134
rect 307606 236898 338090 237134
rect 338326 236898 368810 237134
rect 369046 236898 399530 237134
rect 399766 236898 430250 237134
rect 430486 236898 460970 237134
rect 461206 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 46250 219454
rect 46486 219218 76970 219454
rect 77206 219218 107690 219454
rect 107926 219218 138410 219454
rect 138646 219218 169130 219454
rect 169366 219218 199850 219454
rect 200086 219218 230570 219454
rect 230806 219218 261290 219454
rect 261526 219218 292010 219454
rect 292246 219218 322730 219454
rect 322966 219218 353450 219454
rect 353686 219218 384170 219454
rect 384406 219218 414890 219454
rect 415126 219218 445610 219454
rect 445846 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 46250 219134
rect 46486 218898 76970 219134
rect 77206 218898 107690 219134
rect 107926 218898 138410 219134
rect 138646 218898 169130 219134
rect 169366 218898 199850 219134
rect 200086 218898 230570 219134
rect 230806 218898 261290 219134
rect 261526 218898 292010 219134
rect 292246 218898 322730 219134
rect 322966 218898 353450 219134
rect 353686 218898 384170 219134
rect 384406 218898 414890 219134
rect 415126 218898 445610 219134
rect 445846 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 61610 201454
rect 61846 201218 92330 201454
rect 92566 201218 123050 201454
rect 123286 201218 153770 201454
rect 154006 201218 184490 201454
rect 184726 201218 215210 201454
rect 215446 201218 245930 201454
rect 246166 201218 276650 201454
rect 276886 201218 307370 201454
rect 307606 201218 338090 201454
rect 338326 201218 368810 201454
rect 369046 201218 399530 201454
rect 399766 201218 430250 201454
rect 430486 201218 460970 201454
rect 461206 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 61610 201134
rect 61846 200898 92330 201134
rect 92566 200898 123050 201134
rect 123286 200898 153770 201134
rect 154006 200898 184490 201134
rect 184726 200898 215210 201134
rect 215446 200898 245930 201134
rect 246166 200898 276650 201134
rect 276886 200898 307370 201134
rect 307606 200898 338090 201134
rect 338326 200898 368810 201134
rect 369046 200898 399530 201134
rect 399766 200898 430250 201134
rect 430486 200898 460970 201134
rect 461206 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 46250 183454
rect 46486 183218 76970 183454
rect 77206 183218 107690 183454
rect 107926 183218 138410 183454
rect 138646 183218 169130 183454
rect 169366 183218 199850 183454
rect 200086 183218 230570 183454
rect 230806 183218 261290 183454
rect 261526 183218 292010 183454
rect 292246 183218 322730 183454
rect 322966 183218 353450 183454
rect 353686 183218 384170 183454
rect 384406 183218 414890 183454
rect 415126 183218 445610 183454
rect 445846 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 46250 183134
rect 46486 182898 76970 183134
rect 77206 182898 107690 183134
rect 107926 182898 138410 183134
rect 138646 182898 169130 183134
rect 169366 182898 199850 183134
rect 200086 182898 230570 183134
rect 230806 182898 261290 183134
rect 261526 182898 292010 183134
rect 292246 182898 322730 183134
rect 322966 182898 353450 183134
rect 353686 182898 384170 183134
rect 384406 182898 414890 183134
rect 415126 182898 445610 183134
rect 445846 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 61610 165454
rect 61846 165218 92330 165454
rect 92566 165218 123050 165454
rect 123286 165218 153770 165454
rect 154006 165218 184490 165454
rect 184726 165218 215210 165454
rect 215446 165218 245930 165454
rect 246166 165218 276650 165454
rect 276886 165218 307370 165454
rect 307606 165218 338090 165454
rect 338326 165218 368810 165454
rect 369046 165218 399530 165454
rect 399766 165218 430250 165454
rect 430486 165218 460970 165454
rect 461206 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 61610 165134
rect 61846 164898 92330 165134
rect 92566 164898 123050 165134
rect 123286 164898 153770 165134
rect 154006 164898 184490 165134
rect 184726 164898 215210 165134
rect 215446 164898 245930 165134
rect 246166 164898 276650 165134
rect 276886 164898 307370 165134
rect 307606 164898 338090 165134
rect 338326 164898 368810 165134
rect 369046 164898 399530 165134
rect 399766 164898 430250 165134
rect 430486 164898 460970 165134
rect 461206 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 46250 147454
rect 46486 147218 76970 147454
rect 77206 147218 107690 147454
rect 107926 147218 138410 147454
rect 138646 147218 169130 147454
rect 169366 147218 199850 147454
rect 200086 147218 230570 147454
rect 230806 147218 261290 147454
rect 261526 147218 292010 147454
rect 292246 147218 322730 147454
rect 322966 147218 353450 147454
rect 353686 147218 384170 147454
rect 384406 147218 414890 147454
rect 415126 147218 445610 147454
rect 445846 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 46250 147134
rect 46486 146898 76970 147134
rect 77206 146898 107690 147134
rect 107926 146898 138410 147134
rect 138646 146898 169130 147134
rect 169366 146898 199850 147134
rect 200086 146898 230570 147134
rect 230806 146898 261290 147134
rect 261526 146898 292010 147134
rect 292246 146898 322730 147134
rect 322966 146898 353450 147134
rect 353686 146898 384170 147134
rect 384406 146898 414890 147134
rect 415126 146898 445610 147134
rect 445846 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 61610 129454
rect 61846 129218 92330 129454
rect 92566 129218 123050 129454
rect 123286 129218 153770 129454
rect 154006 129218 184490 129454
rect 184726 129218 215210 129454
rect 215446 129218 245930 129454
rect 246166 129218 276650 129454
rect 276886 129218 307370 129454
rect 307606 129218 338090 129454
rect 338326 129218 368810 129454
rect 369046 129218 399530 129454
rect 399766 129218 430250 129454
rect 430486 129218 460970 129454
rect 461206 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 61610 129134
rect 61846 128898 92330 129134
rect 92566 128898 123050 129134
rect 123286 128898 153770 129134
rect 154006 128898 184490 129134
rect 184726 128898 215210 129134
rect 215446 128898 245930 129134
rect 246166 128898 276650 129134
rect 276886 128898 307370 129134
rect 307606 128898 338090 129134
rect 338326 128898 368810 129134
rect 369046 128898 399530 129134
rect 399766 128898 430250 129134
rect 430486 128898 460970 129134
rect 461206 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 46250 111454
rect 46486 111218 76970 111454
rect 77206 111218 107690 111454
rect 107926 111218 138410 111454
rect 138646 111218 169130 111454
rect 169366 111218 199850 111454
rect 200086 111218 230570 111454
rect 230806 111218 261290 111454
rect 261526 111218 292010 111454
rect 292246 111218 322730 111454
rect 322966 111218 353450 111454
rect 353686 111218 384170 111454
rect 384406 111218 414890 111454
rect 415126 111218 445610 111454
rect 445846 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 46250 111134
rect 46486 110898 76970 111134
rect 77206 110898 107690 111134
rect 107926 110898 138410 111134
rect 138646 110898 169130 111134
rect 169366 110898 199850 111134
rect 200086 110898 230570 111134
rect 230806 110898 261290 111134
rect 261526 110898 292010 111134
rect 292246 110898 322730 111134
rect 322966 110898 353450 111134
rect 353686 110898 384170 111134
rect 384406 110898 414890 111134
rect 415126 110898 445610 111134
rect 445846 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 61610 93454
rect 61846 93218 92330 93454
rect 92566 93218 123050 93454
rect 123286 93218 153770 93454
rect 154006 93218 184490 93454
rect 184726 93218 215210 93454
rect 215446 93218 245930 93454
rect 246166 93218 276650 93454
rect 276886 93218 307370 93454
rect 307606 93218 338090 93454
rect 338326 93218 368810 93454
rect 369046 93218 399530 93454
rect 399766 93218 430250 93454
rect 430486 93218 460970 93454
rect 461206 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 61610 93134
rect 61846 92898 92330 93134
rect 92566 92898 123050 93134
rect 123286 92898 153770 93134
rect 154006 92898 184490 93134
rect 184726 92898 215210 93134
rect 215446 92898 245930 93134
rect 246166 92898 276650 93134
rect 276886 92898 307370 93134
rect 307606 92898 338090 93134
rect 338326 92898 368810 93134
rect 369046 92898 399530 93134
rect 399766 92898 430250 93134
rect 430486 92898 460970 93134
rect 461206 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 46250 75454
rect 46486 75218 76970 75454
rect 77206 75218 107690 75454
rect 107926 75218 138410 75454
rect 138646 75218 169130 75454
rect 169366 75218 199850 75454
rect 200086 75218 230570 75454
rect 230806 75218 261290 75454
rect 261526 75218 292010 75454
rect 292246 75218 322730 75454
rect 322966 75218 353450 75454
rect 353686 75218 384170 75454
rect 384406 75218 414890 75454
rect 415126 75218 445610 75454
rect 445846 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 46250 75134
rect 46486 74898 76970 75134
rect 77206 74898 107690 75134
rect 107926 74898 138410 75134
rect 138646 74898 169130 75134
rect 169366 74898 199850 75134
rect 200086 74898 230570 75134
rect 230806 74898 261290 75134
rect 261526 74898 292010 75134
rect 292246 74898 322730 75134
rect 322966 74898 353450 75134
rect 353686 74898 384170 75134
rect 384406 74898 414890 75134
rect 415126 74898 445610 75134
rect 445846 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 61610 57454
rect 61846 57218 92330 57454
rect 92566 57218 123050 57454
rect 123286 57218 153770 57454
rect 154006 57218 184490 57454
rect 184726 57218 215210 57454
rect 215446 57218 245930 57454
rect 246166 57218 276650 57454
rect 276886 57218 307370 57454
rect 307606 57218 338090 57454
rect 338326 57218 368810 57454
rect 369046 57218 399530 57454
rect 399766 57218 430250 57454
rect 430486 57218 460970 57454
rect 461206 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 61610 57134
rect 61846 56898 92330 57134
rect 92566 56898 123050 57134
rect 123286 56898 153770 57134
rect 154006 56898 184490 57134
rect 184726 56898 215210 57134
rect 215446 56898 245930 57134
rect 246166 56898 276650 57134
rect 276886 56898 307370 57134
rect 307606 56898 338090 57134
rect 338326 56898 368810 57134
rect 369046 56898 399530 57134
rect 399766 56898 430250 57134
rect 430486 56898 460970 57134
rect 461206 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1636387369
transform 1 0 42000 0 1 42000
box 382 0 424551 426704
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 40000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 470704 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 470704 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 470704 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 470704 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 470704 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 470704 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 470704 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 470704 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 470704 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 470704 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 470704 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 40000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 470704 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 470704 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 470704 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 470704 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 470704 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 470704 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 470704 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 470704 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 470704 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 470704 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 470704 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 470704 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 40000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 470704 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 470704 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 470704 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 470704 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 470704 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 470704 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 470704 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 470704 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 470704 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 470704 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 470704 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 470704 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 40000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 470704 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 470704 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 470704 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 470704 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 470704 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 470704 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 470704 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 470704 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 470704 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 470704 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 470704 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 470704 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 40000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 470704 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 470704 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 470704 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 470704 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 470704 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 470704 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 470704 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 470704 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 470704 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 470704 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 470704 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 470704 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 40000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 470704 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 470704 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 470704 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 470704 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 470704 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 470704 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 470704 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 470704 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 470704 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 470704 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 470704 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 470704 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 40000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 470704 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 470704 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 470704 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 470704 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 470704 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 470704 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 470704 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 470704 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 470704 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 470704 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 470704 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 470704 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 40000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 470704 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 470704 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 470704 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 470704 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 470704 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 470704 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 470704 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 470704 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 470704 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 470704 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 470704 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 470704 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
