magic
tech sky130A
magscale 1 2
timestamp 1635724552
<< obsli1 >>
rect 1104 289 519403 637585
<< obsm1 >>
rect 474 8 519418 637616
<< metal2 >>
rect 2226 639200 2282 640000
rect 6734 639200 6790 640000
rect 11334 639200 11390 640000
rect 15842 639200 15898 640000
rect 20442 639200 20498 640000
rect 24950 639200 25006 640000
rect 29550 639200 29606 640000
rect 34150 639200 34206 640000
rect 38658 639200 38714 640000
rect 43258 639200 43314 640000
rect 47766 639200 47822 640000
rect 52366 639200 52422 640000
rect 56874 639200 56930 640000
rect 61474 639200 61530 640000
rect 66074 639200 66130 640000
rect 70582 639200 70638 640000
rect 75182 639200 75238 640000
rect 79690 639200 79746 640000
rect 84290 639200 84346 640000
rect 88890 639200 88946 640000
rect 93398 639200 93454 640000
rect 97998 639200 98054 640000
rect 102506 639200 102562 640000
rect 107106 639200 107162 640000
rect 111614 639200 111670 640000
rect 116214 639200 116270 640000
rect 120814 639200 120870 640000
rect 125322 639200 125378 640000
rect 129922 639200 129978 640000
rect 134430 639200 134486 640000
rect 139030 639200 139086 640000
rect 143538 639200 143594 640000
rect 148138 639200 148194 640000
rect 152738 639200 152794 640000
rect 157246 639200 157302 640000
rect 161846 639200 161902 640000
rect 166354 639200 166410 640000
rect 170954 639200 171010 640000
rect 175554 639200 175610 640000
rect 180062 639200 180118 640000
rect 184662 639200 184718 640000
rect 189170 639200 189226 640000
rect 193770 639200 193826 640000
rect 198278 639200 198334 640000
rect 202878 639200 202934 640000
rect 207478 639200 207534 640000
rect 211986 639200 212042 640000
rect 216586 639200 216642 640000
rect 221094 639200 221150 640000
rect 225694 639200 225750 640000
rect 230202 639200 230258 640000
rect 234802 639200 234858 640000
rect 239402 639200 239458 640000
rect 243910 639200 243966 640000
rect 248510 639200 248566 640000
rect 253018 639200 253074 640000
rect 257618 639200 257674 640000
rect 262218 639200 262274 640000
rect 266726 639200 266782 640000
rect 271326 639200 271382 640000
rect 275834 639200 275890 640000
rect 280434 639200 280490 640000
rect 284942 639200 284998 640000
rect 289542 639200 289598 640000
rect 294142 639200 294198 640000
rect 298650 639200 298706 640000
rect 303250 639200 303306 640000
rect 307758 639200 307814 640000
rect 312358 639200 312414 640000
rect 316866 639200 316922 640000
rect 321466 639200 321522 640000
rect 326066 639200 326122 640000
rect 330574 639200 330630 640000
rect 335174 639200 335230 640000
rect 339682 639200 339738 640000
rect 344282 639200 344338 640000
rect 348882 639200 348938 640000
rect 353390 639200 353446 640000
rect 357990 639200 358046 640000
rect 362498 639200 362554 640000
rect 367098 639200 367154 640000
rect 371606 639200 371662 640000
rect 376206 639200 376262 640000
rect 380806 639200 380862 640000
rect 385314 639200 385370 640000
rect 389914 639200 389970 640000
rect 394422 639200 394478 640000
rect 399022 639200 399078 640000
rect 403530 639200 403586 640000
rect 408130 639200 408186 640000
rect 412730 639200 412786 640000
rect 417238 639200 417294 640000
rect 421838 639200 421894 640000
rect 426346 639200 426402 640000
rect 430946 639200 431002 640000
rect 435546 639200 435602 640000
rect 440054 639200 440110 640000
rect 444654 639200 444710 640000
rect 449162 639200 449218 640000
rect 453762 639200 453818 640000
rect 458270 639200 458326 640000
rect 462870 639200 462926 640000
rect 467470 639200 467526 640000
rect 471978 639200 472034 640000
rect 476578 639200 476634 640000
rect 481086 639200 481142 640000
rect 485686 639200 485742 640000
rect 490194 639200 490250 640000
rect 494794 639200 494850 640000
rect 499394 639200 499450 640000
rect 503902 639200 503958 640000
rect 508502 639200 508558 640000
rect 513010 639200 513066 640000
rect 517610 639200 517666 640000
rect 478 0 534 800
rect 1490 0 1546 800
rect 2502 0 2558 800
rect 3606 0 3662 800
rect 4618 0 4674 800
rect 5722 0 5778 800
rect 6734 0 6790 800
rect 7838 0 7894 800
rect 8850 0 8906 800
rect 9954 0 10010 800
rect 10966 0 11022 800
rect 12070 0 12126 800
rect 13082 0 13138 800
rect 14186 0 14242 800
rect 15198 0 15254 800
rect 16210 0 16266 800
rect 17314 0 17370 800
rect 18326 0 18382 800
rect 19430 0 19486 800
rect 20442 0 20498 800
rect 21546 0 21602 800
rect 22558 0 22614 800
rect 23662 0 23718 800
rect 24674 0 24730 800
rect 25778 0 25834 800
rect 26790 0 26846 800
rect 27894 0 27950 800
rect 28906 0 28962 800
rect 30010 0 30066 800
rect 31022 0 31078 800
rect 32034 0 32090 800
rect 33138 0 33194 800
rect 34150 0 34206 800
rect 35254 0 35310 800
rect 36266 0 36322 800
rect 37370 0 37426 800
rect 38382 0 38438 800
rect 39486 0 39542 800
rect 40498 0 40554 800
rect 41602 0 41658 800
rect 42614 0 42670 800
rect 43718 0 43774 800
rect 44730 0 44786 800
rect 45742 0 45798 800
rect 46846 0 46902 800
rect 47858 0 47914 800
rect 48962 0 49018 800
rect 49974 0 50030 800
rect 51078 0 51134 800
rect 52090 0 52146 800
rect 53194 0 53250 800
rect 54206 0 54262 800
rect 55310 0 55366 800
rect 56322 0 56378 800
rect 57426 0 57482 800
rect 58438 0 58494 800
rect 59542 0 59598 800
rect 60554 0 60610 800
rect 61566 0 61622 800
rect 62670 0 62726 800
rect 63682 0 63738 800
rect 64786 0 64842 800
rect 65798 0 65854 800
rect 66902 0 66958 800
rect 67914 0 67970 800
rect 69018 0 69074 800
rect 70030 0 70086 800
rect 71134 0 71190 800
rect 72146 0 72202 800
rect 73250 0 73306 800
rect 74262 0 74318 800
rect 75274 0 75330 800
rect 76378 0 76434 800
rect 77390 0 77446 800
rect 78494 0 78550 800
rect 79506 0 79562 800
rect 80610 0 80666 800
rect 81622 0 81678 800
rect 82726 0 82782 800
rect 83738 0 83794 800
rect 84842 0 84898 800
rect 85854 0 85910 800
rect 86958 0 87014 800
rect 87970 0 88026 800
rect 89074 0 89130 800
rect 90086 0 90142 800
rect 91098 0 91154 800
rect 92202 0 92258 800
rect 93214 0 93270 800
rect 94318 0 94374 800
rect 95330 0 95386 800
rect 96434 0 96490 800
rect 97446 0 97502 800
rect 98550 0 98606 800
rect 99562 0 99618 800
rect 100666 0 100722 800
rect 101678 0 101734 800
rect 102782 0 102838 800
rect 103794 0 103850 800
rect 104806 0 104862 800
rect 105910 0 105966 800
rect 106922 0 106978 800
rect 108026 0 108082 800
rect 109038 0 109094 800
rect 110142 0 110198 800
rect 111154 0 111210 800
rect 112258 0 112314 800
rect 113270 0 113326 800
rect 114374 0 114430 800
rect 115386 0 115442 800
rect 116490 0 116546 800
rect 117502 0 117558 800
rect 118606 0 118662 800
rect 119618 0 119674 800
rect 120630 0 120686 800
rect 121734 0 121790 800
rect 122746 0 122802 800
rect 123850 0 123906 800
rect 124862 0 124918 800
rect 125966 0 126022 800
rect 126978 0 127034 800
rect 128082 0 128138 800
rect 129094 0 129150 800
rect 130198 0 130254 800
rect 131210 0 131266 800
rect 132314 0 132370 800
rect 133326 0 133382 800
rect 134338 0 134394 800
rect 135442 0 135498 800
rect 136454 0 136510 800
rect 137558 0 137614 800
rect 138570 0 138626 800
rect 139674 0 139730 800
rect 140686 0 140742 800
rect 141790 0 141846 800
rect 142802 0 142858 800
rect 143906 0 143962 800
rect 144918 0 144974 800
rect 146022 0 146078 800
rect 147034 0 147090 800
rect 148138 0 148194 800
rect 149150 0 149206 800
rect 150162 0 150218 800
rect 151266 0 151322 800
rect 152278 0 152334 800
rect 153382 0 153438 800
rect 154394 0 154450 800
rect 155498 0 155554 800
rect 156510 0 156566 800
rect 157614 0 157670 800
rect 158626 0 158682 800
rect 159730 0 159786 800
rect 160742 0 160798 800
rect 161846 0 161902 800
rect 162858 0 162914 800
rect 163870 0 163926 800
rect 164974 0 165030 800
rect 165986 0 166042 800
rect 167090 0 167146 800
rect 168102 0 168158 800
rect 169206 0 169262 800
rect 170218 0 170274 800
rect 171322 0 171378 800
rect 172334 0 172390 800
rect 173438 0 173494 800
rect 174450 0 174506 800
rect 175554 0 175610 800
rect 176566 0 176622 800
rect 177670 0 177726 800
rect 178682 0 178738 800
rect 179694 0 179750 800
rect 180798 0 180854 800
rect 181810 0 181866 800
rect 182914 0 182970 800
rect 183926 0 183982 800
rect 185030 0 185086 800
rect 186042 0 186098 800
rect 187146 0 187202 800
rect 188158 0 188214 800
rect 189262 0 189318 800
rect 190274 0 190330 800
rect 191378 0 191434 800
rect 192390 0 192446 800
rect 193494 0 193550 800
rect 194506 0 194562 800
rect 195518 0 195574 800
rect 196622 0 196678 800
rect 197634 0 197690 800
rect 198738 0 198794 800
rect 199750 0 199806 800
rect 200854 0 200910 800
rect 201866 0 201922 800
rect 202970 0 203026 800
rect 203982 0 204038 800
rect 205086 0 205142 800
rect 206098 0 206154 800
rect 207202 0 207258 800
rect 208214 0 208270 800
rect 209226 0 209282 800
rect 210330 0 210386 800
rect 211342 0 211398 800
rect 212446 0 212502 800
rect 213458 0 213514 800
rect 214562 0 214618 800
rect 215574 0 215630 800
rect 216678 0 216734 800
rect 217690 0 217746 800
rect 218794 0 218850 800
rect 219806 0 219862 800
rect 220910 0 220966 800
rect 221922 0 221978 800
rect 223026 0 223082 800
rect 224038 0 224094 800
rect 225050 0 225106 800
rect 226154 0 226210 800
rect 227166 0 227222 800
rect 228270 0 228326 800
rect 229282 0 229338 800
rect 230386 0 230442 800
rect 231398 0 231454 800
rect 232502 0 232558 800
rect 233514 0 233570 800
rect 234618 0 234674 800
rect 235630 0 235686 800
rect 236734 0 236790 800
rect 237746 0 237802 800
rect 238758 0 238814 800
rect 239862 0 239918 800
rect 240874 0 240930 800
rect 241978 0 242034 800
rect 242990 0 243046 800
rect 244094 0 244150 800
rect 245106 0 245162 800
rect 246210 0 246266 800
rect 247222 0 247278 800
rect 248326 0 248382 800
rect 249338 0 249394 800
rect 250442 0 250498 800
rect 251454 0 251510 800
rect 252558 0 252614 800
rect 253570 0 253626 800
rect 254582 0 254638 800
rect 255686 0 255742 800
rect 256698 0 256754 800
rect 257802 0 257858 800
rect 258814 0 258870 800
rect 259918 0 259974 800
rect 260930 0 260986 800
rect 262034 0 262090 800
rect 263046 0 263102 800
rect 264150 0 264206 800
rect 265162 0 265218 800
rect 266266 0 266322 800
rect 267278 0 267334 800
rect 268290 0 268346 800
rect 269394 0 269450 800
rect 270406 0 270462 800
rect 271510 0 271566 800
rect 272522 0 272578 800
rect 273626 0 273682 800
rect 274638 0 274694 800
rect 275742 0 275798 800
rect 276754 0 276810 800
rect 277858 0 277914 800
rect 278870 0 278926 800
rect 279974 0 280030 800
rect 280986 0 281042 800
rect 282090 0 282146 800
rect 283102 0 283158 800
rect 284114 0 284170 800
rect 285218 0 285274 800
rect 286230 0 286286 800
rect 287334 0 287390 800
rect 288346 0 288402 800
rect 289450 0 289506 800
rect 290462 0 290518 800
rect 291566 0 291622 800
rect 292578 0 292634 800
rect 293682 0 293738 800
rect 294694 0 294750 800
rect 295798 0 295854 800
rect 296810 0 296866 800
rect 297822 0 297878 800
rect 298926 0 298982 800
rect 299938 0 299994 800
rect 301042 0 301098 800
rect 302054 0 302110 800
rect 303158 0 303214 800
rect 304170 0 304226 800
rect 305274 0 305330 800
rect 306286 0 306342 800
rect 307390 0 307446 800
rect 308402 0 308458 800
rect 309506 0 309562 800
rect 310518 0 310574 800
rect 311622 0 311678 800
rect 312634 0 312690 800
rect 313646 0 313702 800
rect 314750 0 314806 800
rect 315762 0 315818 800
rect 316866 0 316922 800
rect 317878 0 317934 800
rect 318982 0 319038 800
rect 319994 0 320050 800
rect 321098 0 321154 800
rect 322110 0 322166 800
rect 323214 0 323270 800
rect 324226 0 324282 800
rect 325330 0 325386 800
rect 326342 0 326398 800
rect 327354 0 327410 800
rect 328458 0 328514 800
rect 329470 0 329526 800
rect 330574 0 330630 800
rect 331586 0 331642 800
rect 332690 0 332746 800
rect 333702 0 333758 800
rect 334806 0 334862 800
rect 335818 0 335874 800
rect 336922 0 336978 800
rect 337934 0 337990 800
rect 339038 0 339094 800
rect 340050 0 340106 800
rect 341154 0 341210 800
rect 342166 0 342222 800
rect 343178 0 343234 800
rect 344282 0 344338 800
rect 345294 0 345350 800
rect 346398 0 346454 800
rect 347410 0 347466 800
rect 348514 0 348570 800
rect 349526 0 349582 800
rect 350630 0 350686 800
rect 351642 0 351698 800
rect 352746 0 352802 800
rect 353758 0 353814 800
rect 354862 0 354918 800
rect 355874 0 355930 800
rect 356978 0 357034 800
rect 357990 0 358046 800
rect 359002 0 359058 800
rect 360106 0 360162 800
rect 361118 0 361174 800
rect 362222 0 362278 800
rect 363234 0 363290 800
rect 364338 0 364394 800
rect 365350 0 365406 800
rect 366454 0 366510 800
rect 367466 0 367522 800
rect 368570 0 368626 800
rect 369582 0 369638 800
rect 370686 0 370742 800
rect 371698 0 371754 800
rect 372710 0 372766 800
rect 373814 0 373870 800
rect 374826 0 374882 800
rect 375930 0 375986 800
rect 376942 0 376998 800
rect 378046 0 378102 800
rect 379058 0 379114 800
rect 380162 0 380218 800
rect 381174 0 381230 800
rect 382278 0 382334 800
rect 383290 0 383346 800
rect 384394 0 384450 800
rect 385406 0 385462 800
rect 386510 0 386566 800
rect 387522 0 387578 800
rect 388534 0 388590 800
rect 389638 0 389694 800
rect 390650 0 390706 800
rect 391754 0 391810 800
rect 392766 0 392822 800
rect 393870 0 393926 800
rect 394882 0 394938 800
rect 395986 0 396042 800
rect 396998 0 397054 800
rect 398102 0 398158 800
rect 399114 0 399170 800
rect 400218 0 400274 800
rect 401230 0 401286 800
rect 402242 0 402298 800
rect 403346 0 403402 800
rect 404358 0 404414 800
rect 405462 0 405518 800
rect 406474 0 406530 800
rect 407578 0 407634 800
rect 408590 0 408646 800
rect 409694 0 409750 800
rect 410706 0 410762 800
rect 411810 0 411866 800
rect 412822 0 412878 800
rect 413926 0 413982 800
rect 414938 0 414994 800
rect 416042 0 416098 800
rect 417054 0 417110 800
rect 418066 0 418122 800
rect 419170 0 419226 800
rect 420182 0 420238 800
rect 421286 0 421342 800
rect 422298 0 422354 800
rect 423402 0 423458 800
rect 424414 0 424470 800
rect 425518 0 425574 800
rect 426530 0 426586 800
rect 427634 0 427690 800
rect 428646 0 428702 800
rect 429750 0 429806 800
rect 430762 0 430818 800
rect 431774 0 431830 800
rect 432878 0 432934 800
rect 433890 0 433946 800
rect 434994 0 435050 800
rect 436006 0 436062 800
rect 437110 0 437166 800
rect 438122 0 438178 800
rect 439226 0 439282 800
rect 440238 0 440294 800
rect 441342 0 441398 800
rect 442354 0 442410 800
rect 443458 0 443514 800
rect 444470 0 444526 800
rect 445574 0 445630 800
rect 446586 0 446642 800
rect 447598 0 447654 800
rect 448702 0 448758 800
rect 449714 0 449770 800
rect 450818 0 450874 800
rect 451830 0 451886 800
rect 452934 0 452990 800
rect 453946 0 454002 800
rect 455050 0 455106 800
rect 456062 0 456118 800
rect 457166 0 457222 800
rect 458178 0 458234 800
rect 459282 0 459338 800
rect 460294 0 460350 800
rect 461306 0 461362 800
rect 462410 0 462466 800
rect 463422 0 463478 800
rect 464526 0 464582 800
rect 465538 0 465594 800
rect 466642 0 466698 800
rect 467654 0 467710 800
rect 468758 0 468814 800
rect 469770 0 469826 800
rect 470874 0 470930 800
rect 471886 0 471942 800
rect 472990 0 473046 800
rect 474002 0 474058 800
rect 475106 0 475162 800
rect 476118 0 476174 800
rect 477130 0 477186 800
rect 478234 0 478290 800
rect 479246 0 479302 800
rect 480350 0 480406 800
rect 481362 0 481418 800
rect 482466 0 482522 800
rect 483478 0 483534 800
rect 484582 0 484638 800
rect 485594 0 485650 800
rect 486698 0 486754 800
rect 487710 0 487766 800
rect 488814 0 488870 800
rect 489826 0 489882 800
rect 490838 0 490894 800
rect 491942 0 491998 800
rect 492954 0 493010 800
rect 494058 0 494114 800
rect 495070 0 495126 800
rect 496174 0 496230 800
rect 497186 0 497242 800
rect 498290 0 498346 800
rect 499302 0 499358 800
rect 500406 0 500462 800
rect 501418 0 501474 800
rect 502522 0 502578 800
rect 503534 0 503590 800
rect 504638 0 504694 800
rect 505650 0 505706 800
rect 506662 0 506718 800
rect 507766 0 507822 800
rect 508778 0 508834 800
rect 509882 0 509938 800
rect 510894 0 510950 800
rect 511998 0 512054 800
rect 513010 0 513066 800
rect 514114 0 514170 800
rect 515126 0 515182 800
rect 516230 0 516286 800
rect 517242 0 517298 800
rect 518346 0 518402 800
rect 519358 0 519414 800
<< obsm2 >>
rect 480 639144 2170 639282
rect 2338 639144 6678 639282
rect 6846 639144 11278 639282
rect 11446 639144 15786 639282
rect 15954 639144 20386 639282
rect 20554 639144 24894 639282
rect 25062 639144 29494 639282
rect 29662 639144 34094 639282
rect 34262 639144 38602 639282
rect 38770 639144 43202 639282
rect 43370 639144 47710 639282
rect 47878 639144 52310 639282
rect 52478 639144 56818 639282
rect 56986 639144 61418 639282
rect 61586 639144 66018 639282
rect 66186 639144 70526 639282
rect 70694 639144 75126 639282
rect 75294 639144 79634 639282
rect 79802 639144 84234 639282
rect 84402 639144 88834 639282
rect 89002 639144 93342 639282
rect 93510 639144 97942 639282
rect 98110 639144 102450 639282
rect 102618 639144 107050 639282
rect 107218 639144 111558 639282
rect 111726 639144 116158 639282
rect 116326 639144 120758 639282
rect 120926 639144 125266 639282
rect 125434 639144 129866 639282
rect 130034 639144 134374 639282
rect 134542 639144 138974 639282
rect 139142 639144 143482 639282
rect 143650 639144 148082 639282
rect 148250 639144 152682 639282
rect 152850 639144 157190 639282
rect 157358 639144 161790 639282
rect 161958 639144 166298 639282
rect 166466 639144 170898 639282
rect 171066 639144 175498 639282
rect 175666 639144 180006 639282
rect 180174 639144 184606 639282
rect 184774 639144 189114 639282
rect 189282 639144 193714 639282
rect 193882 639144 198222 639282
rect 198390 639144 202822 639282
rect 202990 639144 207422 639282
rect 207590 639144 211930 639282
rect 212098 639144 216530 639282
rect 216698 639144 221038 639282
rect 221206 639144 225638 639282
rect 225806 639144 230146 639282
rect 230314 639144 234746 639282
rect 234914 639144 239346 639282
rect 239514 639144 243854 639282
rect 244022 639144 248454 639282
rect 248622 639144 252962 639282
rect 253130 639144 257562 639282
rect 257730 639144 262162 639282
rect 262330 639144 266670 639282
rect 266838 639144 271270 639282
rect 271438 639144 275778 639282
rect 275946 639144 280378 639282
rect 280546 639144 284886 639282
rect 285054 639144 289486 639282
rect 289654 639144 294086 639282
rect 294254 639144 298594 639282
rect 298762 639144 303194 639282
rect 303362 639144 307702 639282
rect 307870 639144 312302 639282
rect 312470 639144 316810 639282
rect 316978 639144 321410 639282
rect 321578 639144 326010 639282
rect 326178 639144 330518 639282
rect 330686 639144 335118 639282
rect 335286 639144 339626 639282
rect 339794 639144 344226 639282
rect 344394 639144 348826 639282
rect 348994 639144 353334 639282
rect 353502 639144 357934 639282
rect 358102 639144 362442 639282
rect 362610 639144 367042 639282
rect 367210 639144 371550 639282
rect 371718 639144 376150 639282
rect 376318 639144 380750 639282
rect 380918 639144 385258 639282
rect 385426 639144 389858 639282
rect 390026 639144 394366 639282
rect 394534 639144 398966 639282
rect 399134 639144 403474 639282
rect 403642 639144 408074 639282
rect 408242 639144 412674 639282
rect 412842 639144 417182 639282
rect 417350 639144 421782 639282
rect 421950 639144 426290 639282
rect 426458 639144 430890 639282
rect 431058 639144 435490 639282
rect 435658 639144 439998 639282
rect 440166 639144 444598 639282
rect 444766 639144 449106 639282
rect 449274 639144 453706 639282
rect 453874 639144 458214 639282
rect 458382 639144 462814 639282
rect 462982 639144 467414 639282
rect 467582 639144 471922 639282
rect 472090 639144 476522 639282
rect 476690 639144 481030 639282
rect 481198 639144 485630 639282
rect 485798 639144 490138 639282
rect 490306 639144 494738 639282
rect 494906 639144 499338 639282
rect 499506 639144 503846 639282
rect 504014 639144 508446 639282
rect 508614 639144 512954 639282
rect 513122 639144 517554 639282
rect 517722 639144 519412 639282
rect 480 856 519412 639144
rect 590 2 1434 856
rect 1602 2 2446 856
rect 2614 2 3550 856
rect 3718 2 4562 856
rect 4730 2 5666 856
rect 5834 2 6678 856
rect 6846 2 7782 856
rect 7950 2 8794 856
rect 8962 2 9898 856
rect 10066 2 10910 856
rect 11078 2 12014 856
rect 12182 2 13026 856
rect 13194 2 14130 856
rect 14298 2 15142 856
rect 15310 2 16154 856
rect 16322 2 17258 856
rect 17426 2 18270 856
rect 18438 2 19374 856
rect 19542 2 20386 856
rect 20554 2 21490 856
rect 21658 2 22502 856
rect 22670 2 23606 856
rect 23774 2 24618 856
rect 24786 2 25722 856
rect 25890 2 26734 856
rect 26902 2 27838 856
rect 28006 2 28850 856
rect 29018 2 29954 856
rect 30122 2 30966 856
rect 31134 2 31978 856
rect 32146 2 33082 856
rect 33250 2 34094 856
rect 34262 2 35198 856
rect 35366 2 36210 856
rect 36378 2 37314 856
rect 37482 2 38326 856
rect 38494 2 39430 856
rect 39598 2 40442 856
rect 40610 2 41546 856
rect 41714 2 42558 856
rect 42726 2 43662 856
rect 43830 2 44674 856
rect 44842 2 45686 856
rect 45854 2 46790 856
rect 46958 2 47802 856
rect 47970 2 48906 856
rect 49074 2 49918 856
rect 50086 2 51022 856
rect 51190 2 52034 856
rect 52202 2 53138 856
rect 53306 2 54150 856
rect 54318 2 55254 856
rect 55422 2 56266 856
rect 56434 2 57370 856
rect 57538 2 58382 856
rect 58550 2 59486 856
rect 59654 2 60498 856
rect 60666 2 61510 856
rect 61678 2 62614 856
rect 62782 2 63626 856
rect 63794 2 64730 856
rect 64898 2 65742 856
rect 65910 2 66846 856
rect 67014 2 67858 856
rect 68026 2 68962 856
rect 69130 2 69974 856
rect 70142 2 71078 856
rect 71246 2 72090 856
rect 72258 2 73194 856
rect 73362 2 74206 856
rect 74374 2 75218 856
rect 75386 2 76322 856
rect 76490 2 77334 856
rect 77502 2 78438 856
rect 78606 2 79450 856
rect 79618 2 80554 856
rect 80722 2 81566 856
rect 81734 2 82670 856
rect 82838 2 83682 856
rect 83850 2 84786 856
rect 84954 2 85798 856
rect 85966 2 86902 856
rect 87070 2 87914 856
rect 88082 2 89018 856
rect 89186 2 90030 856
rect 90198 2 91042 856
rect 91210 2 92146 856
rect 92314 2 93158 856
rect 93326 2 94262 856
rect 94430 2 95274 856
rect 95442 2 96378 856
rect 96546 2 97390 856
rect 97558 2 98494 856
rect 98662 2 99506 856
rect 99674 2 100610 856
rect 100778 2 101622 856
rect 101790 2 102726 856
rect 102894 2 103738 856
rect 103906 2 104750 856
rect 104918 2 105854 856
rect 106022 2 106866 856
rect 107034 2 107970 856
rect 108138 2 108982 856
rect 109150 2 110086 856
rect 110254 2 111098 856
rect 111266 2 112202 856
rect 112370 2 113214 856
rect 113382 2 114318 856
rect 114486 2 115330 856
rect 115498 2 116434 856
rect 116602 2 117446 856
rect 117614 2 118550 856
rect 118718 2 119562 856
rect 119730 2 120574 856
rect 120742 2 121678 856
rect 121846 2 122690 856
rect 122858 2 123794 856
rect 123962 2 124806 856
rect 124974 2 125910 856
rect 126078 2 126922 856
rect 127090 2 128026 856
rect 128194 2 129038 856
rect 129206 2 130142 856
rect 130310 2 131154 856
rect 131322 2 132258 856
rect 132426 2 133270 856
rect 133438 2 134282 856
rect 134450 2 135386 856
rect 135554 2 136398 856
rect 136566 2 137502 856
rect 137670 2 138514 856
rect 138682 2 139618 856
rect 139786 2 140630 856
rect 140798 2 141734 856
rect 141902 2 142746 856
rect 142914 2 143850 856
rect 144018 2 144862 856
rect 145030 2 145966 856
rect 146134 2 146978 856
rect 147146 2 148082 856
rect 148250 2 149094 856
rect 149262 2 150106 856
rect 150274 2 151210 856
rect 151378 2 152222 856
rect 152390 2 153326 856
rect 153494 2 154338 856
rect 154506 2 155442 856
rect 155610 2 156454 856
rect 156622 2 157558 856
rect 157726 2 158570 856
rect 158738 2 159674 856
rect 159842 2 160686 856
rect 160854 2 161790 856
rect 161958 2 162802 856
rect 162970 2 163814 856
rect 163982 2 164918 856
rect 165086 2 165930 856
rect 166098 2 167034 856
rect 167202 2 168046 856
rect 168214 2 169150 856
rect 169318 2 170162 856
rect 170330 2 171266 856
rect 171434 2 172278 856
rect 172446 2 173382 856
rect 173550 2 174394 856
rect 174562 2 175498 856
rect 175666 2 176510 856
rect 176678 2 177614 856
rect 177782 2 178626 856
rect 178794 2 179638 856
rect 179806 2 180742 856
rect 180910 2 181754 856
rect 181922 2 182858 856
rect 183026 2 183870 856
rect 184038 2 184974 856
rect 185142 2 185986 856
rect 186154 2 187090 856
rect 187258 2 188102 856
rect 188270 2 189206 856
rect 189374 2 190218 856
rect 190386 2 191322 856
rect 191490 2 192334 856
rect 192502 2 193438 856
rect 193606 2 194450 856
rect 194618 2 195462 856
rect 195630 2 196566 856
rect 196734 2 197578 856
rect 197746 2 198682 856
rect 198850 2 199694 856
rect 199862 2 200798 856
rect 200966 2 201810 856
rect 201978 2 202914 856
rect 203082 2 203926 856
rect 204094 2 205030 856
rect 205198 2 206042 856
rect 206210 2 207146 856
rect 207314 2 208158 856
rect 208326 2 209170 856
rect 209338 2 210274 856
rect 210442 2 211286 856
rect 211454 2 212390 856
rect 212558 2 213402 856
rect 213570 2 214506 856
rect 214674 2 215518 856
rect 215686 2 216622 856
rect 216790 2 217634 856
rect 217802 2 218738 856
rect 218906 2 219750 856
rect 219918 2 220854 856
rect 221022 2 221866 856
rect 222034 2 222970 856
rect 223138 2 223982 856
rect 224150 2 224994 856
rect 225162 2 226098 856
rect 226266 2 227110 856
rect 227278 2 228214 856
rect 228382 2 229226 856
rect 229394 2 230330 856
rect 230498 2 231342 856
rect 231510 2 232446 856
rect 232614 2 233458 856
rect 233626 2 234562 856
rect 234730 2 235574 856
rect 235742 2 236678 856
rect 236846 2 237690 856
rect 237858 2 238702 856
rect 238870 2 239806 856
rect 239974 2 240818 856
rect 240986 2 241922 856
rect 242090 2 242934 856
rect 243102 2 244038 856
rect 244206 2 245050 856
rect 245218 2 246154 856
rect 246322 2 247166 856
rect 247334 2 248270 856
rect 248438 2 249282 856
rect 249450 2 250386 856
rect 250554 2 251398 856
rect 251566 2 252502 856
rect 252670 2 253514 856
rect 253682 2 254526 856
rect 254694 2 255630 856
rect 255798 2 256642 856
rect 256810 2 257746 856
rect 257914 2 258758 856
rect 258926 2 259862 856
rect 260030 2 260874 856
rect 261042 2 261978 856
rect 262146 2 262990 856
rect 263158 2 264094 856
rect 264262 2 265106 856
rect 265274 2 266210 856
rect 266378 2 267222 856
rect 267390 2 268234 856
rect 268402 2 269338 856
rect 269506 2 270350 856
rect 270518 2 271454 856
rect 271622 2 272466 856
rect 272634 2 273570 856
rect 273738 2 274582 856
rect 274750 2 275686 856
rect 275854 2 276698 856
rect 276866 2 277802 856
rect 277970 2 278814 856
rect 278982 2 279918 856
rect 280086 2 280930 856
rect 281098 2 282034 856
rect 282202 2 283046 856
rect 283214 2 284058 856
rect 284226 2 285162 856
rect 285330 2 286174 856
rect 286342 2 287278 856
rect 287446 2 288290 856
rect 288458 2 289394 856
rect 289562 2 290406 856
rect 290574 2 291510 856
rect 291678 2 292522 856
rect 292690 2 293626 856
rect 293794 2 294638 856
rect 294806 2 295742 856
rect 295910 2 296754 856
rect 296922 2 297766 856
rect 297934 2 298870 856
rect 299038 2 299882 856
rect 300050 2 300986 856
rect 301154 2 301998 856
rect 302166 2 303102 856
rect 303270 2 304114 856
rect 304282 2 305218 856
rect 305386 2 306230 856
rect 306398 2 307334 856
rect 307502 2 308346 856
rect 308514 2 309450 856
rect 309618 2 310462 856
rect 310630 2 311566 856
rect 311734 2 312578 856
rect 312746 2 313590 856
rect 313758 2 314694 856
rect 314862 2 315706 856
rect 315874 2 316810 856
rect 316978 2 317822 856
rect 317990 2 318926 856
rect 319094 2 319938 856
rect 320106 2 321042 856
rect 321210 2 322054 856
rect 322222 2 323158 856
rect 323326 2 324170 856
rect 324338 2 325274 856
rect 325442 2 326286 856
rect 326454 2 327298 856
rect 327466 2 328402 856
rect 328570 2 329414 856
rect 329582 2 330518 856
rect 330686 2 331530 856
rect 331698 2 332634 856
rect 332802 2 333646 856
rect 333814 2 334750 856
rect 334918 2 335762 856
rect 335930 2 336866 856
rect 337034 2 337878 856
rect 338046 2 338982 856
rect 339150 2 339994 856
rect 340162 2 341098 856
rect 341266 2 342110 856
rect 342278 2 343122 856
rect 343290 2 344226 856
rect 344394 2 345238 856
rect 345406 2 346342 856
rect 346510 2 347354 856
rect 347522 2 348458 856
rect 348626 2 349470 856
rect 349638 2 350574 856
rect 350742 2 351586 856
rect 351754 2 352690 856
rect 352858 2 353702 856
rect 353870 2 354806 856
rect 354974 2 355818 856
rect 355986 2 356922 856
rect 357090 2 357934 856
rect 358102 2 358946 856
rect 359114 2 360050 856
rect 360218 2 361062 856
rect 361230 2 362166 856
rect 362334 2 363178 856
rect 363346 2 364282 856
rect 364450 2 365294 856
rect 365462 2 366398 856
rect 366566 2 367410 856
rect 367578 2 368514 856
rect 368682 2 369526 856
rect 369694 2 370630 856
rect 370798 2 371642 856
rect 371810 2 372654 856
rect 372822 2 373758 856
rect 373926 2 374770 856
rect 374938 2 375874 856
rect 376042 2 376886 856
rect 377054 2 377990 856
rect 378158 2 379002 856
rect 379170 2 380106 856
rect 380274 2 381118 856
rect 381286 2 382222 856
rect 382390 2 383234 856
rect 383402 2 384338 856
rect 384506 2 385350 856
rect 385518 2 386454 856
rect 386622 2 387466 856
rect 387634 2 388478 856
rect 388646 2 389582 856
rect 389750 2 390594 856
rect 390762 2 391698 856
rect 391866 2 392710 856
rect 392878 2 393814 856
rect 393982 2 394826 856
rect 394994 2 395930 856
rect 396098 2 396942 856
rect 397110 2 398046 856
rect 398214 2 399058 856
rect 399226 2 400162 856
rect 400330 2 401174 856
rect 401342 2 402186 856
rect 402354 2 403290 856
rect 403458 2 404302 856
rect 404470 2 405406 856
rect 405574 2 406418 856
rect 406586 2 407522 856
rect 407690 2 408534 856
rect 408702 2 409638 856
rect 409806 2 410650 856
rect 410818 2 411754 856
rect 411922 2 412766 856
rect 412934 2 413870 856
rect 414038 2 414882 856
rect 415050 2 415986 856
rect 416154 2 416998 856
rect 417166 2 418010 856
rect 418178 2 419114 856
rect 419282 2 420126 856
rect 420294 2 421230 856
rect 421398 2 422242 856
rect 422410 2 423346 856
rect 423514 2 424358 856
rect 424526 2 425462 856
rect 425630 2 426474 856
rect 426642 2 427578 856
rect 427746 2 428590 856
rect 428758 2 429694 856
rect 429862 2 430706 856
rect 430874 2 431718 856
rect 431886 2 432822 856
rect 432990 2 433834 856
rect 434002 2 434938 856
rect 435106 2 435950 856
rect 436118 2 437054 856
rect 437222 2 438066 856
rect 438234 2 439170 856
rect 439338 2 440182 856
rect 440350 2 441286 856
rect 441454 2 442298 856
rect 442466 2 443402 856
rect 443570 2 444414 856
rect 444582 2 445518 856
rect 445686 2 446530 856
rect 446698 2 447542 856
rect 447710 2 448646 856
rect 448814 2 449658 856
rect 449826 2 450762 856
rect 450930 2 451774 856
rect 451942 2 452878 856
rect 453046 2 453890 856
rect 454058 2 454994 856
rect 455162 2 456006 856
rect 456174 2 457110 856
rect 457278 2 458122 856
rect 458290 2 459226 856
rect 459394 2 460238 856
rect 460406 2 461250 856
rect 461418 2 462354 856
rect 462522 2 463366 856
rect 463534 2 464470 856
rect 464638 2 465482 856
rect 465650 2 466586 856
rect 466754 2 467598 856
rect 467766 2 468702 856
rect 468870 2 469714 856
rect 469882 2 470818 856
rect 470986 2 471830 856
rect 471998 2 472934 856
rect 473102 2 473946 856
rect 474114 2 475050 856
rect 475218 2 476062 856
rect 476230 2 477074 856
rect 477242 2 478178 856
rect 478346 2 479190 856
rect 479358 2 480294 856
rect 480462 2 481306 856
rect 481474 2 482410 856
rect 482578 2 483422 856
rect 483590 2 484526 856
rect 484694 2 485538 856
rect 485706 2 486642 856
rect 486810 2 487654 856
rect 487822 2 488758 856
rect 488926 2 489770 856
rect 489938 2 490782 856
rect 490950 2 491886 856
rect 492054 2 492898 856
rect 493066 2 494002 856
rect 494170 2 495014 856
rect 495182 2 496118 856
rect 496286 2 497130 856
rect 497298 2 498234 856
rect 498402 2 499246 856
rect 499414 2 500350 856
rect 500518 2 501362 856
rect 501530 2 502466 856
rect 502634 2 503478 856
rect 503646 2 504582 856
rect 504750 2 505594 856
rect 505762 2 506606 856
rect 506774 2 507710 856
rect 507878 2 508722 856
rect 508890 2 509826 856
rect 509994 2 510838 856
rect 511006 2 511942 856
rect 512110 2 512954 856
rect 513122 2 514058 856
rect 514226 2 515070 856
rect 515238 2 516174 856
rect 516342 2 517186 856
rect 517354 2 518290 856
rect 518458 2 519302 856
<< obsm3 >>
rect 3141 35 517763 637601
<< metal4 >>
rect 4208 2128 4528 637616
rect 19568 2128 19888 637616
rect 34928 2128 35248 637616
rect 50288 2128 50608 637616
rect 65648 2128 65968 637616
rect 81008 2128 81328 637616
rect 96368 2128 96688 637616
rect 111728 2128 112048 637616
rect 127088 2128 127408 637616
rect 142448 2128 142768 637616
rect 157808 2128 158128 637616
rect 173168 2128 173488 637616
rect 188528 2128 188848 637616
rect 203888 2128 204208 637616
rect 219248 2128 219568 637616
rect 234608 2128 234928 637616
rect 249968 2128 250288 637616
rect 265328 2128 265648 637616
rect 280688 2128 281008 637616
rect 296048 2128 296368 637616
rect 311408 2128 311728 637616
rect 326768 2128 327088 637616
rect 342128 2128 342448 637616
rect 357488 2128 357808 637616
rect 372848 2128 373168 637616
rect 388208 2128 388528 637616
rect 403568 2128 403888 637616
rect 418928 2128 419248 637616
rect 434288 2128 434608 637616
rect 449648 2128 449968 637616
rect 465008 2128 465328 637616
rect 480368 2128 480688 637616
rect 495728 2128 496048 637616
rect 511088 2128 511408 637616
<< obsm4 >>
rect 19379 3163 19488 637261
rect 19968 3163 34848 637261
rect 35328 3163 50208 637261
rect 50688 3163 65568 637261
rect 66048 3163 80928 637261
rect 81408 3163 96288 637261
rect 96768 3163 111648 637261
rect 112128 3163 127008 637261
rect 127488 3163 142368 637261
rect 142848 3163 157728 637261
rect 158208 3163 173088 637261
rect 173568 3163 188448 637261
rect 188928 3163 203808 637261
rect 204288 3163 219168 637261
rect 219648 3163 234528 637261
rect 235008 3163 249888 637261
rect 250368 3163 265248 637261
rect 265728 3163 280608 637261
rect 281088 3163 295968 637261
rect 296448 3163 311328 637261
rect 311808 3163 326688 637261
rect 327168 3163 342048 637261
rect 342528 3163 357408 637261
rect 357888 3163 372768 637261
rect 373248 3163 388128 637261
rect 388608 3163 403488 637261
rect 403968 3163 418848 637261
rect 419328 3163 434208 637261
rect 434688 3163 449568 637261
rect 450048 3163 464928 637261
rect 465408 3163 480288 637261
rect 480768 3163 495648 637261
rect 496128 3163 511008 637261
rect 511488 3163 516429 637261
<< labels >>
rlabel metal2 s 2226 639200 2282 640000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 139030 639200 139086 640000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 152738 639200 152794 640000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 166354 639200 166410 640000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 180062 639200 180118 640000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 193770 639200 193826 640000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 207478 639200 207534 640000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 221094 639200 221150 640000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 234802 639200 234858 640000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 248510 639200 248566 640000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 262218 639200 262274 640000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 15842 639200 15898 640000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 275834 639200 275890 640000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 289542 639200 289598 640000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 303250 639200 303306 640000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 316866 639200 316922 640000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 330574 639200 330630 640000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 344282 639200 344338 640000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 357990 639200 358046 640000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 371606 639200 371662 640000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 385314 639200 385370 640000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 399022 639200 399078 640000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 29550 639200 29606 640000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 412730 639200 412786 640000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 426346 639200 426402 640000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 440054 639200 440110 640000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 453762 639200 453818 640000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 467470 639200 467526 640000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 481086 639200 481142 640000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 494794 639200 494850 640000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 508502 639200 508558 640000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 43258 639200 43314 640000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 56874 639200 56930 640000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 70582 639200 70638 640000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 84290 639200 84346 640000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 97998 639200 98054 640000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 111614 639200 111670 640000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 125322 639200 125378 640000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6734 639200 6790 640000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 143538 639200 143594 640000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 157246 639200 157302 640000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 170954 639200 171010 640000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 184662 639200 184718 640000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 198278 639200 198334 640000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 211986 639200 212042 640000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 225694 639200 225750 640000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 239402 639200 239458 640000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 253018 639200 253074 640000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 266726 639200 266782 640000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 20442 639200 20498 640000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 280434 639200 280490 640000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 294142 639200 294198 640000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 307758 639200 307814 640000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 321466 639200 321522 640000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 335174 639200 335230 640000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 348882 639200 348938 640000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 362498 639200 362554 640000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 376206 639200 376262 640000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 389914 639200 389970 640000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 403530 639200 403586 640000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 34150 639200 34206 640000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 417238 639200 417294 640000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 430946 639200 431002 640000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 444654 639200 444710 640000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 458270 639200 458326 640000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 471978 639200 472034 640000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 485686 639200 485742 640000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 499394 639200 499450 640000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 513010 639200 513066 640000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 47766 639200 47822 640000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 61474 639200 61530 640000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 75182 639200 75238 640000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 88890 639200 88946 640000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 102506 639200 102562 640000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 116214 639200 116270 640000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 129922 639200 129978 640000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 11334 639200 11390 640000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 148138 639200 148194 640000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 161846 639200 161902 640000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 175554 639200 175610 640000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 189170 639200 189226 640000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 202878 639200 202934 640000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 216586 639200 216642 640000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 230202 639200 230258 640000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 243910 639200 243966 640000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 257618 639200 257674 640000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 271326 639200 271382 640000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 24950 639200 25006 640000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 284942 639200 284998 640000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 298650 639200 298706 640000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 312358 639200 312414 640000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 326066 639200 326122 640000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 339682 639200 339738 640000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 353390 639200 353446 640000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 367098 639200 367154 640000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 380806 639200 380862 640000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 394422 639200 394478 640000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 408130 639200 408186 640000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 38658 639200 38714 640000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 421838 639200 421894 640000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 435546 639200 435602 640000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 449162 639200 449218 640000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 462870 639200 462926 640000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 476578 639200 476634 640000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 490194 639200 490250 640000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 503902 639200 503958 640000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 517610 639200 517666 640000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 52366 639200 52422 640000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 66074 639200 66130 640000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 79690 639200 79746 640000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 93398 639200 93454 640000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 107106 639200 107162 640000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 120814 639200 120870 640000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 134430 639200 134486 640000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 517242 0 517298 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 518346 0 518402 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 519358 0 519414 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 428646 0 428702 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 431774 0 431830 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 434994 0 435050 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 438122 0 438178 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 441342 0 441398 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 444470 0 444526 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 447598 0 447654 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 450818 0 450874 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 453946 0 454002 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 457166 0 457222 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 460294 0 460350 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 463422 0 463478 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 466642 0 466698 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 469770 0 469826 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 472990 0 473046 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 476118 0 476174 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 479246 0 479302 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 482466 0 482522 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 485594 0 485650 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 488814 0 488870 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 491942 0 491998 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 495070 0 495126 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 498290 0 498346 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 501418 0 501474 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 504638 0 504694 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 507766 0 507822 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 510894 0 510950 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 514114 0 514170 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 181810 0 181866 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 185030 0 185086 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 203982 0 204038 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 216678 0 216734 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 219806 0 219862 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 223026 0 223082 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 226154 0 226210 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 238758 0 238814 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 245106 0 245162 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 248326 0 248382 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 251454 0 251510 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 254582 0 254638 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 257802 0 257858 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 260930 0 260986 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 264150 0 264206 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 267278 0 267334 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 270406 0 270462 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 273626 0 273682 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 276754 0 276810 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 283102 0 283158 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 286230 0 286286 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 289450 0 289506 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 292578 0 292634 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 295798 0 295854 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 298926 0 298982 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 302054 0 302110 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 305274 0 305330 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 308402 0 308458 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 311622 0 311678 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 314750 0 314806 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 317878 0 317934 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 321098 0 321154 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 324226 0 324282 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 327354 0 327410 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 330574 0 330630 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 333702 0 333758 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 336922 0 336978 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 343178 0 343234 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 346398 0 346454 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 349526 0 349582 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 352746 0 352802 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 355874 0 355930 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 359002 0 359058 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 362222 0 362278 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 365350 0 365406 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 368570 0 368626 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 371698 0 371754 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 374826 0 374882 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 378046 0 378102 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 381174 0 381230 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 384394 0 384450 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 387522 0 387578 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 390650 0 390706 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 393870 0 393926 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 396998 0 397054 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 400218 0 400274 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 403346 0 403402 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 406474 0 406530 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 409694 0 409750 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 412822 0 412878 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 416042 0 416098 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 419170 0 419226 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 422298 0 422354 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 425518 0 425574 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 429750 0 429806 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 432878 0 432934 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 436006 0 436062 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 439226 0 439282 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 442354 0 442410 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 445574 0 445630 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 448702 0 448758 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 451830 0 451886 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 455050 0 455106 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 458178 0 458234 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 461306 0 461362 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 464526 0 464582 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 467654 0 467710 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 470874 0 470930 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 474002 0 474058 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 477130 0 477186 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 480350 0 480406 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 483478 0 483534 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 486698 0 486754 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 489826 0 489882 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 492954 0 493010 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 496174 0 496230 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 499302 0 499358 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 502522 0 502578 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 505650 0 505706 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 508778 0 508834 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 511998 0 512054 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 515126 0 515182 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 151266 0 151322 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 160742 0 160798 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 167090 0 167146 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 170218 0 170274 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 173438 0 173494 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 182914 0 182970 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 186042 0 186098 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 189262 0 189318 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 192390 0 192446 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 195518 0 195574 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 198738 0 198794 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 201866 0 201922 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 205086 0 205142 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 208214 0 208270 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 211342 0 211398 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 214562 0 214618 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 220910 0 220966 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 227166 0 227222 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 230386 0 230442 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 233514 0 233570 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 236734 0 236790 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 239862 0 239918 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 242990 0 243046 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 246210 0 246266 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 249338 0 249394 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 252558 0 252614 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 255686 0 255742 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 258814 0 258870 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 262034 0 262090 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 265162 0 265218 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 268290 0 268346 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 271510 0 271566 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 274638 0 274694 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 277858 0 277914 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 280986 0 281042 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 284114 0 284170 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 287334 0 287390 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 290462 0 290518 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 293682 0 293738 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 296810 0 296866 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 299938 0 299994 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 303158 0 303214 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 306286 0 306342 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 309506 0 309562 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 312634 0 312690 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 315762 0 315818 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 318982 0 319038 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 322110 0 322166 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 325330 0 325386 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 328458 0 328514 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 331586 0 331642 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 334806 0 334862 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 337934 0 337990 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 341154 0 341210 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 344282 0 344338 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 347410 0 347466 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 350630 0 350686 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 353758 0 353814 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 356978 0 357034 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 360106 0 360162 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 363234 0 363290 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 366454 0 366510 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 369582 0 369638 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 372710 0 372766 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 375930 0 375986 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 379058 0 379114 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 382278 0 382334 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 385406 0 385462 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 388534 0 388590 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 391754 0 391810 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 394882 0 394938 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 398102 0 398158 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 401230 0 401286 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 404358 0 404414 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 407578 0 407634 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 410706 0 410762 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 413926 0 413982 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 417054 0 417110 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 420182 0 420238 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 423402 0 423458 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 426530 0 426586 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 430762 0 430818 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 433890 0 433946 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 437110 0 437166 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 440238 0 440294 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 443458 0 443514 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 446586 0 446642 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 449714 0 449770 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 452934 0 452990 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 456062 0 456118 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 459282 0 459338 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 462410 0 462466 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 465538 0 465594 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 468758 0 468814 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 471886 0 471942 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 475106 0 475162 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 478234 0 478290 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 481362 0 481418 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 484582 0 484638 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 487710 0 487766 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 490838 0 490894 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 494058 0 494114 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 497186 0 497242 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 500406 0 500462 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 503534 0 503590 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 506662 0 506718 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 509882 0 509938 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 513010 0 513066 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 516230 0 516286 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 202970 0 203026 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 209226 0 209282 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 215574 0 215630 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 221922 0 221978 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 231398 0 231454 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 234618 0 234674 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 237746 0 237802 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 240874 0 240930 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 247222 0 247278 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 250442 0 250498 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 253570 0 253626 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 256698 0 256754 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 259918 0 259974 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 266266 0 266322 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 269394 0 269450 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 272522 0 272578 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 278870 0 278926 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 282090 0 282146 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 285218 0 285274 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 288346 0 288402 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 294694 0 294750 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 301042 0 301098 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 304170 0 304226 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 307390 0 307446 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 310518 0 310574 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 313646 0 313702 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 316866 0 316922 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 319994 0 320050 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 323214 0 323270 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 326342 0 326398 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 329470 0 329526 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 332690 0 332746 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 335818 0 335874 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 339038 0 339094 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 342166 0 342222 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 345294 0 345350 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 348514 0 348570 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 351642 0 351698 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 354862 0 354918 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 357990 0 358046 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 361118 0 361174 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 364338 0 364394 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 367466 0 367522 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 370686 0 370742 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 373814 0 373870 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 376942 0 376998 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 380162 0 380218 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 383290 0 383346 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 386510 0 386566 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 389638 0 389694 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 392766 0 392822 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 395986 0 396042 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 399114 0 399170 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 402242 0 402298 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 405462 0 405518 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 408590 0 408646 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 411810 0 411866 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 414938 0 414994 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 418066 0 418122 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 421286 0 421342 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 424414 0 424470 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 427634 0 427690 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 434288 2128 434608 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 465008 2128 465328 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 495728 2128 496048 637616 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 418928 2128 419248 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 449648 2128 449968 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 480368 2128 480688 637616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 511088 2128 511408 637616 6 vssd1
port 503 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 520000 640000
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 894537314
string GDS_START 1479438
<< end >>

